magic
tech gf180mcuC
magscale 1 10
timestamp 1676577649
<< error_p >>
rect -27407 3555 -27363 3563
rect -27307 3555 -27263 3563
rect -27207 3555 -27163 3563
rect -27107 3555 -27063 3563
rect -27007 3555 -26963 3563
rect -26907 3555 -26863 3563
rect -26807 3555 -26763 3563
rect -26707 3555 -26663 3563
rect -26607 3555 -26563 3563
rect -26507 3555 -26463 3563
rect -26407 3555 -26363 3563
rect -26307 3555 -26263 3563
rect -26207 3555 -26163 3563
rect -26107 3555 -26063 3563
rect -26007 3555 -25963 3563
rect -25907 3555 -25863 3563
rect -25407 3555 -25363 3563
rect -25307 3555 -25263 3563
rect -25207 3555 -25163 3563
rect -25107 3555 -25063 3563
rect -25007 3555 -24963 3563
rect -24907 3555 -24863 3563
rect -24807 3555 -24763 3563
rect -24707 3555 -24663 3563
rect -24607 3555 -24563 3563
rect -24507 3555 -24463 3563
rect -24407 3555 -24363 3563
rect -24307 3555 -24263 3563
rect -24207 3555 -24163 3563
rect -24107 3555 -24063 3563
rect -24007 3555 -23963 3563
rect -23907 3555 -23863 3563
rect -23407 3555 -23363 3563
rect -23307 3555 -23263 3563
rect -23207 3555 -23163 3563
rect -23107 3555 -23063 3563
rect -23007 3555 -22963 3563
rect -22907 3555 -22863 3563
rect -22807 3555 -22763 3563
rect -22707 3555 -22663 3563
rect -22607 3555 -22563 3563
rect -22507 3555 -22463 3563
rect -22407 3555 -22363 3563
rect -22307 3555 -22263 3563
rect -22207 3555 -22163 3563
rect -22107 3555 -22063 3563
rect -22007 3555 -21963 3563
rect -21907 3555 -21863 3563
rect -21407 3555 -21363 3563
rect -21307 3555 -21263 3563
rect -21207 3555 -21163 3563
rect -21107 3555 -21063 3563
rect -21007 3555 -20963 3563
rect -20907 3555 -20863 3563
rect -20807 3555 -20763 3563
rect -20707 3555 -20663 3563
rect -20607 3555 -20563 3563
rect -20507 3555 -20463 3563
rect -20407 3555 -20363 3563
rect -20307 3555 -20263 3563
rect -20207 3555 -20163 3563
rect -20107 3555 -20063 3563
rect -20007 3555 -19963 3563
rect -19907 3555 -19863 3563
rect -27363 3511 -27355 3555
rect -27263 3511 -27255 3555
rect -27163 3511 -27155 3555
rect -27063 3511 -27055 3555
rect -26963 3511 -26955 3555
rect -26863 3511 -26855 3555
rect -26763 3511 -26755 3555
rect -26663 3511 -26655 3555
rect -26563 3511 -26555 3555
rect -26463 3511 -26455 3555
rect -26363 3511 -26355 3555
rect -26263 3511 -26255 3555
rect -26163 3511 -26155 3555
rect -26063 3511 -26055 3555
rect -25963 3511 -25955 3555
rect -25863 3511 -25855 3555
rect -25363 3511 -25355 3555
rect -25263 3511 -25255 3555
rect -25163 3511 -25155 3555
rect -25063 3511 -25055 3555
rect -24963 3511 -24955 3555
rect -24863 3511 -24855 3555
rect -24763 3511 -24755 3555
rect -24663 3511 -24655 3555
rect -24563 3511 -24555 3555
rect -24463 3511 -24455 3555
rect -24363 3511 -24355 3555
rect -24263 3511 -24255 3555
rect -24163 3511 -24155 3555
rect -24063 3511 -24055 3555
rect -23963 3511 -23955 3555
rect -23863 3511 -23855 3555
rect -23363 3511 -23355 3555
rect -23263 3511 -23255 3555
rect -23163 3511 -23155 3555
rect -23063 3511 -23055 3555
rect -22963 3511 -22955 3555
rect -22863 3511 -22855 3555
rect -22763 3511 -22755 3555
rect -22663 3511 -22655 3555
rect -22563 3511 -22555 3555
rect -22463 3511 -22455 3555
rect -22363 3511 -22355 3555
rect -22263 3511 -22255 3555
rect -22163 3511 -22155 3555
rect -22063 3511 -22055 3555
rect -21963 3511 -21955 3555
rect -21863 3511 -21855 3555
rect -21363 3511 -21355 3555
rect -21263 3511 -21255 3555
rect -21163 3511 -21155 3555
rect -21063 3511 -21055 3555
rect -20963 3511 -20955 3555
rect -20863 3511 -20855 3555
rect -20763 3511 -20755 3555
rect -20663 3511 -20655 3555
rect -20563 3511 -20555 3555
rect -20463 3511 -20455 3555
rect -20363 3511 -20355 3555
rect -20263 3511 -20255 3555
rect -20163 3511 -20155 3555
rect -20063 3511 -20055 3555
rect -19963 3511 -19955 3555
rect -19863 3511 -19855 3555
rect -27407 3455 -27363 3463
rect -27307 3455 -27263 3463
rect -27207 3455 -27163 3463
rect -27107 3455 -27063 3463
rect -27007 3455 -26963 3463
rect -26907 3455 -26863 3463
rect -26807 3455 -26763 3463
rect -26707 3455 -26663 3463
rect -26607 3455 -26563 3463
rect -26507 3455 -26463 3463
rect -26407 3455 -26363 3463
rect -26307 3455 -26263 3463
rect -26207 3455 -26163 3463
rect -26107 3455 -26063 3463
rect -26007 3455 -25963 3463
rect -25907 3455 -25863 3463
rect -25407 3455 -25363 3463
rect -25307 3455 -25263 3463
rect -25207 3455 -25163 3463
rect -25107 3455 -25063 3463
rect -25007 3455 -24963 3463
rect -24907 3455 -24863 3463
rect -24807 3455 -24763 3463
rect -24707 3455 -24663 3463
rect -24607 3455 -24563 3463
rect -24507 3455 -24463 3463
rect -24407 3455 -24363 3463
rect -24307 3455 -24263 3463
rect -24207 3455 -24163 3463
rect -24107 3455 -24063 3463
rect -24007 3455 -23963 3463
rect -23907 3455 -23863 3463
rect -23407 3455 -23363 3463
rect -23307 3455 -23263 3463
rect -23207 3455 -23163 3463
rect -23107 3455 -23063 3463
rect -23007 3455 -22963 3463
rect -22907 3455 -22863 3463
rect -22807 3455 -22763 3463
rect -22707 3455 -22663 3463
rect -22607 3455 -22563 3463
rect -22507 3455 -22463 3463
rect -22407 3455 -22363 3463
rect -22307 3455 -22263 3463
rect -22207 3455 -22163 3463
rect -22107 3455 -22063 3463
rect -22007 3455 -21963 3463
rect -21907 3455 -21863 3463
rect -21407 3455 -21363 3463
rect -21307 3455 -21263 3463
rect -21207 3455 -21163 3463
rect -21107 3455 -21063 3463
rect -21007 3455 -20963 3463
rect -20907 3455 -20863 3463
rect -20807 3455 -20763 3463
rect -20707 3455 -20663 3463
rect -20607 3455 -20563 3463
rect -20507 3455 -20463 3463
rect -20407 3455 -20363 3463
rect -20307 3455 -20263 3463
rect -20207 3455 -20163 3463
rect -20107 3455 -20063 3463
rect -20007 3455 -19963 3463
rect -19907 3455 -19863 3463
rect -27363 3411 -27355 3455
rect -27263 3411 -27255 3455
rect -27163 3411 -27155 3455
rect -27063 3411 -27055 3455
rect -26963 3411 -26955 3455
rect -26863 3411 -26855 3455
rect -26763 3411 -26755 3455
rect -26663 3411 -26655 3455
rect -26563 3411 -26555 3455
rect -26463 3411 -26455 3455
rect -26363 3411 -26355 3455
rect -26263 3411 -26255 3455
rect -26163 3411 -26155 3455
rect -26063 3411 -26055 3455
rect -25963 3411 -25955 3455
rect -25863 3411 -25855 3455
rect -25363 3411 -25355 3455
rect -25263 3411 -25255 3455
rect -25163 3411 -25155 3455
rect -25063 3411 -25055 3455
rect -24963 3411 -24955 3455
rect -24863 3411 -24855 3455
rect -24763 3411 -24755 3455
rect -24663 3411 -24655 3455
rect -24563 3411 -24555 3455
rect -24463 3411 -24455 3455
rect -24363 3411 -24355 3455
rect -24263 3411 -24255 3455
rect -24163 3411 -24155 3455
rect -24063 3411 -24055 3455
rect -23963 3411 -23955 3455
rect -23863 3411 -23855 3455
rect -23363 3411 -23355 3455
rect -23263 3411 -23255 3455
rect -23163 3411 -23155 3455
rect -23063 3411 -23055 3455
rect -22963 3411 -22955 3455
rect -22863 3411 -22855 3455
rect -22763 3411 -22755 3455
rect -22663 3411 -22655 3455
rect -22563 3411 -22555 3455
rect -22463 3411 -22455 3455
rect -22363 3411 -22355 3455
rect -22263 3411 -22255 3455
rect -22163 3411 -22155 3455
rect -22063 3411 -22055 3455
rect -21963 3411 -21955 3455
rect -21863 3411 -21855 3455
rect -21363 3411 -21355 3455
rect -21263 3411 -21255 3455
rect -21163 3411 -21155 3455
rect -21063 3411 -21055 3455
rect -20963 3411 -20955 3455
rect -20863 3411 -20855 3455
rect -20763 3411 -20755 3455
rect -20663 3411 -20655 3455
rect -20563 3411 -20555 3455
rect -20463 3411 -20455 3455
rect -20363 3411 -20355 3455
rect -20263 3411 -20255 3455
rect -20163 3411 -20155 3455
rect -20063 3411 -20055 3455
rect -19963 3411 -19955 3455
rect -19863 3411 -19855 3455
rect -27407 3355 -27363 3363
rect -27307 3355 -27263 3363
rect -27207 3355 -27163 3363
rect -27107 3355 -27063 3363
rect -27007 3355 -26963 3363
rect -26907 3355 -26863 3363
rect -26807 3355 -26763 3363
rect -26707 3355 -26663 3363
rect -26607 3355 -26563 3363
rect -26507 3355 -26463 3363
rect -26407 3355 -26363 3363
rect -26307 3355 -26263 3363
rect -26207 3355 -26163 3363
rect -26107 3355 -26063 3363
rect -26007 3355 -25963 3363
rect -25907 3355 -25863 3363
rect -25407 3355 -25363 3363
rect -25307 3355 -25263 3363
rect -25207 3355 -25163 3363
rect -25107 3355 -25063 3363
rect -25007 3355 -24963 3363
rect -24907 3355 -24863 3363
rect -24807 3355 -24763 3363
rect -24707 3355 -24663 3363
rect -24607 3355 -24563 3363
rect -24507 3355 -24463 3363
rect -24407 3355 -24363 3363
rect -24307 3355 -24263 3363
rect -24207 3355 -24163 3363
rect -24107 3355 -24063 3363
rect -24007 3355 -23963 3363
rect -23907 3355 -23863 3363
rect -23407 3355 -23363 3363
rect -23307 3355 -23263 3363
rect -23207 3355 -23163 3363
rect -23107 3355 -23063 3363
rect -23007 3355 -22963 3363
rect -22907 3355 -22863 3363
rect -22807 3355 -22763 3363
rect -22707 3355 -22663 3363
rect -22607 3355 -22563 3363
rect -22507 3355 -22463 3363
rect -22407 3355 -22363 3363
rect -22307 3355 -22263 3363
rect -22207 3355 -22163 3363
rect -22107 3355 -22063 3363
rect -22007 3355 -21963 3363
rect -21907 3355 -21863 3363
rect -21407 3355 -21363 3363
rect -21307 3355 -21263 3363
rect -21207 3355 -21163 3363
rect -21107 3355 -21063 3363
rect -21007 3355 -20963 3363
rect -20907 3355 -20863 3363
rect -20807 3355 -20763 3363
rect -20707 3355 -20663 3363
rect -20607 3355 -20563 3363
rect -20507 3355 -20463 3363
rect -20407 3355 -20363 3363
rect -20307 3355 -20263 3363
rect -20207 3355 -20163 3363
rect -20107 3355 -20063 3363
rect -20007 3355 -19963 3363
rect -19907 3355 -19863 3363
rect -27363 3311 -27355 3355
rect -27263 3311 -27255 3355
rect -27163 3311 -27155 3355
rect -27063 3311 -27055 3355
rect -26963 3311 -26955 3355
rect -26863 3311 -26855 3355
rect -26763 3311 -26755 3355
rect -26663 3311 -26655 3355
rect -26563 3311 -26555 3355
rect -26463 3311 -26455 3355
rect -26363 3311 -26355 3355
rect -26263 3311 -26255 3355
rect -26163 3311 -26155 3355
rect -26063 3311 -26055 3355
rect -25963 3311 -25955 3355
rect -25863 3311 -25855 3355
rect -25363 3311 -25355 3355
rect -25263 3311 -25255 3355
rect -25163 3311 -25155 3355
rect -25063 3311 -25055 3355
rect -24963 3311 -24955 3355
rect -24863 3311 -24855 3355
rect -24763 3311 -24755 3355
rect -24663 3311 -24655 3355
rect -24563 3311 -24555 3355
rect -24463 3311 -24455 3355
rect -24363 3311 -24355 3355
rect -24263 3311 -24255 3355
rect -24163 3311 -24155 3355
rect -24063 3311 -24055 3355
rect -23963 3311 -23955 3355
rect -23863 3311 -23855 3355
rect -23363 3311 -23355 3355
rect -23263 3311 -23255 3355
rect -23163 3311 -23155 3355
rect -23063 3311 -23055 3355
rect -22963 3311 -22955 3355
rect -22863 3311 -22855 3355
rect -22763 3311 -22755 3355
rect -22663 3311 -22655 3355
rect -22563 3311 -22555 3355
rect -22463 3311 -22455 3355
rect -22363 3311 -22355 3355
rect -22263 3311 -22255 3355
rect -22163 3311 -22155 3355
rect -22063 3311 -22055 3355
rect -21963 3311 -21955 3355
rect -21863 3311 -21855 3355
rect -21363 3311 -21355 3355
rect -21263 3311 -21255 3355
rect -21163 3311 -21155 3355
rect -21063 3311 -21055 3355
rect -20963 3311 -20955 3355
rect -20863 3311 -20855 3355
rect -20763 3311 -20755 3355
rect -20663 3311 -20655 3355
rect -20563 3311 -20555 3355
rect -20463 3311 -20455 3355
rect -20363 3311 -20355 3355
rect -20263 3311 -20255 3355
rect -20163 3311 -20155 3355
rect -20063 3311 -20055 3355
rect -19963 3311 -19955 3355
rect -19863 3311 -19855 3355
rect -27407 3255 -27363 3263
rect -27307 3255 -27263 3263
rect -27207 3255 -27163 3263
rect -27107 3255 -27063 3263
rect -27007 3255 -26963 3263
rect -26907 3255 -26863 3263
rect -26807 3255 -26763 3263
rect -26707 3255 -26663 3263
rect -26607 3255 -26563 3263
rect -26507 3255 -26463 3263
rect -26407 3255 -26363 3263
rect -26307 3255 -26263 3263
rect -26207 3255 -26163 3263
rect -26107 3255 -26063 3263
rect -26007 3255 -25963 3263
rect -25907 3255 -25863 3263
rect -25407 3255 -25363 3263
rect -25307 3255 -25263 3263
rect -25207 3255 -25163 3263
rect -25107 3255 -25063 3263
rect -25007 3255 -24963 3263
rect -24907 3255 -24863 3263
rect -24807 3255 -24763 3263
rect -24707 3255 -24663 3263
rect -24607 3255 -24563 3263
rect -24507 3255 -24463 3263
rect -24407 3255 -24363 3263
rect -24307 3255 -24263 3263
rect -24207 3255 -24163 3263
rect -24107 3255 -24063 3263
rect -24007 3255 -23963 3263
rect -23907 3255 -23863 3263
rect -23407 3255 -23363 3263
rect -23307 3255 -23263 3263
rect -23207 3255 -23163 3263
rect -23107 3255 -23063 3263
rect -23007 3255 -22963 3263
rect -22907 3255 -22863 3263
rect -22807 3255 -22763 3263
rect -22707 3255 -22663 3263
rect -22607 3255 -22563 3263
rect -22507 3255 -22463 3263
rect -22407 3255 -22363 3263
rect -22307 3255 -22263 3263
rect -22207 3255 -22163 3263
rect -22107 3255 -22063 3263
rect -22007 3255 -21963 3263
rect -21907 3255 -21863 3263
rect -21407 3255 -21363 3263
rect -21307 3255 -21263 3263
rect -21207 3255 -21163 3263
rect -21107 3255 -21063 3263
rect -21007 3255 -20963 3263
rect -20907 3255 -20863 3263
rect -20807 3255 -20763 3263
rect -20707 3255 -20663 3263
rect -20607 3255 -20563 3263
rect -20507 3255 -20463 3263
rect -20407 3255 -20363 3263
rect -20307 3255 -20263 3263
rect -20207 3255 -20163 3263
rect -20107 3255 -20063 3263
rect -20007 3255 -19963 3263
rect -19907 3255 -19863 3263
rect -27363 3211 -27355 3255
rect -27263 3211 -27255 3255
rect -27163 3211 -27155 3255
rect -27063 3211 -27055 3255
rect -26963 3211 -26955 3255
rect -26863 3211 -26855 3255
rect -26763 3211 -26755 3255
rect -26663 3211 -26655 3255
rect -26563 3211 -26555 3255
rect -26463 3211 -26455 3255
rect -26363 3211 -26355 3255
rect -26263 3211 -26255 3255
rect -26163 3211 -26155 3255
rect -26063 3211 -26055 3255
rect -25963 3211 -25955 3255
rect -25863 3211 -25855 3255
rect -25363 3211 -25355 3255
rect -25263 3211 -25255 3255
rect -25163 3211 -25155 3255
rect -25063 3211 -25055 3255
rect -24963 3211 -24955 3255
rect -24863 3211 -24855 3255
rect -24763 3211 -24755 3255
rect -24663 3211 -24655 3255
rect -24563 3211 -24555 3255
rect -24463 3211 -24455 3255
rect -24363 3211 -24355 3255
rect -24263 3211 -24255 3255
rect -24163 3211 -24155 3255
rect -24063 3211 -24055 3255
rect -23963 3211 -23955 3255
rect -23863 3211 -23855 3255
rect -23363 3211 -23355 3255
rect -23263 3211 -23255 3255
rect -23163 3211 -23155 3255
rect -23063 3211 -23055 3255
rect -22963 3211 -22955 3255
rect -22863 3211 -22855 3255
rect -22763 3211 -22755 3255
rect -22663 3211 -22655 3255
rect -22563 3211 -22555 3255
rect -22463 3211 -22455 3255
rect -22363 3211 -22355 3255
rect -22263 3211 -22255 3255
rect -22163 3211 -22155 3255
rect -22063 3211 -22055 3255
rect -21963 3211 -21955 3255
rect -21863 3211 -21855 3255
rect -21363 3211 -21355 3255
rect -21263 3211 -21255 3255
rect -21163 3211 -21155 3255
rect -21063 3211 -21055 3255
rect -20963 3211 -20955 3255
rect -20863 3211 -20855 3255
rect -20763 3211 -20755 3255
rect -20663 3211 -20655 3255
rect -20563 3211 -20555 3255
rect -20463 3211 -20455 3255
rect -20363 3211 -20355 3255
rect -20263 3211 -20255 3255
rect -20163 3211 -20155 3255
rect -20063 3211 -20055 3255
rect -19963 3211 -19955 3255
rect -19863 3211 -19855 3255
rect -27407 3155 -27363 3163
rect -27307 3155 -27263 3163
rect -27207 3155 -27163 3163
rect -27107 3155 -27063 3163
rect -27007 3155 -26963 3163
rect -26907 3155 -26863 3163
rect -26807 3155 -26763 3163
rect -26707 3155 -26663 3163
rect -26607 3155 -26563 3163
rect -26507 3155 -26463 3163
rect -26407 3155 -26363 3163
rect -26307 3155 -26263 3163
rect -26207 3155 -26163 3163
rect -26107 3155 -26063 3163
rect -26007 3155 -25963 3163
rect -25907 3155 -25863 3163
rect -25407 3155 -25363 3163
rect -25307 3155 -25263 3163
rect -25207 3155 -25163 3163
rect -25107 3155 -25063 3163
rect -25007 3155 -24963 3163
rect -24907 3155 -24863 3163
rect -24807 3155 -24763 3163
rect -24707 3155 -24663 3163
rect -24607 3155 -24563 3163
rect -24507 3155 -24463 3163
rect -24407 3155 -24363 3163
rect -24307 3155 -24263 3163
rect -24207 3155 -24163 3163
rect -24107 3155 -24063 3163
rect -24007 3155 -23963 3163
rect -23907 3155 -23863 3163
rect -23407 3155 -23363 3163
rect -23307 3155 -23263 3163
rect -23207 3155 -23163 3163
rect -23107 3155 -23063 3163
rect -23007 3155 -22963 3163
rect -22907 3155 -22863 3163
rect -22807 3155 -22763 3163
rect -22707 3155 -22663 3163
rect -22607 3155 -22563 3163
rect -22507 3155 -22463 3163
rect -22407 3155 -22363 3163
rect -22307 3155 -22263 3163
rect -22207 3155 -22163 3163
rect -22107 3155 -22063 3163
rect -22007 3155 -21963 3163
rect -21907 3155 -21863 3163
rect -21407 3155 -21363 3163
rect -21307 3155 -21263 3163
rect -21207 3155 -21163 3163
rect -21107 3155 -21063 3163
rect -21007 3155 -20963 3163
rect -20907 3155 -20863 3163
rect -20807 3155 -20763 3163
rect -20707 3155 -20663 3163
rect -20607 3155 -20563 3163
rect -20507 3155 -20463 3163
rect -20407 3155 -20363 3163
rect -20307 3155 -20263 3163
rect -20207 3155 -20163 3163
rect -20107 3155 -20063 3163
rect -20007 3155 -19963 3163
rect -19907 3155 -19863 3163
rect -27363 3111 -27355 3155
rect -27263 3111 -27255 3155
rect -27163 3111 -27155 3155
rect -27063 3111 -27055 3155
rect -26963 3111 -26955 3155
rect -26863 3111 -26855 3155
rect -26763 3111 -26755 3155
rect -26663 3111 -26655 3155
rect -26563 3111 -26555 3155
rect -26463 3111 -26455 3155
rect -26363 3111 -26355 3155
rect -26263 3111 -26255 3155
rect -26163 3111 -26155 3155
rect -26063 3111 -26055 3155
rect -25963 3111 -25955 3155
rect -25863 3111 -25855 3155
rect -25363 3111 -25355 3155
rect -25263 3111 -25255 3155
rect -25163 3111 -25155 3155
rect -25063 3111 -25055 3155
rect -24963 3111 -24955 3155
rect -24863 3111 -24855 3155
rect -24763 3111 -24755 3155
rect -24663 3111 -24655 3155
rect -24563 3111 -24555 3155
rect -24463 3111 -24455 3155
rect -24363 3111 -24355 3155
rect -24263 3111 -24255 3155
rect -24163 3111 -24155 3155
rect -24063 3111 -24055 3155
rect -23963 3111 -23955 3155
rect -23863 3111 -23855 3155
rect -23363 3111 -23355 3155
rect -23263 3111 -23255 3155
rect -23163 3111 -23155 3155
rect -23063 3111 -23055 3155
rect -22963 3111 -22955 3155
rect -22863 3111 -22855 3155
rect -22763 3111 -22755 3155
rect -22663 3111 -22655 3155
rect -22563 3111 -22555 3155
rect -22463 3111 -22455 3155
rect -22363 3111 -22355 3155
rect -22263 3111 -22255 3155
rect -22163 3111 -22155 3155
rect -22063 3111 -22055 3155
rect -21963 3111 -21955 3155
rect -21863 3111 -21855 3155
rect -21363 3111 -21355 3155
rect -21263 3111 -21255 3155
rect -21163 3111 -21155 3155
rect -21063 3111 -21055 3155
rect -20963 3111 -20955 3155
rect -20863 3111 -20855 3155
rect -20763 3111 -20755 3155
rect -20663 3111 -20655 3155
rect -20563 3111 -20555 3155
rect -20463 3111 -20455 3155
rect -20363 3111 -20355 3155
rect -20263 3111 -20255 3155
rect -20163 3111 -20155 3155
rect -20063 3111 -20055 3155
rect -19963 3111 -19955 3155
rect -19863 3111 -19855 3155
rect -27407 3055 -27363 3063
rect -27307 3055 -27263 3063
rect -27207 3055 -27163 3063
rect -27107 3055 -27063 3063
rect -27007 3055 -26963 3063
rect -26907 3055 -26863 3063
rect -26807 3055 -26763 3063
rect -26707 3055 -26663 3063
rect -26607 3055 -26563 3063
rect -26507 3055 -26463 3063
rect -26407 3055 -26363 3063
rect -26307 3055 -26263 3063
rect -26207 3055 -26163 3063
rect -26107 3055 -26063 3063
rect -26007 3055 -25963 3063
rect -25907 3055 -25863 3063
rect -25407 3055 -25363 3063
rect -25307 3055 -25263 3063
rect -25207 3055 -25163 3063
rect -25107 3055 -25063 3063
rect -25007 3055 -24963 3063
rect -24907 3055 -24863 3063
rect -24807 3055 -24763 3063
rect -24707 3055 -24663 3063
rect -24607 3055 -24563 3063
rect -24507 3055 -24463 3063
rect -24407 3055 -24363 3063
rect -24307 3055 -24263 3063
rect -24207 3055 -24163 3063
rect -24107 3055 -24063 3063
rect -24007 3055 -23963 3063
rect -23907 3055 -23863 3063
rect -23407 3055 -23363 3063
rect -23307 3055 -23263 3063
rect -23207 3055 -23163 3063
rect -23107 3055 -23063 3063
rect -23007 3055 -22963 3063
rect -22907 3055 -22863 3063
rect -22807 3055 -22763 3063
rect -22707 3055 -22663 3063
rect -22607 3055 -22563 3063
rect -22507 3055 -22463 3063
rect -22407 3055 -22363 3063
rect -22307 3055 -22263 3063
rect -22207 3055 -22163 3063
rect -22107 3055 -22063 3063
rect -22007 3055 -21963 3063
rect -21907 3055 -21863 3063
rect -21407 3055 -21363 3063
rect -21307 3055 -21263 3063
rect -21207 3055 -21163 3063
rect -21107 3055 -21063 3063
rect -21007 3055 -20963 3063
rect -20907 3055 -20863 3063
rect -20807 3055 -20763 3063
rect -20707 3055 -20663 3063
rect -20607 3055 -20563 3063
rect -20507 3055 -20463 3063
rect -20407 3055 -20363 3063
rect -20307 3055 -20263 3063
rect -20207 3055 -20163 3063
rect -20107 3055 -20063 3063
rect -20007 3055 -19963 3063
rect -19907 3055 -19863 3063
rect -27363 3011 -27355 3055
rect -27263 3011 -27255 3055
rect -27163 3011 -27155 3055
rect -27063 3011 -27055 3055
rect -26963 3011 -26955 3055
rect -26863 3011 -26855 3055
rect -26763 3011 -26755 3055
rect -26663 3011 -26655 3055
rect -26563 3011 -26555 3055
rect -26463 3011 -26455 3055
rect -26363 3011 -26355 3055
rect -26263 3011 -26255 3055
rect -26163 3011 -26155 3055
rect -26063 3011 -26055 3055
rect -25963 3011 -25955 3055
rect -25863 3011 -25855 3055
rect -25363 3011 -25355 3055
rect -25263 3011 -25255 3055
rect -25163 3011 -25155 3055
rect -25063 3011 -25055 3055
rect -24963 3011 -24955 3055
rect -24863 3011 -24855 3055
rect -24763 3011 -24755 3055
rect -24663 3011 -24655 3055
rect -24563 3011 -24555 3055
rect -24463 3011 -24455 3055
rect -24363 3011 -24355 3055
rect -24263 3011 -24255 3055
rect -24163 3011 -24155 3055
rect -24063 3011 -24055 3055
rect -23963 3011 -23955 3055
rect -23863 3011 -23855 3055
rect -23363 3011 -23355 3055
rect -23263 3011 -23255 3055
rect -23163 3011 -23155 3055
rect -23063 3011 -23055 3055
rect -22963 3011 -22955 3055
rect -22863 3011 -22855 3055
rect -22763 3011 -22755 3055
rect -22663 3011 -22655 3055
rect -22563 3011 -22555 3055
rect -22463 3011 -22455 3055
rect -22363 3011 -22355 3055
rect -22263 3011 -22255 3055
rect -22163 3011 -22155 3055
rect -22063 3011 -22055 3055
rect -21963 3011 -21955 3055
rect -21863 3011 -21855 3055
rect -21363 3011 -21355 3055
rect -21263 3011 -21255 3055
rect -21163 3011 -21155 3055
rect -21063 3011 -21055 3055
rect -20963 3011 -20955 3055
rect -20863 3011 -20855 3055
rect -20763 3011 -20755 3055
rect -20663 3011 -20655 3055
rect -20563 3011 -20555 3055
rect -20463 3011 -20455 3055
rect -20363 3011 -20355 3055
rect -20263 3011 -20255 3055
rect -20163 3011 -20155 3055
rect -20063 3011 -20055 3055
rect -19963 3011 -19955 3055
rect -19863 3011 -19855 3055
rect -27407 2955 -27363 2963
rect -27307 2955 -27263 2963
rect -27207 2955 -27163 2963
rect -27107 2955 -27063 2963
rect -27007 2955 -26963 2963
rect -26907 2955 -26863 2963
rect -26807 2955 -26763 2963
rect -26707 2955 -26663 2963
rect -26607 2955 -26563 2963
rect -26507 2955 -26463 2963
rect -26407 2955 -26363 2963
rect -26307 2955 -26263 2963
rect -26207 2955 -26163 2963
rect -26107 2955 -26063 2963
rect -26007 2955 -25963 2963
rect -25907 2955 -25863 2963
rect -25407 2955 -25363 2963
rect -25307 2955 -25263 2963
rect -25207 2955 -25163 2963
rect -25107 2955 -25063 2963
rect -25007 2955 -24963 2963
rect -24907 2955 -24863 2963
rect -24807 2955 -24763 2963
rect -24707 2955 -24663 2963
rect -24607 2955 -24563 2963
rect -24507 2955 -24463 2963
rect -24407 2955 -24363 2963
rect -24307 2955 -24263 2963
rect -24207 2955 -24163 2963
rect -24107 2955 -24063 2963
rect -24007 2955 -23963 2963
rect -23907 2955 -23863 2963
rect -23407 2955 -23363 2963
rect -23307 2955 -23263 2963
rect -23207 2955 -23163 2963
rect -23107 2955 -23063 2963
rect -23007 2955 -22963 2963
rect -22907 2955 -22863 2963
rect -22807 2955 -22763 2963
rect -22707 2955 -22663 2963
rect -22607 2955 -22563 2963
rect -22507 2955 -22463 2963
rect -22407 2955 -22363 2963
rect -22307 2955 -22263 2963
rect -22207 2955 -22163 2963
rect -22107 2955 -22063 2963
rect -22007 2955 -21963 2963
rect -21907 2955 -21863 2963
rect -21407 2955 -21363 2963
rect -21307 2955 -21263 2963
rect -21207 2955 -21163 2963
rect -21107 2955 -21063 2963
rect -21007 2955 -20963 2963
rect -20907 2955 -20863 2963
rect -20807 2955 -20763 2963
rect -20707 2955 -20663 2963
rect -20607 2955 -20563 2963
rect -20507 2955 -20463 2963
rect -20407 2955 -20363 2963
rect -20307 2955 -20263 2963
rect -20207 2955 -20163 2963
rect -20107 2955 -20063 2963
rect -20007 2955 -19963 2963
rect -19907 2955 -19863 2963
rect -27363 2911 -27355 2955
rect -27263 2911 -27255 2955
rect -27163 2911 -27155 2955
rect -27063 2911 -27055 2955
rect -26963 2911 -26955 2955
rect -26863 2911 -26855 2955
rect -26763 2911 -26755 2955
rect -26663 2911 -26655 2955
rect -26563 2911 -26555 2955
rect -26463 2911 -26455 2955
rect -26363 2911 -26355 2955
rect -26263 2911 -26255 2955
rect -26163 2911 -26155 2955
rect -26063 2911 -26055 2955
rect -25963 2911 -25955 2955
rect -25863 2911 -25855 2955
rect -25363 2911 -25355 2955
rect -25263 2911 -25255 2955
rect -25163 2911 -25155 2955
rect -25063 2911 -25055 2955
rect -24963 2911 -24955 2955
rect -24863 2911 -24855 2955
rect -24763 2911 -24755 2955
rect -24663 2911 -24655 2955
rect -24563 2911 -24555 2955
rect -24463 2911 -24455 2955
rect -24363 2911 -24355 2955
rect -24263 2911 -24255 2955
rect -24163 2911 -24155 2955
rect -24063 2911 -24055 2955
rect -23963 2911 -23955 2955
rect -23863 2911 -23855 2955
rect -23363 2911 -23355 2955
rect -23263 2911 -23255 2955
rect -23163 2911 -23155 2955
rect -23063 2911 -23055 2955
rect -22963 2911 -22955 2955
rect -22863 2911 -22855 2955
rect -22763 2911 -22755 2955
rect -22663 2911 -22655 2955
rect -22563 2911 -22555 2955
rect -22463 2911 -22455 2955
rect -22363 2911 -22355 2955
rect -22263 2911 -22255 2955
rect -22163 2911 -22155 2955
rect -22063 2911 -22055 2955
rect -21963 2911 -21955 2955
rect -21863 2911 -21855 2955
rect -21363 2911 -21355 2955
rect -21263 2911 -21255 2955
rect -21163 2911 -21155 2955
rect -21063 2911 -21055 2955
rect -20963 2911 -20955 2955
rect -20863 2911 -20855 2955
rect -20763 2911 -20755 2955
rect -20663 2911 -20655 2955
rect -20563 2911 -20555 2955
rect -20463 2911 -20455 2955
rect -20363 2911 -20355 2955
rect -20263 2911 -20255 2955
rect -20163 2911 -20155 2955
rect -20063 2911 -20055 2955
rect -19963 2911 -19955 2955
rect -19863 2911 -19855 2955
rect -27407 2855 -27363 2863
rect -27307 2855 -27263 2863
rect -27207 2855 -27163 2863
rect -27107 2855 -27063 2863
rect -27007 2855 -26963 2863
rect -26907 2855 -26863 2863
rect -26807 2855 -26763 2863
rect -26707 2855 -26663 2863
rect -26607 2855 -26563 2863
rect -26507 2855 -26463 2863
rect -26407 2855 -26363 2863
rect -26307 2855 -26263 2863
rect -26207 2855 -26163 2863
rect -26107 2855 -26063 2863
rect -26007 2855 -25963 2863
rect -25907 2855 -25863 2863
rect -25407 2855 -25363 2863
rect -25307 2855 -25263 2863
rect -25207 2855 -25163 2863
rect -25107 2855 -25063 2863
rect -25007 2855 -24963 2863
rect -24907 2855 -24863 2863
rect -24807 2855 -24763 2863
rect -24707 2855 -24663 2863
rect -24607 2855 -24563 2863
rect -24507 2855 -24463 2863
rect -24407 2855 -24363 2863
rect -24307 2855 -24263 2863
rect -24207 2855 -24163 2863
rect -24107 2855 -24063 2863
rect -24007 2855 -23963 2863
rect -23907 2855 -23863 2863
rect -23407 2855 -23363 2863
rect -23307 2855 -23263 2863
rect -23207 2855 -23163 2863
rect -23107 2855 -23063 2863
rect -23007 2855 -22963 2863
rect -22907 2855 -22863 2863
rect -22807 2855 -22763 2863
rect -22707 2855 -22663 2863
rect -22607 2855 -22563 2863
rect -22507 2855 -22463 2863
rect -22407 2855 -22363 2863
rect -22307 2855 -22263 2863
rect -22207 2855 -22163 2863
rect -22107 2855 -22063 2863
rect -22007 2855 -21963 2863
rect -21907 2855 -21863 2863
rect -21407 2855 -21363 2863
rect -21307 2855 -21263 2863
rect -21207 2855 -21163 2863
rect -21107 2855 -21063 2863
rect -21007 2855 -20963 2863
rect -20907 2855 -20863 2863
rect -20807 2855 -20763 2863
rect -20707 2855 -20663 2863
rect -20607 2855 -20563 2863
rect -20507 2855 -20463 2863
rect -20407 2855 -20363 2863
rect -20307 2855 -20263 2863
rect -20207 2855 -20163 2863
rect -20107 2855 -20063 2863
rect -20007 2855 -19963 2863
rect -19907 2855 -19863 2863
rect -27363 2811 -27355 2855
rect -27263 2811 -27255 2855
rect -27163 2811 -27155 2855
rect -27063 2811 -27055 2855
rect -26963 2811 -26955 2855
rect -26863 2811 -26855 2855
rect -26763 2811 -26755 2855
rect -26663 2811 -26655 2855
rect -26563 2811 -26555 2855
rect -26463 2811 -26455 2855
rect -26363 2811 -26355 2855
rect -26263 2811 -26255 2855
rect -26163 2811 -26155 2855
rect -26063 2811 -26055 2855
rect -25963 2811 -25955 2855
rect -25863 2811 -25855 2855
rect -25363 2811 -25355 2855
rect -25263 2811 -25255 2855
rect -25163 2811 -25155 2855
rect -25063 2811 -25055 2855
rect -24963 2811 -24955 2855
rect -24863 2811 -24855 2855
rect -24763 2811 -24755 2855
rect -24663 2811 -24655 2855
rect -24563 2811 -24555 2855
rect -24463 2811 -24455 2855
rect -24363 2811 -24355 2855
rect -24263 2811 -24255 2855
rect -24163 2811 -24155 2855
rect -24063 2811 -24055 2855
rect -23963 2811 -23955 2855
rect -23863 2811 -23855 2855
rect -23363 2811 -23355 2855
rect -23263 2811 -23255 2855
rect -23163 2811 -23155 2855
rect -23063 2811 -23055 2855
rect -22963 2811 -22955 2855
rect -22863 2811 -22855 2855
rect -22763 2811 -22755 2855
rect -22663 2811 -22655 2855
rect -22563 2811 -22555 2855
rect -22463 2811 -22455 2855
rect -22363 2811 -22355 2855
rect -22263 2811 -22255 2855
rect -22163 2811 -22155 2855
rect -22063 2811 -22055 2855
rect -21963 2811 -21955 2855
rect -21863 2811 -21855 2855
rect -21363 2811 -21355 2855
rect -21263 2811 -21255 2855
rect -21163 2811 -21155 2855
rect -21063 2811 -21055 2855
rect -20963 2811 -20955 2855
rect -20863 2811 -20855 2855
rect -20763 2811 -20755 2855
rect -20663 2811 -20655 2855
rect -20563 2811 -20555 2855
rect -20463 2811 -20455 2855
rect -20363 2811 -20355 2855
rect -20263 2811 -20255 2855
rect -20163 2811 -20155 2855
rect -20063 2811 -20055 2855
rect -19963 2811 -19955 2855
rect -19863 2811 -19855 2855
rect -27407 2755 -27363 2763
rect -27307 2755 -27263 2763
rect -27207 2755 -27163 2763
rect -27107 2755 -27063 2763
rect -27007 2755 -26963 2763
rect -26907 2755 -26863 2763
rect -26807 2755 -26763 2763
rect -26707 2755 -26663 2763
rect -26607 2755 -26563 2763
rect -26507 2755 -26463 2763
rect -26407 2755 -26363 2763
rect -26307 2755 -26263 2763
rect -26207 2755 -26163 2763
rect -26107 2755 -26063 2763
rect -26007 2755 -25963 2763
rect -25907 2755 -25863 2763
rect -25407 2755 -25363 2763
rect -25307 2755 -25263 2763
rect -25207 2755 -25163 2763
rect -25107 2755 -25063 2763
rect -25007 2755 -24963 2763
rect -24907 2755 -24863 2763
rect -24807 2755 -24763 2763
rect -24707 2755 -24663 2763
rect -24607 2755 -24563 2763
rect -24507 2755 -24463 2763
rect -24407 2755 -24363 2763
rect -24307 2755 -24263 2763
rect -24207 2755 -24163 2763
rect -24107 2755 -24063 2763
rect -24007 2755 -23963 2763
rect -23907 2755 -23863 2763
rect -23407 2755 -23363 2763
rect -23307 2755 -23263 2763
rect -23207 2755 -23163 2763
rect -23107 2755 -23063 2763
rect -23007 2755 -22963 2763
rect -22907 2755 -22863 2763
rect -22807 2755 -22763 2763
rect -22707 2755 -22663 2763
rect -22607 2755 -22563 2763
rect -22507 2755 -22463 2763
rect -22407 2755 -22363 2763
rect -22307 2755 -22263 2763
rect -22207 2755 -22163 2763
rect -22107 2755 -22063 2763
rect -22007 2755 -21963 2763
rect -21907 2755 -21863 2763
rect -21407 2755 -21363 2763
rect -21307 2755 -21263 2763
rect -21207 2755 -21163 2763
rect -21107 2755 -21063 2763
rect -21007 2755 -20963 2763
rect -20907 2755 -20863 2763
rect -20807 2755 -20763 2763
rect -20707 2755 -20663 2763
rect -20607 2755 -20563 2763
rect -20507 2755 -20463 2763
rect -20407 2755 -20363 2763
rect -20307 2755 -20263 2763
rect -20207 2755 -20163 2763
rect -20107 2755 -20063 2763
rect -20007 2755 -19963 2763
rect -19907 2755 -19863 2763
rect -27363 2711 -27355 2755
rect -27263 2711 -27255 2755
rect -27163 2711 -27155 2755
rect -27063 2711 -27055 2755
rect -26963 2711 -26955 2755
rect -26863 2711 -26855 2755
rect -26763 2711 -26755 2755
rect -26663 2711 -26655 2755
rect -26563 2711 -26555 2755
rect -26463 2711 -26455 2755
rect -26363 2711 -26355 2755
rect -26263 2711 -26255 2755
rect -26163 2711 -26155 2755
rect -26063 2711 -26055 2755
rect -25963 2711 -25955 2755
rect -25863 2711 -25855 2755
rect -25363 2711 -25355 2755
rect -25263 2711 -25255 2755
rect -25163 2711 -25155 2755
rect -25063 2711 -25055 2755
rect -24963 2711 -24955 2755
rect -24863 2711 -24855 2755
rect -24763 2711 -24755 2755
rect -24663 2711 -24655 2755
rect -24563 2711 -24555 2755
rect -24463 2711 -24455 2755
rect -24363 2711 -24355 2755
rect -24263 2711 -24255 2755
rect -24163 2711 -24155 2755
rect -24063 2711 -24055 2755
rect -23963 2711 -23955 2755
rect -23863 2711 -23855 2755
rect -23363 2711 -23355 2755
rect -23263 2711 -23255 2755
rect -23163 2711 -23155 2755
rect -23063 2711 -23055 2755
rect -22963 2711 -22955 2755
rect -22863 2711 -22855 2755
rect -22763 2711 -22755 2755
rect -22663 2711 -22655 2755
rect -22563 2711 -22555 2755
rect -22463 2711 -22455 2755
rect -22363 2711 -22355 2755
rect -22263 2711 -22255 2755
rect -22163 2711 -22155 2755
rect -22063 2711 -22055 2755
rect -21963 2711 -21955 2755
rect -21863 2711 -21855 2755
rect -21363 2711 -21355 2755
rect -21263 2711 -21255 2755
rect -21163 2711 -21155 2755
rect -21063 2711 -21055 2755
rect -20963 2711 -20955 2755
rect -20863 2711 -20855 2755
rect -20763 2711 -20755 2755
rect -20663 2711 -20655 2755
rect -20563 2711 -20555 2755
rect -20463 2711 -20455 2755
rect -20363 2711 -20355 2755
rect -20263 2711 -20255 2755
rect -20163 2711 -20155 2755
rect -20063 2711 -20055 2755
rect -19963 2711 -19955 2755
rect -19863 2711 -19855 2755
rect -27407 2655 -27363 2663
rect -27307 2655 -27263 2663
rect -27207 2655 -27163 2663
rect -27107 2655 -27063 2663
rect -27007 2655 -26963 2663
rect -26907 2655 -26863 2663
rect -26807 2655 -26763 2663
rect -26707 2655 -26663 2663
rect -26607 2655 -26563 2663
rect -26507 2655 -26463 2663
rect -26407 2655 -26363 2663
rect -26307 2655 -26263 2663
rect -26207 2655 -26163 2663
rect -26107 2655 -26063 2663
rect -26007 2655 -25963 2663
rect -25907 2655 -25863 2663
rect -25407 2655 -25363 2663
rect -25307 2655 -25263 2663
rect -25207 2655 -25163 2663
rect -25107 2655 -25063 2663
rect -25007 2655 -24963 2663
rect -24907 2655 -24863 2663
rect -24807 2655 -24763 2663
rect -24707 2655 -24663 2663
rect -24607 2655 -24563 2663
rect -24507 2655 -24463 2663
rect -24407 2655 -24363 2663
rect -24307 2655 -24263 2663
rect -24207 2655 -24163 2663
rect -24107 2655 -24063 2663
rect -24007 2655 -23963 2663
rect -23907 2655 -23863 2663
rect -23407 2655 -23363 2663
rect -23307 2655 -23263 2663
rect -23207 2655 -23163 2663
rect -23107 2655 -23063 2663
rect -23007 2655 -22963 2663
rect -22907 2655 -22863 2663
rect -22807 2655 -22763 2663
rect -22707 2655 -22663 2663
rect -22607 2655 -22563 2663
rect -22507 2655 -22463 2663
rect -22407 2655 -22363 2663
rect -22307 2655 -22263 2663
rect -22207 2655 -22163 2663
rect -22107 2655 -22063 2663
rect -22007 2655 -21963 2663
rect -21907 2655 -21863 2663
rect -21407 2655 -21363 2663
rect -21307 2655 -21263 2663
rect -21207 2655 -21163 2663
rect -21107 2655 -21063 2663
rect -21007 2655 -20963 2663
rect -20907 2655 -20863 2663
rect -20807 2655 -20763 2663
rect -20707 2655 -20663 2663
rect -20607 2655 -20563 2663
rect -20507 2655 -20463 2663
rect -20407 2655 -20363 2663
rect -20307 2655 -20263 2663
rect -20207 2655 -20163 2663
rect -20107 2655 -20063 2663
rect -20007 2655 -19963 2663
rect -19907 2655 -19863 2663
rect -27363 2611 -27355 2655
rect -27263 2611 -27255 2655
rect -27163 2611 -27155 2655
rect -27063 2611 -27055 2655
rect -26963 2611 -26955 2655
rect -26863 2611 -26855 2655
rect -26763 2611 -26755 2655
rect -26663 2611 -26655 2655
rect -26563 2611 -26555 2655
rect -26463 2611 -26455 2655
rect -26363 2611 -26355 2655
rect -26263 2611 -26255 2655
rect -26163 2611 -26155 2655
rect -26063 2611 -26055 2655
rect -25963 2611 -25955 2655
rect -25863 2611 -25855 2655
rect -25363 2611 -25355 2655
rect -25263 2611 -25255 2655
rect -25163 2611 -25155 2655
rect -25063 2611 -25055 2655
rect -24963 2611 -24955 2655
rect -24863 2611 -24855 2655
rect -24763 2611 -24755 2655
rect -24663 2611 -24655 2655
rect -24563 2611 -24555 2655
rect -24463 2611 -24455 2655
rect -24363 2611 -24355 2655
rect -24263 2611 -24255 2655
rect -24163 2611 -24155 2655
rect -24063 2611 -24055 2655
rect -23963 2611 -23955 2655
rect -23863 2611 -23855 2655
rect -23363 2611 -23355 2655
rect -23263 2611 -23255 2655
rect -23163 2611 -23155 2655
rect -23063 2611 -23055 2655
rect -22963 2611 -22955 2655
rect -22863 2611 -22855 2655
rect -22763 2611 -22755 2655
rect -22663 2611 -22655 2655
rect -22563 2611 -22555 2655
rect -22463 2611 -22455 2655
rect -22363 2611 -22355 2655
rect -22263 2611 -22255 2655
rect -22163 2611 -22155 2655
rect -22063 2611 -22055 2655
rect -21963 2611 -21955 2655
rect -21863 2611 -21855 2655
rect -21363 2611 -21355 2655
rect -21263 2611 -21255 2655
rect -21163 2611 -21155 2655
rect -21063 2611 -21055 2655
rect -20963 2611 -20955 2655
rect -20863 2611 -20855 2655
rect -20763 2611 -20755 2655
rect -20663 2611 -20655 2655
rect -20563 2611 -20555 2655
rect -20463 2611 -20455 2655
rect -20363 2611 -20355 2655
rect -20263 2611 -20255 2655
rect -20163 2611 -20155 2655
rect -20063 2611 -20055 2655
rect -19963 2611 -19955 2655
rect -19863 2611 -19855 2655
rect -27407 2555 -27363 2563
rect -27307 2555 -27263 2563
rect -27207 2555 -27163 2563
rect -27107 2555 -27063 2563
rect -27007 2555 -26963 2563
rect -26907 2555 -26863 2563
rect -26807 2555 -26763 2563
rect -26707 2555 -26663 2563
rect -26607 2555 -26563 2563
rect -26507 2555 -26463 2563
rect -26407 2555 -26363 2563
rect -26307 2555 -26263 2563
rect -26207 2555 -26163 2563
rect -26107 2555 -26063 2563
rect -26007 2555 -25963 2563
rect -25907 2555 -25863 2563
rect -25407 2555 -25363 2563
rect -25307 2555 -25263 2563
rect -25207 2555 -25163 2563
rect -25107 2555 -25063 2563
rect -25007 2555 -24963 2563
rect -24907 2555 -24863 2563
rect -24807 2555 -24763 2563
rect -24707 2555 -24663 2563
rect -24607 2555 -24563 2563
rect -24507 2555 -24463 2563
rect -24407 2555 -24363 2563
rect -24307 2555 -24263 2563
rect -24207 2555 -24163 2563
rect -24107 2555 -24063 2563
rect -24007 2555 -23963 2563
rect -23907 2555 -23863 2563
rect -23407 2555 -23363 2563
rect -23307 2555 -23263 2563
rect -23207 2555 -23163 2563
rect -23107 2555 -23063 2563
rect -23007 2555 -22963 2563
rect -22907 2555 -22863 2563
rect -22807 2555 -22763 2563
rect -22707 2555 -22663 2563
rect -22607 2555 -22563 2563
rect -22507 2555 -22463 2563
rect -22407 2555 -22363 2563
rect -22307 2555 -22263 2563
rect -22207 2555 -22163 2563
rect -22107 2555 -22063 2563
rect -22007 2555 -21963 2563
rect -21907 2555 -21863 2563
rect -21407 2555 -21363 2563
rect -21307 2555 -21263 2563
rect -21207 2555 -21163 2563
rect -21107 2555 -21063 2563
rect -21007 2555 -20963 2563
rect -20907 2555 -20863 2563
rect -20807 2555 -20763 2563
rect -20707 2555 -20663 2563
rect -20607 2555 -20563 2563
rect -20507 2555 -20463 2563
rect -20407 2555 -20363 2563
rect -20307 2555 -20263 2563
rect -20207 2555 -20163 2563
rect -20107 2555 -20063 2563
rect -20007 2555 -19963 2563
rect -19907 2555 -19863 2563
rect -27363 2511 -27355 2555
rect -27263 2511 -27255 2555
rect -27163 2511 -27155 2555
rect -27063 2511 -27055 2555
rect -26963 2511 -26955 2555
rect -26863 2511 -26855 2555
rect -26763 2511 -26755 2555
rect -26663 2511 -26655 2555
rect -26563 2511 -26555 2555
rect -26463 2511 -26455 2555
rect -26363 2511 -26355 2555
rect -26263 2511 -26255 2555
rect -26163 2511 -26155 2555
rect -26063 2511 -26055 2555
rect -25963 2511 -25955 2555
rect -25863 2511 -25855 2555
rect -25363 2511 -25355 2555
rect -25263 2511 -25255 2555
rect -25163 2511 -25155 2555
rect -25063 2511 -25055 2555
rect -24963 2511 -24955 2555
rect -24863 2511 -24855 2555
rect -24763 2511 -24755 2555
rect -24663 2511 -24655 2555
rect -24563 2511 -24555 2555
rect -24463 2511 -24455 2555
rect -24363 2511 -24355 2555
rect -24263 2511 -24255 2555
rect -24163 2511 -24155 2555
rect -24063 2511 -24055 2555
rect -23963 2511 -23955 2555
rect -23863 2511 -23855 2555
rect -23363 2511 -23355 2555
rect -23263 2511 -23255 2555
rect -23163 2511 -23155 2555
rect -23063 2511 -23055 2555
rect -22963 2511 -22955 2555
rect -22863 2511 -22855 2555
rect -22763 2511 -22755 2555
rect -22663 2511 -22655 2555
rect -22563 2511 -22555 2555
rect -22463 2511 -22455 2555
rect -22363 2511 -22355 2555
rect -22263 2511 -22255 2555
rect -22163 2511 -22155 2555
rect -22063 2511 -22055 2555
rect -21963 2511 -21955 2555
rect -21863 2511 -21855 2555
rect -21363 2511 -21355 2555
rect -21263 2511 -21255 2555
rect -21163 2511 -21155 2555
rect -21063 2511 -21055 2555
rect -20963 2511 -20955 2555
rect -20863 2511 -20855 2555
rect -20763 2511 -20755 2555
rect -20663 2511 -20655 2555
rect -20563 2511 -20555 2555
rect -20463 2511 -20455 2555
rect -20363 2511 -20355 2555
rect -20263 2511 -20255 2555
rect -20163 2511 -20155 2555
rect -20063 2511 -20055 2555
rect -19963 2511 -19955 2555
rect -19863 2511 -19855 2555
rect -27407 2455 -27363 2463
rect -27307 2455 -27263 2463
rect -27207 2455 -27163 2463
rect -27107 2455 -27063 2463
rect -27007 2455 -26963 2463
rect -26907 2455 -26863 2463
rect -26807 2455 -26763 2463
rect -26707 2455 -26663 2463
rect -26607 2455 -26563 2463
rect -26507 2455 -26463 2463
rect -26407 2455 -26363 2463
rect -26307 2455 -26263 2463
rect -26207 2455 -26163 2463
rect -26107 2455 -26063 2463
rect -26007 2455 -25963 2463
rect -25907 2455 -25863 2463
rect -25407 2455 -25363 2463
rect -25307 2455 -25263 2463
rect -25207 2455 -25163 2463
rect -25107 2455 -25063 2463
rect -25007 2455 -24963 2463
rect -24907 2455 -24863 2463
rect -24807 2455 -24763 2463
rect -24707 2455 -24663 2463
rect -24607 2455 -24563 2463
rect -24507 2455 -24463 2463
rect -24407 2455 -24363 2463
rect -24307 2455 -24263 2463
rect -24207 2455 -24163 2463
rect -24107 2455 -24063 2463
rect -24007 2455 -23963 2463
rect -23907 2455 -23863 2463
rect -23407 2455 -23363 2463
rect -23307 2455 -23263 2463
rect -23207 2455 -23163 2463
rect -23107 2455 -23063 2463
rect -23007 2455 -22963 2463
rect -22907 2455 -22863 2463
rect -22807 2455 -22763 2463
rect -22707 2455 -22663 2463
rect -22607 2455 -22563 2463
rect -22507 2455 -22463 2463
rect -22407 2455 -22363 2463
rect -22307 2455 -22263 2463
rect -22207 2455 -22163 2463
rect -22107 2455 -22063 2463
rect -22007 2455 -21963 2463
rect -21907 2455 -21863 2463
rect -21407 2455 -21363 2463
rect -21307 2455 -21263 2463
rect -21207 2455 -21163 2463
rect -21107 2455 -21063 2463
rect -21007 2455 -20963 2463
rect -20907 2455 -20863 2463
rect -20807 2455 -20763 2463
rect -20707 2455 -20663 2463
rect -20607 2455 -20563 2463
rect -20507 2455 -20463 2463
rect -20407 2455 -20363 2463
rect -20307 2455 -20263 2463
rect -20207 2455 -20163 2463
rect -20107 2455 -20063 2463
rect -20007 2455 -19963 2463
rect -19907 2455 -19863 2463
rect -27363 2411 -27355 2455
rect -27263 2411 -27255 2455
rect -27163 2411 -27155 2455
rect -27063 2411 -27055 2455
rect -26963 2411 -26955 2455
rect -26863 2411 -26855 2455
rect -26763 2411 -26755 2455
rect -26663 2411 -26655 2455
rect -26563 2411 -26555 2455
rect -26463 2411 -26455 2455
rect -26363 2411 -26355 2455
rect -26263 2411 -26255 2455
rect -26163 2411 -26155 2455
rect -26063 2411 -26055 2455
rect -25963 2411 -25955 2455
rect -25863 2411 -25855 2455
rect -25363 2411 -25355 2455
rect -25263 2411 -25255 2455
rect -25163 2411 -25155 2455
rect -25063 2411 -25055 2455
rect -24963 2411 -24955 2455
rect -24863 2411 -24855 2455
rect -24763 2411 -24755 2455
rect -24663 2411 -24655 2455
rect -24563 2411 -24555 2455
rect -24463 2411 -24455 2455
rect -24363 2411 -24355 2455
rect -24263 2411 -24255 2455
rect -24163 2411 -24155 2455
rect -24063 2411 -24055 2455
rect -23963 2411 -23955 2455
rect -23863 2411 -23855 2455
rect -23363 2411 -23355 2455
rect -23263 2411 -23255 2455
rect -23163 2411 -23155 2455
rect -23063 2411 -23055 2455
rect -22963 2411 -22955 2455
rect -22863 2411 -22855 2455
rect -22763 2411 -22755 2455
rect -22663 2411 -22655 2455
rect -22563 2411 -22555 2455
rect -22463 2411 -22455 2455
rect -22363 2411 -22355 2455
rect -22263 2411 -22255 2455
rect -22163 2411 -22155 2455
rect -22063 2411 -22055 2455
rect -21963 2411 -21955 2455
rect -21863 2411 -21855 2455
rect -21363 2411 -21355 2455
rect -21263 2411 -21255 2455
rect -21163 2411 -21155 2455
rect -21063 2411 -21055 2455
rect -20963 2411 -20955 2455
rect -20863 2411 -20855 2455
rect -20763 2411 -20755 2455
rect -20663 2411 -20655 2455
rect -20563 2411 -20555 2455
rect -20463 2411 -20455 2455
rect -20363 2411 -20355 2455
rect -20263 2411 -20255 2455
rect -20163 2411 -20155 2455
rect -20063 2411 -20055 2455
rect -19963 2411 -19955 2455
rect -19863 2411 -19855 2455
rect -27407 2355 -27363 2363
rect -27307 2355 -27263 2363
rect -27207 2355 -27163 2363
rect -27107 2355 -27063 2363
rect -27007 2355 -26963 2363
rect -26907 2355 -26863 2363
rect -26807 2355 -26763 2363
rect -26707 2355 -26663 2363
rect -26607 2355 -26563 2363
rect -26507 2355 -26463 2363
rect -26407 2355 -26363 2363
rect -26307 2355 -26263 2363
rect -26207 2355 -26163 2363
rect -26107 2355 -26063 2363
rect -26007 2355 -25963 2363
rect -25907 2355 -25863 2363
rect -25407 2355 -25363 2363
rect -25307 2355 -25263 2363
rect -25207 2355 -25163 2363
rect -25107 2355 -25063 2363
rect -25007 2355 -24963 2363
rect -24907 2355 -24863 2363
rect -24807 2355 -24763 2363
rect -24707 2355 -24663 2363
rect -24607 2355 -24563 2363
rect -24507 2355 -24463 2363
rect -24407 2355 -24363 2363
rect -24307 2355 -24263 2363
rect -24207 2355 -24163 2363
rect -24107 2355 -24063 2363
rect -24007 2355 -23963 2363
rect -23907 2355 -23863 2363
rect -23407 2355 -23363 2363
rect -23307 2355 -23263 2363
rect -23207 2355 -23163 2363
rect -23107 2355 -23063 2363
rect -23007 2355 -22963 2363
rect -22907 2355 -22863 2363
rect -22807 2355 -22763 2363
rect -22707 2355 -22663 2363
rect -22607 2355 -22563 2363
rect -22507 2355 -22463 2363
rect -22407 2355 -22363 2363
rect -22307 2355 -22263 2363
rect -22207 2355 -22163 2363
rect -22107 2355 -22063 2363
rect -22007 2355 -21963 2363
rect -21907 2355 -21863 2363
rect -21407 2355 -21363 2363
rect -21307 2355 -21263 2363
rect -21207 2355 -21163 2363
rect -21107 2355 -21063 2363
rect -21007 2355 -20963 2363
rect -20907 2355 -20863 2363
rect -20807 2355 -20763 2363
rect -20707 2355 -20663 2363
rect -20607 2355 -20563 2363
rect -20507 2355 -20463 2363
rect -20407 2355 -20363 2363
rect -20307 2355 -20263 2363
rect -20207 2355 -20163 2363
rect -20107 2355 -20063 2363
rect -20007 2355 -19963 2363
rect -19907 2355 -19863 2363
rect -27363 2311 -27355 2355
rect -27263 2311 -27255 2355
rect -27163 2311 -27155 2355
rect -27063 2311 -27055 2355
rect -26963 2311 -26955 2355
rect -26863 2311 -26855 2355
rect -26763 2311 -26755 2355
rect -26663 2311 -26655 2355
rect -26563 2311 -26555 2355
rect -26463 2311 -26455 2355
rect -26363 2311 -26355 2355
rect -26263 2311 -26255 2355
rect -26163 2311 -26155 2355
rect -26063 2311 -26055 2355
rect -25963 2311 -25955 2355
rect -25863 2311 -25855 2355
rect -25363 2311 -25355 2355
rect -25263 2311 -25255 2355
rect -25163 2311 -25155 2355
rect -25063 2311 -25055 2355
rect -24963 2311 -24955 2355
rect -24863 2311 -24855 2355
rect -24763 2311 -24755 2355
rect -24663 2311 -24655 2355
rect -24563 2311 -24555 2355
rect -24463 2311 -24455 2355
rect -24363 2311 -24355 2355
rect -24263 2311 -24255 2355
rect -24163 2311 -24155 2355
rect -24063 2311 -24055 2355
rect -23963 2311 -23955 2355
rect -23863 2311 -23855 2355
rect -23363 2311 -23355 2355
rect -23263 2311 -23255 2355
rect -23163 2311 -23155 2355
rect -23063 2311 -23055 2355
rect -22963 2311 -22955 2355
rect -22863 2311 -22855 2355
rect -22763 2311 -22755 2355
rect -22663 2311 -22655 2355
rect -22563 2311 -22555 2355
rect -22463 2311 -22455 2355
rect -22363 2311 -22355 2355
rect -22263 2311 -22255 2355
rect -22163 2311 -22155 2355
rect -22063 2311 -22055 2355
rect -21963 2311 -21955 2355
rect -21863 2311 -21855 2355
rect -21363 2311 -21355 2355
rect -21263 2311 -21255 2355
rect -21163 2311 -21155 2355
rect -21063 2311 -21055 2355
rect -20963 2311 -20955 2355
rect -20863 2311 -20855 2355
rect -20763 2311 -20755 2355
rect -20663 2311 -20655 2355
rect -20563 2311 -20555 2355
rect -20463 2311 -20455 2355
rect -20363 2311 -20355 2355
rect -20263 2311 -20255 2355
rect -20163 2311 -20155 2355
rect -20063 2311 -20055 2355
rect -19963 2311 -19955 2355
rect -19863 2311 -19855 2355
rect -27407 2255 -27363 2263
rect -27307 2255 -27263 2263
rect -27207 2255 -27163 2263
rect -27107 2255 -27063 2263
rect -27007 2255 -26963 2263
rect -26907 2255 -26863 2263
rect -26807 2255 -26763 2263
rect -26707 2255 -26663 2263
rect -26607 2255 -26563 2263
rect -26507 2255 -26463 2263
rect -26407 2255 -26363 2263
rect -26307 2255 -26263 2263
rect -26207 2255 -26163 2263
rect -26107 2255 -26063 2263
rect -26007 2255 -25963 2263
rect -25907 2255 -25863 2263
rect -25407 2255 -25363 2263
rect -25307 2255 -25263 2263
rect -25207 2255 -25163 2263
rect -25107 2255 -25063 2263
rect -25007 2255 -24963 2263
rect -24907 2255 -24863 2263
rect -24807 2255 -24763 2263
rect -24707 2255 -24663 2263
rect -24607 2255 -24563 2263
rect -24507 2255 -24463 2263
rect -24407 2255 -24363 2263
rect -24307 2255 -24263 2263
rect -24207 2255 -24163 2263
rect -24107 2255 -24063 2263
rect -24007 2255 -23963 2263
rect -23907 2255 -23863 2263
rect -23407 2255 -23363 2263
rect -23307 2255 -23263 2263
rect -23207 2255 -23163 2263
rect -23107 2255 -23063 2263
rect -23007 2255 -22963 2263
rect -22907 2255 -22863 2263
rect -22807 2255 -22763 2263
rect -22707 2255 -22663 2263
rect -22607 2255 -22563 2263
rect -22507 2255 -22463 2263
rect -22407 2255 -22363 2263
rect -22307 2255 -22263 2263
rect -22207 2255 -22163 2263
rect -22107 2255 -22063 2263
rect -22007 2255 -21963 2263
rect -21907 2255 -21863 2263
rect -21407 2255 -21363 2263
rect -21307 2255 -21263 2263
rect -21207 2255 -21163 2263
rect -21107 2255 -21063 2263
rect -21007 2255 -20963 2263
rect -20907 2255 -20863 2263
rect -20807 2255 -20763 2263
rect -20707 2255 -20663 2263
rect -20607 2255 -20563 2263
rect -20507 2255 -20463 2263
rect -20407 2255 -20363 2263
rect -20307 2255 -20263 2263
rect -20207 2255 -20163 2263
rect -20107 2255 -20063 2263
rect -20007 2255 -19963 2263
rect -19907 2255 -19863 2263
rect -27363 2211 -27355 2255
rect -27263 2211 -27255 2255
rect -27163 2211 -27155 2255
rect -27063 2211 -27055 2255
rect -26963 2211 -26955 2255
rect -26863 2211 -26855 2255
rect -26763 2211 -26755 2255
rect -26663 2211 -26655 2255
rect -26563 2211 -26555 2255
rect -26463 2211 -26455 2255
rect -26363 2211 -26355 2255
rect -26263 2211 -26255 2255
rect -26163 2211 -26155 2255
rect -26063 2211 -26055 2255
rect -25963 2211 -25955 2255
rect -25863 2211 -25855 2255
rect -25363 2211 -25355 2255
rect -25263 2211 -25255 2255
rect -25163 2211 -25155 2255
rect -25063 2211 -25055 2255
rect -24963 2211 -24955 2255
rect -24863 2211 -24855 2255
rect -24763 2211 -24755 2255
rect -24663 2211 -24655 2255
rect -24563 2211 -24555 2255
rect -24463 2211 -24455 2255
rect -24363 2211 -24355 2255
rect -24263 2211 -24255 2255
rect -24163 2211 -24155 2255
rect -24063 2211 -24055 2255
rect -23963 2211 -23955 2255
rect -23863 2211 -23855 2255
rect -23363 2211 -23355 2255
rect -23263 2211 -23255 2255
rect -23163 2211 -23155 2255
rect -23063 2211 -23055 2255
rect -22963 2211 -22955 2255
rect -22863 2211 -22855 2255
rect -22763 2211 -22755 2255
rect -22663 2211 -22655 2255
rect -22563 2211 -22555 2255
rect -22463 2211 -22455 2255
rect -22363 2211 -22355 2255
rect -22263 2211 -22255 2255
rect -22163 2211 -22155 2255
rect -22063 2211 -22055 2255
rect -21963 2211 -21955 2255
rect -21863 2211 -21855 2255
rect -21363 2211 -21355 2255
rect -21263 2211 -21255 2255
rect -21163 2211 -21155 2255
rect -21063 2211 -21055 2255
rect -20963 2211 -20955 2255
rect -20863 2211 -20855 2255
rect -20763 2211 -20755 2255
rect -20663 2211 -20655 2255
rect -20563 2211 -20555 2255
rect -20463 2211 -20455 2255
rect -20363 2211 -20355 2255
rect -20263 2211 -20255 2255
rect -20163 2211 -20155 2255
rect -20063 2211 -20055 2255
rect -19963 2211 -19955 2255
rect -19863 2211 -19855 2255
rect -27407 2155 -27363 2163
rect -27307 2155 -27263 2163
rect -27207 2155 -27163 2163
rect -27107 2155 -27063 2163
rect -27007 2155 -26963 2163
rect -26907 2155 -26863 2163
rect -26807 2155 -26763 2163
rect -26707 2155 -26663 2163
rect -26607 2155 -26563 2163
rect -26507 2155 -26463 2163
rect -26407 2155 -26363 2163
rect -26307 2155 -26263 2163
rect -26207 2155 -26163 2163
rect -26107 2155 -26063 2163
rect -26007 2155 -25963 2163
rect -25907 2155 -25863 2163
rect -25407 2155 -25363 2163
rect -25307 2155 -25263 2163
rect -25207 2155 -25163 2163
rect -25107 2155 -25063 2163
rect -25007 2155 -24963 2163
rect -24907 2155 -24863 2163
rect -24807 2155 -24763 2163
rect -24707 2155 -24663 2163
rect -24607 2155 -24563 2163
rect -24507 2155 -24463 2163
rect -24407 2155 -24363 2163
rect -24307 2155 -24263 2163
rect -24207 2155 -24163 2163
rect -24107 2155 -24063 2163
rect -24007 2155 -23963 2163
rect -23907 2155 -23863 2163
rect -23407 2155 -23363 2163
rect -23307 2155 -23263 2163
rect -23207 2155 -23163 2163
rect -23107 2155 -23063 2163
rect -23007 2155 -22963 2163
rect -22907 2155 -22863 2163
rect -22807 2155 -22763 2163
rect -22707 2155 -22663 2163
rect -22607 2155 -22563 2163
rect -22507 2155 -22463 2163
rect -22407 2155 -22363 2163
rect -22307 2155 -22263 2163
rect -22207 2155 -22163 2163
rect -22107 2155 -22063 2163
rect -22007 2155 -21963 2163
rect -21907 2155 -21863 2163
rect -21407 2155 -21363 2163
rect -21307 2155 -21263 2163
rect -21207 2155 -21163 2163
rect -21107 2155 -21063 2163
rect -21007 2155 -20963 2163
rect -20907 2155 -20863 2163
rect -20807 2155 -20763 2163
rect -20707 2155 -20663 2163
rect -20607 2155 -20563 2163
rect -20507 2155 -20463 2163
rect -20407 2155 -20363 2163
rect -20307 2155 -20263 2163
rect -20207 2155 -20163 2163
rect -20107 2155 -20063 2163
rect -20007 2155 -19963 2163
rect -19907 2155 -19863 2163
rect -27363 2111 -27355 2155
rect -27263 2111 -27255 2155
rect -27163 2111 -27155 2155
rect -27063 2111 -27055 2155
rect -26963 2111 -26955 2155
rect -26863 2111 -26855 2155
rect -26763 2111 -26755 2155
rect -26663 2111 -26655 2155
rect -26563 2111 -26555 2155
rect -26463 2111 -26455 2155
rect -26363 2111 -26355 2155
rect -26263 2111 -26255 2155
rect -26163 2111 -26155 2155
rect -26063 2111 -26055 2155
rect -25963 2111 -25955 2155
rect -25863 2111 -25855 2155
rect -25363 2111 -25355 2155
rect -25263 2111 -25255 2155
rect -25163 2111 -25155 2155
rect -25063 2111 -25055 2155
rect -24963 2111 -24955 2155
rect -24863 2111 -24855 2155
rect -24763 2111 -24755 2155
rect -24663 2111 -24655 2155
rect -24563 2111 -24555 2155
rect -24463 2111 -24455 2155
rect -24363 2111 -24355 2155
rect -24263 2111 -24255 2155
rect -24163 2111 -24155 2155
rect -24063 2111 -24055 2155
rect -23963 2111 -23955 2155
rect -23863 2111 -23855 2155
rect -23363 2111 -23355 2155
rect -23263 2111 -23255 2155
rect -23163 2111 -23155 2155
rect -23063 2111 -23055 2155
rect -22963 2111 -22955 2155
rect -22863 2111 -22855 2155
rect -22763 2111 -22755 2155
rect -22663 2111 -22655 2155
rect -22563 2111 -22555 2155
rect -22463 2111 -22455 2155
rect -22363 2111 -22355 2155
rect -22263 2111 -22255 2155
rect -22163 2111 -22155 2155
rect -22063 2111 -22055 2155
rect -21963 2111 -21955 2155
rect -21863 2111 -21855 2155
rect -21363 2111 -21355 2155
rect -21263 2111 -21255 2155
rect -21163 2111 -21155 2155
rect -21063 2111 -21055 2155
rect -20963 2111 -20955 2155
rect -20863 2111 -20855 2155
rect -20763 2111 -20755 2155
rect -20663 2111 -20655 2155
rect -20563 2111 -20555 2155
rect -20463 2111 -20455 2155
rect -20363 2111 -20355 2155
rect -20263 2111 -20255 2155
rect -20163 2111 -20155 2155
rect -20063 2111 -20055 2155
rect -19963 2111 -19955 2155
rect -19863 2111 -19855 2155
rect -27407 2055 -27363 2063
rect -27307 2055 -27263 2063
rect -27207 2055 -27163 2063
rect -27107 2055 -27063 2063
rect -27007 2055 -26963 2063
rect -26907 2055 -26863 2063
rect -26807 2055 -26763 2063
rect -26707 2055 -26663 2063
rect -26607 2055 -26563 2063
rect -26507 2055 -26463 2063
rect -26407 2055 -26363 2063
rect -26307 2055 -26263 2063
rect -26207 2055 -26163 2063
rect -26107 2055 -26063 2063
rect -26007 2055 -25963 2063
rect -25907 2055 -25863 2063
rect -25407 2055 -25363 2063
rect -25307 2055 -25263 2063
rect -25207 2055 -25163 2063
rect -25107 2055 -25063 2063
rect -25007 2055 -24963 2063
rect -24907 2055 -24863 2063
rect -24807 2055 -24763 2063
rect -24707 2055 -24663 2063
rect -24607 2055 -24563 2063
rect -24507 2055 -24463 2063
rect -24407 2055 -24363 2063
rect -24307 2055 -24263 2063
rect -24207 2055 -24163 2063
rect -24107 2055 -24063 2063
rect -24007 2055 -23963 2063
rect -23907 2055 -23863 2063
rect -23407 2055 -23363 2063
rect -23307 2055 -23263 2063
rect -23207 2055 -23163 2063
rect -23107 2055 -23063 2063
rect -23007 2055 -22963 2063
rect -22907 2055 -22863 2063
rect -22807 2055 -22763 2063
rect -22707 2055 -22663 2063
rect -22607 2055 -22563 2063
rect -22507 2055 -22463 2063
rect -22407 2055 -22363 2063
rect -22307 2055 -22263 2063
rect -22207 2055 -22163 2063
rect -22107 2055 -22063 2063
rect -22007 2055 -21963 2063
rect -21907 2055 -21863 2063
rect -21407 2055 -21363 2063
rect -21307 2055 -21263 2063
rect -21207 2055 -21163 2063
rect -21107 2055 -21063 2063
rect -21007 2055 -20963 2063
rect -20907 2055 -20863 2063
rect -20807 2055 -20763 2063
rect -20707 2055 -20663 2063
rect -20607 2055 -20563 2063
rect -20507 2055 -20463 2063
rect -20407 2055 -20363 2063
rect -20307 2055 -20263 2063
rect -20207 2055 -20163 2063
rect -20107 2055 -20063 2063
rect -20007 2055 -19963 2063
rect -19907 2055 -19863 2063
rect -27363 2011 -27355 2055
rect -27263 2011 -27255 2055
rect -27163 2011 -27155 2055
rect -27063 2011 -27055 2055
rect -26963 2011 -26955 2055
rect -26863 2011 -26855 2055
rect -26763 2011 -26755 2055
rect -26663 2011 -26655 2055
rect -26563 2011 -26555 2055
rect -26463 2011 -26455 2055
rect -26363 2011 -26355 2055
rect -26263 2011 -26255 2055
rect -26163 2011 -26155 2055
rect -26063 2011 -26055 2055
rect -25963 2011 -25955 2055
rect -25863 2011 -25855 2055
rect -25363 2011 -25355 2055
rect -25263 2011 -25255 2055
rect -25163 2011 -25155 2055
rect -25063 2011 -25055 2055
rect -24963 2011 -24955 2055
rect -24863 2011 -24855 2055
rect -24763 2011 -24755 2055
rect -24663 2011 -24655 2055
rect -24563 2011 -24555 2055
rect -24463 2011 -24455 2055
rect -24363 2011 -24355 2055
rect -24263 2011 -24255 2055
rect -24163 2011 -24155 2055
rect -24063 2011 -24055 2055
rect -23963 2011 -23955 2055
rect -23863 2011 -23855 2055
rect -23363 2011 -23355 2055
rect -23263 2011 -23255 2055
rect -23163 2011 -23155 2055
rect -23063 2011 -23055 2055
rect -22963 2011 -22955 2055
rect -22863 2011 -22855 2055
rect -22763 2011 -22755 2055
rect -22663 2011 -22655 2055
rect -22563 2011 -22555 2055
rect -22463 2011 -22455 2055
rect -22363 2011 -22355 2055
rect -22263 2011 -22255 2055
rect -22163 2011 -22155 2055
rect -22063 2011 -22055 2055
rect -21963 2011 -21955 2055
rect -21863 2011 -21855 2055
rect -21363 2011 -21355 2055
rect -21263 2011 -21255 2055
rect -21163 2011 -21155 2055
rect -21063 2011 -21055 2055
rect -20963 2011 -20955 2055
rect -20863 2011 -20855 2055
rect -20763 2011 -20755 2055
rect -20663 2011 -20655 2055
rect -20563 2011 -20555 2055
rect -20463 2011 -20455 2055
rect -20363 2011 -20355 2055
rect -20263 2011 -20255 2055
rect -20163 2011 -20155 2055
rect -20063 2011 -20055 2055
rect -19963 2011 -19955 2055
rect -19863 2011 -19855 2055
rect 144904 -17445 144948 -17437
rect 145004 -17445 145048 -17437
rect 145104 -17445 145148 -17437
rect 145204 -17445 145248 -17437
rect 145304 -17445 145348 -17437
rect 145404 -17445 145448 -17437
rect 145504 -17445 145548 -17437
rect 145604 -17445 145648 -17437
rect 145704 -17445 145748 -17437
rect 145804 -17445 145848 -17437
rect 145904 -17445 145948 -17437
rect 146004 -17445 146048 -17437
rect 146104 -17445 146148 -17437
rect 146204 -17445 146248 -17437
rect 146304 -17445 146348 -17437
rect 146404 -17445 146448 -17437
rect 146904 -17445 146948 -17437
rect 147004 -17445 147048 -17437
rect 147104 -17445 147148 -17437
rect 147204 -17445 147248 -17437
rect 147304 -17445 147348 -17437
rect 147404 -17445 147448 -17437
rect 147504 -17445 147548 -17437
rect 147604 -17445 147648 -17437
rect 147704 -17445 147748 -17437
rect 147804 -17445 147848 -17437
rect 147904 -17445 147948 -17437
rect 148004 -17445 148048 -17437
rect 148104 -17445 148148 -17437
rect 148204 -17445 148248 -17437
rect 148304 -17445 148348 -17437
rect 148404 -17445 148448 -17437
rect 148904 -17445 148948 -17437
rect 149004 -17445 149048 -17437
rect 149104 -17445 149148 -17437
rect 149204 -17445 149248 -17437
rect 149304 -17445 149348 -17437
rect 149404 -17445 149448 -17437
rect 149504 -17445 149548 -17437
rect 149604 -17445 149648 -17437
rect 149704 -17445 149748 -17437
rect 149804 -17445 149848 -17437
rect 149904 -17445 149948 -17437
rect 150004 -17445 150048 -17437
rect 150104 -17445 150148 -17437
rect 150204 -17445 150248 -17437
rect 150304 -17445 150348 -17437
rect 150404 -17445 150448 -17437
rect 150904 -17445 150948 -17437
rect 151004 -17445 151048 -17437
rect 151104 -17445 151148 -17437
rect 151204 -17445 151248 -17437
rect 151304 -17445 151348 -17437
rect 151404 -17445 151448 -17437
rect 151504 -17445 151548 -17437
rect 151604 -17445 151648 -17437
rect 151704 -17445 151748 -17437
rect 151804 -17445 151848 -17437
rect 151904 -17445 151948 -17437
rect 152004 -17445 152048 -17437
rect 152104 -17445 152148 -17437
rect 152204 -17445 152248 -17437
rect 152304 -17445 152348 -17437
rect 152404 -17445 152448 -17437
rect 144948 -17489 144956 -17445
rect 145048 -17489 145056 -17445
rect 145148 -17489 145156 -17445
rect 145248 -17489 145256 -17445
rect 145348 -17489 145356 -17445
rect 145448 -17489 145456 -17445
rect 145548 -17489 145556 -17445
rect 145648 -17489 145656 -17445
rect 145748 -17489 145756 -17445
rect 145848 -17489 145856 -17445
rect 145948 -17489 145956 -17445
rect 146048 -17489 146056 -17445
rect 146148 -17489 146156 -17445
rect 146248 -17489 146256 -17445
rect 146348 -17489 146356 -17445
rect 146448 -17489 146456 -17445
rect 146948 -17489 146956 -17445
rect 147048 -17489 147056 -17445
rect 147148 -17489 147156 -17445
rect 147248 -17489 147256 -17445
rect 147348 -17489 147356 -17445
rect 147448 -17489 147456 -17445
rect 147548 -17489 147556 -17445
rect 147648 -17489 147656 -17445
rect 147748 -17489 147756 -17445
rect 147848 -17489 147856 -17445
rect 147948 -17489 147956 -17445
rect 148048 -17489 148056 -17445
rect 148148 -17489 148156 -17445
rect 148248 -17489 148256 -17445
rect 148348 -17489 148356 -17445
rect 148448 -17489 148456 -17445
rect 148948 -17489 148956 -17445
rect 149048 -17489 149056 -17445
rect 149148 -17489 149156 -17445
rect 149248 -17489 149256 -17445
rect 149348 -17489 149356 -17445
rect 149448 -17489 149456 -17445
rect 149548 -17489 149556 -17445
rect 149648 -17489 149656 -17445
rect 149748 -17489 149756 -17445
rect 149848 -17489 149856 -17445
rect 149948 -17489 149956 -17445
rect 150048 -17489 150056 -17445
rect 150148 -17489 150156 -17445
rect 150248 -17489 150256 -17445
rect 150348 -17489 150356 -17445
rect 150448 -17489 150456 -17445
rect 150948 -17489 150956 -17445
rect 151048 -17489 151056 -17445
rect 151148 -17489 151156 -17445
rect 151248 -17489 151256 -17445
rect 151348 -17489 151356 -17445
rect 151448 -17489 151456 -17445
rect 151548 -17489 151556 -17445
rect 151648 -17489 151656 -17445
rect 151748 -17489 151756 -17445
rect 151848 -17489 151856 -17445
rect 151948 -17489 151956 -17445
rect 152048 -17489 152056 -17445
rect 152148 -17489 152156 -17445
rect 152248 -17489 152256 -17445
rect 152348 -17489 152356 -17445
rect 152448 -17489 152456 -17445
rect 144904 -17545 144948 -17537
rect 145004 -17545 145048 -17537
rect 145104 -17545 145148 -17537
rect 145204 -17545 145248 -17537
rect 145304 -17545 145348 -17537
rect 145404 -17545 145448 -17537
rect 145504 -17545 145548 -17537
rect 145604 -17545 145648 -17537
rect 145704 -17545 145748 -17537
rect 145804 -17545 145848 -17537
rect 145904 -17545 145948 -17537
rect 146004 -17545 146048 -17537
rect 146104 -17545 146148 -17537
rect 146204 -17545 146248 -17537
rect 146304 -17545 146348 -17537
rect 146404 -17545 146448 -17537
rect 146904 -17545 146948 -17537
rect 147004 -17545 147048 -17537
rect 147104 -17545 147148 -17537
rect 147204 -17545 147248 -17537
rect 147304 -17545 147348 -17537
rect 147404 -17545 147448 -17537
rect 147504 -17545 147548 -17537
rect 147604 -17545 147648 -17537
rect 147704 -17545 147748 -17537
rect 147804 -17545 147848 -17537
rect 147904 -17545 147948 -17537
rect 148004 -17545 148048 -17537
rect 148104 -17545 148148 -17537
rect 148204 -17545 148248 -17537
rect 148304 -17545 148348 -17537
rect 148404 -17545 148448 -17537
rect 148904 -17545 148948 -17537
rect 149004 -17545 149048 -17537
rect 149104 -17545 149148 -17537
rect 149204 -17545 149248 -17537
rect 149304 -17545 149348 -17537
rect 149404 -17545 149448 -17537
rect 149504 -17545 149548 -17537
rect 149604 -17545 149648 -17537
rect 149704 -17545 149748 -17537
rect 149804 -17545 149848 -17537
rect 149904 -17545 149948 -17537
rect 150004 -17545 150048 -17537
rect 150104 -17545 150148 -17537
rect 150204 -17545 150248 -17537
rect 150304 -17545 150348 -17537
rect 150404 -17545 150448 -17537
rect 150904 -17545 150948 -17537
rect 151004 -17545 151048 -17537
rect 151104 -17545 151148 -17537
rect 151204 -17545 151248 -17537
rect 151304 -17545 151348 -17537
rect 151404 -17545 151448 -17537
rect 151504 -17545 151548 -17537
rect 151604 -17545 151648 -17537
rect 151704 -17545 151748 -17537
rect 151804 -17545 151848 -17537
rect 151904 -17545 151948 -17537
rect 152004 -17545 152048 -17537
rect 152104 -17545 152148 -17537
rect 152204 -17545 152248 -17537
rect 152304 -17545 152348 -17537
rect 152404 -17545 152448 -17537
rect 144948 -17589 144956 -17545
rect 145048 -17589 145056 -17545
rect 145148 -17589 145156 -17545
rect 145248 -17589 145256 -17545
rect 145348 -17589 145356 -17545
rect 145448 -17589 145456 -17545
rect 145548 -17589 145556 -17545
rect 145648 -17589 145656 -17545
rect 145748 -17589 145756 -17545
rect 145848 -17589 145856 -17545
rect 145948 -17589 145956 -17545
rect 146048 -17589 146056 -17545
rect 146148 -17589 146156 -17545
rect 146248 -17589 146256 -17545
rect 146348 -17589 146356 -17545
rect 146448 -17589 146456 -17545
rect 146948 -17589 146956 -17545
rect 147048 -17589 147056 -17545
rect 147148 -17589 147156 -17545
rect 147248 -17589 147256 -17545
rect 147348 -17589 147356 -17545
rect 147448 -17589 147456 -17545
rect 147548 -17589 147556 -17545
rect 147648 -17589 147656 -17545
rect 147748 -17589 147756 -17545
rect 147848 -17589 147856 -17545
rect 147948 -17589 147956 -17545
rect 148048 -17589 148056 -17545
rect 148148 -17589 148156 -17545
rect 148248 -17589 148256 -17545
rect 148348 -17589 148356 -17545
rect 148448 -17589 148456 -17545
rect 148948 -17589 148956 -17545
rect 149048 -17589 149056 -17545
rect 149148 -17589 149156 -17545
rect 149248 -17589 149256 -17545
rect 149348 -17589 149356 -17545
rect 149448 -17589 149456 -17545
rect 149548 -17589 149556 -17545
rect 149648 -17589 149656 -17545
rect 149748 -17589 149756 -17545
rect 149848 -17589 149856 -17545
rect 149948 -17589 149956 -17545
rect 150048 -17589 150056 -17545
rect 150148 -17589 150156 -17545
rect 150248 -17589 150256 -17545
rect 150348 -17589 150356 -17545
rect 150448 -17589 150456 -17545
rect 150948 -17589 150956 -17545
rect 151048 -17589 151056 -17545
rect 151148 -17589 151156 -17545
rect 151248 -17589 151256 -17545
rect 151348 -17589 151356 -17545
rect 151448 -17589 151456 -17545
rect 151548 -17589 151556 -17545
rect 151648 -17589 151656 -17545
rect 151748 -17589 151756 -17545
rect 151848 -17589 151856 -17545
rect 151948 -17589 151956 -17545
rect 152048 -17589 152056 -17545
rect 152148 -17589 152156 -17545
rect 152248 -17589 152256 -17545
rect 152348 -17589 152356 -17545
rect 152448 -17589 152456 -17545
rect 144904 -17645 144948 -17637
rect 145004 -17645 145048 -17637
rect 145104 -17645 145148 -17637
rect 145204 -17645 145248 -17637
rect 145304 -17645 145348 -17637
rect 145404 -17645 145448 -17637
rect 145504 -17645 145548 -17637
rect 145604 -17645 145648 -17637
rect 145704 -17645 145748 -17637
rect 145804 -17645 145848 -17637
rect 145904 -17645 145948 -17637
rect 146004 -17645 146048 -17637
rect 146104 -17645 146148 -17637
rect 146204 -17645 146248 -17637
rect 146304 -17645 146348 -17637
rect 146404 -17645 146448 -17637
rect 146904 -17645 146948 -17637
rect 147004 -17645 147048 -17637
rect 147104 -17645 147148 -17637
rect 147204 -17645 147248 -17637
rect 147304 -17645 147348 -17637
rect 147404 -17645 147448 -17637
rect 147504 -17645 147548 -17637
rect 147604 -17645 147648 -17637
rect 147704 -17645 147748 -17637
rect 147804 -17645 147848 -17637
rect 147904 -17645 147948 -17637
rect 148004 -17645 148048 -17637
rect 148104 -17645 148148 -17637
rect 148204 -17645 148248 -17637
rect 148304 -17645 148348 -17637
rect 148404 -17645 148448 -17637
rect 148904 -17645 148948 -17637
rect 149004 -17645 149048 -17637
rect 149104 -17645 149148 -17637
rect 149204 -17645 149248 -17637
rect 149304 -17645 149348 -17637
rect 149404 -17645 149448 -17637
rect 149504 -17645 149548 -17637
rect 149604 -17645 149648 -17637
rect 149704 -17645 149748 -17637
rect 149804 -17645 149848 -17637
rect 149904 -17645 149948 -17637
rect 150004 -17645 150048 -17637
rect 150104 -17645 150148 -17637
rect 150204 -17645 150248 -17637
rect 150304 -17645 150348 -17637
rect 150404 -17645 150448 -17637
rect 150904 -17645 150948 -17637
rect 151004 -17645 151048 -17637
rect 151104 -17645 151148 -17637
rect 151204 -17645 151248 -17637
rect 151304 -17645 151348 -17637
rect 151404 -17645 151448 -17637
rect 151504 -17645 151548 -17637
rect 151604 -17645 151648 -17637
rect 151704 -17645 151748 -17637
rect 151804 -17645 151848 -17637
rect 151904 -17645 151948 -17637
rect 152004 -17645 152048 -17637
rect 152104 -17645 152148 -17637
rect 152204 -17645 152248 -17637
rect 152304 -17645 152348 -17637
rect 152404 -17645 152448 -17637
rect 144948 -17689 144956 -17645
rect 145048 -17689 145056 -17645
rect 145148 -17689 145156 -17645
rect 145248 -17689 145256 -17645
rect 145348 -17689 145356 -17645
rect 145448 -17689 145456 -17645
rect 145548 -17689 145556 -17645
rect 145648 -17689 145656 -17645
rect 145748 -17689 145756 -17645
rect 145848 -17689 145856 -17645
rect 145948 -17689 145956 -17645
rect 146048 -17689 146056 -17645
rect 146148 -17689 146156 -17645
rect 146248 -17689 146256 -17645
rect 146348 -17689 146356 -17645
rect 146448 -17689 146456 -17645
rect 146948 -17689 146956 -17645
rect 147048 -17689 147056 -17645
rect 147148 -17689 147156 -17645
rect 147248 -17689 147256 -17645
rect 147348 -17689 147356 -17645
rect 147448 -17689 147456 -17645
rect 147548 -17689 147556 -17645
rect 147648 -17689 147656 -17645
rect 147748 -17689 147756 -17645
rect 147848 -17689 147856 -17645
rect 147948 -17689 147956 -17645
rect 148048 -17689 148056 -17645
rect 148148 -17689 148156 -17645
rect 148248 -17689 148256 -17645
rect 148348 -17689 148356 -17645
rect 148448 -17689 148456 -17645
rect 148948 -17689 148956 -17645
rect 149048 -17689 149056 -17645
rect 149148 -17689 149156 -17645
rect 149248 -17689 149256 -17645
rect 149348 -17689 149356 -17645
rect 149448 -17689 149456 -17645
rect 149548 -17689 149556 -17645
rect 149648 -17689 149656 -17645
rect 149748 -17689 149756 -17645
rect 149848 -17689 149856 -17645
rect 149948 -17689 149956 -17645
rect 150048 -17689 150056 -17645
rect 150148 -17689 150156 -17645
rect 150248 -17689 150256 -17645
rect 150348 -17689 150356 -17645
rect 150448 -17689 150456 -17645
rect 150948 -17689 150956 -17645
rect 151048 -17689 151056 -17645
rect 151148 -17689 151156 -17645
rect 151248 -17689 151256 -17645
rect 151348 -17689 151356 -17645
rect 151448 -17689 151456 -17645
rect 151548 -17689 151556 -17645
rect 151648 -17689 151656 -17645
rect 151748 -17689 151756 -17645
rect 151848 -17689 151856 -17645
rect 151948 -17689 151956 -17645
rect 152048 -17689 152056 -17645
rect 152148 -17689 152156 -17645
rect 152248 -17689 152256 -17645
rect 152348 -17689 152356 -17645
rect 152448 -17689 152456 -17645
rect 144904 -17745 144948 -17737
rect 145004 -17745 145048 -17737
rect 145104 -17745 145148 -17737
rect 145204 -17745 145248 -17737
rect 145304 -17745 145348 -17737
rect 145404 -17745 145448 -17737
rect 145504 -17745 145548 -17737
rect 145604 -17745 145648 -17737
rect 145704 -17745 145748 -17737
rect 145804 -17745 145848 -17737
rect 145904 -17745 145948 -17737
rect 146004 -17745 146048 -17737
rect 146104 -17745 146148 -17737
rect 146204 -17745 146248 -17737
rect 146304 -17745 146348 -17737
rect 146404 -17745 146448 -17737
rect 146904 -17745 146948 -17737
rect 147004 -17745 147048 -17737
rect 147104 -17745 147148 -17737
rect 147204 -17745 147248 -17737
rect 147304 -17745 147348 -17737
rect 147404 -17745 147448 -17737
rect 147504 -17745 147548 -17737
rect 147604 -17745 147648 -17737
rect 147704 -17745 147748 -17737
rect 147804 -17745 147848 -17737
rect 147904 -17745 147948 -17737
rect 148004 -17745 148048 -17737
rect 148104 -17745 148148 -17737
rect 148204 -17745 148248 -17737
rect 148304 -17745 148348 -17737
rect 148404 -17745 148448 -17737
rect 148904 -17745 148948 -17737
rect 149004 -17745 149048 -17737
rect 149104 -17745 149148 -17737
rect 149204 -17745 149248 -17737
rect 149304 -17745 149348 -17737
rect 149404 -17745 149448 -17737
rect 149504 -17745 149548 -17737
rect 149604 -17745 149648 -17737
rect 149704 -17745 149748 -17737
rect 149804 -17745 149848 -17737
rect 149904 -17745 149948 -17737
rect 150004 -17745 150048 -17737
rect 150104 -17745 150148 -17737
rect 150204 -17745 150248 -17737
rect 150304 -17745 150348 -17737
rect 150404 -17745 150448 -17737
rect 150904 -17745 150948 -17737
rect 151004 -17745 151048 -17737
rect 151104 -17745 151148 -17737
rect 151204 -17745 151248 -17737
rect 151304 -17745 151348 -17737
rect 151404 -17745 151448 -17737
rect 151504 -17745 151548 -17737
rect 151604 -17745 151648 -17737
rect 151704 -17745 151748 -17737
rect 151804 -17745 151848 -17737
rect 151904 -17745 151948 -17737
rect 152004 -17745 152048 -17737
rect 152104 -17745 152148 -17737
rect 152204 -17745 152248 -17737
rect 152304 -17745 152348 -17737
rect 152404 -17745 152448 -17737
rect 144948 -17789 144956 -17745
rect 145048 -17789 145056 -17745
rect 145148 -17789 145156 -17745
rect 145248 -17789 145256 -17745
rect 145348 -17789 145356 -17745
rect 145448 -17789 145456 -17745
rect 145548 -17789 145556 -17745
rect 145648 -17789 145656 -17745
rect 145748 -17789 145756 -17745
rect 145848 -17789 145856 -17745
rect 145948 -17789 145956 -17745
rect 146048 -17789 146056 -17745
rect 146148 -17789 146156 -17745
rect 146248 -17789 146256 -17745
rect 146348 -17789 146356 -17745
rect 146448 -17789 146456 -17745
rect 146948 -17789 146956 -17745
rect 147048 -17789 147056 -17745
rect 147148 -17789 147156 -17745
rect 147248 -17789 147256 -17745
rect 147348 -17789 147356 -17745
rect 147448 -17789 147456 -17745
rect 147548 -17789 147556 -17745
rect 147648 -17789 147656 -17745
rect 147748 -17789 147756 -17745
rect 147848 -17789 147856 -17745
rect 147948 -17789 147956 -17745
rect 148048 -17789 148056 -17745
rect 148148 -17789 148156 -17745
rect 148248 -17789 148256 -17745
rect 148348 -17789 148356 -17745
rect 148448 -17789 148456 -17745
rect 148948 -17789 148956 -17745
rect 149048 -17789 149056 -17745
rect 149148 -17789 149156 -17745
rect 149248 -17789 149256 -17745
rect 149348 -17789 149356 -17745
rect 149448 -17789 149456 -17745
rect 149548 -17789 149556 -17745
rect 149648 -17789 149656 -17745
rect 149748 -17789 149756 -17745
rect 149848 -17789 149856 -17745
rect 149948 -17789 149956 -17745
rect 150048 -17789 150056 -17745
rect 150148 -17789 150156 -17745
rect 150248 -17789 150256 -17745
rect 150348 -17789 150356 -17745
rect 150448 -17789 150456 -17745
rect 150948 -17789 150956 -17745
rect 151048 -17789 151056 -17745
rect 151148 -17789 151156 -17745
rect 151248 -17789 151256 -17745
rect 151348 -17789 151356 -17745
rect 151448 -17789 151456 -17745
rect 151548 -17789 151556 -17745
rect 151648 -17789 151656 -17745
rect 151748 -17789 151756 -17745
rect 151848 -17789 151856 -17745
rect 151948 -17789 151956 -17745
rect 152048 -17789 152056 -17745
rect 152148 -17789 152156 -17745
rect 152248 -17789 152256 -17745
rect 152348 -17789 152356 -17745
rect 152448 -17789 152456 -17745
rect 144904 -17845 144948 -17837
rect 145004 -17845 145048 -17837
rect 145104 -17845 145148 -17837
rect 145204 -17845 145248 -17837
rect 145304 -17845 145348 -17837
rect 145404 -17845 145448 -17837
rect 145504 -17845 145548 -17837
rect 145604 -17845 145648 -17837
rect 145704 -17845 145748 -17837
rect 145804 -17845 145848 -17837
rect 145904 -17845 145948 -17837
rect 146004 -17845 146048 -17837
rect 146104 -17845 146148 -17837
rect 146204 -17845 146248 -17837
rect 146304 -17845 146348 -17837
rect 146404 -17845 146448 -17837
rect 146904 -17845 146948 -17837
rect 147004 -17845 147048 -17837
rect 147104 -17845 147148 -17837
rect 147204 -17845 147248 -17837
rect 147304 -17845 147348 -17837
rect 147404 -17845 147448 -17837
rect 147504 -17845 147548 -17837
rect 147604 -17845 147648 -17837
rect 147704 -17845 147748 -17837
rect 147804 -17845 147848 -17837
rect 147904 -17845 147948 -17837
rect 148004 -17845 148048 -17837
rect 148104 -17845 148148 -17837
rect 148204 -17845 148248 -17837
rect 148304 -17845 148348 -17837
rect 148404 -17845 148448 -17837
rect 148904 -17845 148948 -17837
rect 149004 -17845 149048 -17837
rect 149104 -17845 149148 -17837
rect 149204 -17845 149248 -17837
rect 149304 -17845 149348 -17837
rect 149404 -17845 149448 -17837
rect 149504 -17845 149548 -17837
rect 149604 -17845 149648 -17837
rect 149704 -17845 149748 -17837
rect 149804 -17845 149848 -17837
rect 149904 -17845 149948 -17837
rect 150004 -17845 150048 -17837
rect 150104 -17845 150148 -17837
rect 150204 -17845 150248 -17837
rect 150304 -17845 150348 -17837
rect 150404 -17845 150448 -17837
rect 150904 -17845 150948 -17837
rect 151004 -17845 151048 -17837
rect 151104 -17845 151148 -17837
rect 151204 -17845 151248 -17837
rect 151304 -17845 151348 -17837
rect 151404 -17845 151448 -17837
rect 151504 -17845 151548 -17837
rect 151604 -17845 151648 -17837
rect 151704 -17845 151748 -17837
rect 151804 -17845 151848 -17837
rect 151904 -17845 151948 -17837
rect 152004 -17845 152048 -17837
rect 152104 -17845 152148 -17837
rect 152204 -17845 152248 -17837
rect 152304 -17845 152348 -17837
rect 152404 -17845 152448 -17837
rect 144948 -17889 144956 -17845
rect 145048 -17889 145056 -17845
rect 145148 -17889 145156 -17845
rect 145248 -17889 145256 -17845
rect 145348 -17889 145356 -17845
rect 145448 -17889 145456 -17845
rect 145548 -17889 145556 -17845
rect 145648 -17889 145656 -17845
rect 145748 -17889 145756 -17845
rect 145848 -17889 145856 -17845
rect 145948 -17889 145956 -17845
rect 146048 -17889 146056 -17845
rect 146148 -17889 146156 -17845
rect 146248 -17889 146256 -17845
rect 146348 -17889 146356 -17845
rect 146448 -17889 146456 -17845
rect 146948 -17889 146956 -17845
rect 147048 -17889 147056 -17845
rect 147148 -17889 147156 -17845
rect 147248 -17889 147256 -17845
rect 147348 -17889 147356 -17845
rect 147448 -17889 147456 -17845
rect 147548 -17889 147556 -17845
rect 147648 -17889 147656 -17845
rect 147748 -17889 147756 -17845
rect 147848 -17889 147856 -17845
rect 147948 -17889 147956 -17845
rect 148048 -17889 148056 -17845
rect 148148 -17889 148156 -17845
rect 148248 -17889 148256 -17845
rect 148348 -17889 148356 -17845
rect 148448 -17889 148456 -17845
rect 148948 -17889 148956 -17845
rect 149048 -17889 149056 -17845
rect 149148 -17889 149156 -17845
rect 149248 -17889 149256 -17845
rect 149348 -17889 149356 -17845
rect 149448 -17889 149456 -17845
rect 149548 -17889 149556 -17845
rect 149648 -17889 149656 -17845
rect 149748 -17889 149756 -17845
rect 149848 -17889 149856 -17845
rect 149948 -17889 149956 -17845
rect 150048 -17889 150056 -17845
rect 150148 -17889 150156 -17845
rect 150248 -17889 150256 -17845
rect 150348 -17889 150356 -17845
rect 150448 -17889 150456 -17845
rect 150948 -17889 150956 -17845
rect 151048 -17889 151056 -17845
rect 151148 -17889 151156 -17845
rect 151248 -17889 151256 -17845
rect 151348 -17889 151356 -17845
rect 151448 -17889 151456 -17845
rect 151548 -17889 151556 -17845
rect 151648 -17889 151656 -17845
rect 151748 -17889 151756 -17845
rect 151848 -17889 151856 -17845
rect 151948 -17889 151956 -17845
rect 152048 -17889 152056 -17845
rect 152148 -17889 152156 -17845
rect 152248 -17889 152256 -17845
rect 152348 -17889 152356 -17845
rect 152448 -17889 152456 -17845
rect 144904 -17945 144948 -17937
rect 145004 -17945 145048 -17937
rect 145104 -17945 145148 -17937
rect 145204 -17945 145248 -17937
rect 145304 -17945 145348 -17937
rect 145404 -17945 145448 -17937
rect 145504 -17945 145548 -17937
rect 145604 -17945 145648 -17937
rect 145704 -17945 145748 -17937
rect 145804 -17945 145848 -17937
rect 145904 -17945 145948 -17937
rect 146004 -17945 146048 -17937
rect 146104 -17945 146148 -17937
rect 146204 -17945 146248 -17937
rect 146304 -17945 146348 -17937
rect 146404 -17945 146448 -17937
rect 146904 -17945 146948 -17937
rect 147004 -17945 147048 -17937
rect 147104 -17945 147148 -17937
rect 147204 -17945 147248 -17937
rect 147304 -17945 147348 -17937
rect 147404 -17945 147448 -17937
rect 147504 -17945 147548 -17937
rect 147604 -17945 147648 -17937
rect 147704 -17945 147748 -17937
rect 147804 -17945 147848 -17937
rect 147904 -17945 147948 -17937
rect 148004 -17945 148048 -17937
rect 148104 -17945 148148 -17937
rect 148204 -17945 148248 -17937
rect 148304 -17945 148348 -17937
rect 148404 -17945 148448 -17937
rect 148904 -17945 148948 -17937
rect 149004 -17945 149048 -17937
rect 149104 -17945 149148 -17937
rect 149204 -17945 149248 -17937
rect 149304 -17945 149348 -17937
rect 149404 -17945 149448 -17937
rect 149504 -17945 149548 -17937
rect 149604 -17945 149648 -17937
rect 149704 -17945 149748 -17937
rect 149804 -17945 149848 -17937
rect 149904 -17945 149948 -17937
rect 150004 -17945 150048 -17937
rect 150104 -17945 150148 -17937
rect 150204 -17945 150248 -17937
rect 150304 -17945 150348 -17937
rect 150404 -17945 150448 -17937
rect 150904 -17945 150948 -17937
rect 151004 -17945 151048 -17937
rect 151104 -17945 151148 -17937
rect 151204 -17945 151248 -17937
rect 151304 -17945 151348 -17937
rect 151404 -17945 151448 -17937
rect 151504 -17945 151548 -17937
rect 151604 -17945 151648 -17937
rect 151704 -17945 151748 -17937
rect 151804 -17945 151848 -17937
rect 151904 -17945 151948 -17937
rect 152004 -17945 152048 -17937
rect 152104 -17945 152148 -17937
rect 152204 -17945 152248 -17937
rect 152304 -17945 152348 -17937
rect 152404 -17945 152448 -17937
rect 144948 -17989 144956 -17945
rect 145048 -17989 145056 -17945
rect 145148 -17989 145156 -17945
rect 145248 -17989 145256 -17945
rect 145348 -17989 145356 -17945
rect 145448 -17989 145456 -17945
rect 145548 -17989 145556 -17945
rect 145648 -17989 145656 -17945
rect 145748 -17989 145756 -17945
rect 145848 -17989 145856 -17945
rect 145948 -17989 145956 -17945
rect 146048 -17989 146056 -17945
rect 146148 -17989 146156 -17945
rect 146248 -17989 146256 -17945
rect 146348 -17989 146356 -17945
rect 146448 -17989 146456 -17945
rect 146948 -17989 146956 -17945
rect 147048 -17989 147056 -17945
rect 147148 -17989 147156 -17945
rect 147248 -17989 147256 -17945
rect 147348 -17989 147356 -17945
rect 147448 -17989 147456 -17945
rect 147548 -17989 147556 -17945
rect 147648 -17989 147656 -17945
rect 147748 -17989 147756 -17945
rect 147848 -17989 147856 -17945
rect 147948 -17989 147956 -17945
rect 148048 -17989 148056 -17945
rect 148148 -17989 148156 -17945
rect 148248 -17989 148256 -17945
rect 148348 -17989 148356 -17945
rect 148448 -17989 148456 -17945
rect 148948 -17989 148956 -17945
rect 149048 -17989 149056 -17945
rect 149148 -17989 149156 -17945
rect 149248 -17989 149256 -17945
rect 149348 -17989 149356 -17945
rect 149448 -17989 149456 -17945
rect 149548 -17989 149556 -17945
rect 149648 -17989 149656 -17945
rect 149748 -17989 149756 -17945
rect 149848 -17989 149856 -17945
rect 149948 -17989 149956 -17945
rect 150048 -17989 150056 -17945
rect 150148 -17989 150156 -17945
rect 150248 -17989 150256 -17945
rect 150348 -17989 150356 -17945
rect 150448 -17989 150456 -17945
rect 150948 -17989 150956 -17945
rect 151048 -17989 151056 -17945
rect 151148 -17989 151156 -17945
rect 151248 -17989 151256 -17945
rect 151348 -17989 151356 -17945
rect 151448 -17989 151456 -17945
rect 151548 -17989 151556 -17945
rect 151648 -17989 151656 -17945
rect 151748 -17989 151756 -17945
rect 151848 -17989 151856 -17945
rect 151948 -17989 151956 -17945
rect 152048 -17989 152056 -17945
rect 152148 -17989 152156 -17945
rect 152248 -17989 152256 -17945
rect 152348 -17989 152356 -17945
rect 152448 -17989 152456 -17945
rect 144904 -18045 144948 -18037
rect 145004 -18045 145048 -18037
rect 145104 -18045 145148 -18037
rect 145204 -18045 145248 -18037
rect 145304 -18045 145348 -18037
rect 145404 -18045 145448 -18037
rect 145504 -18045 145548 -18037
rect 145604 -18045 145648 -18037
rect 145704 -18045 145748 -18037
rect 145804 -18045 145848 -18037
rect 145904 -18045 145948 -18037
rect 146004 -18045 146048 -18037
rect 146104 -18045 146148 -18037
rect 146204 -18045 146248 -18037
rect 146304 -18045 146348 -18037
rect 146404 -18045 146448 -18037
rect 146904 -18045 146948 -18037
rect 147004 -18045 147048 -18037
rect 147104 -18045 147148 -18037
rect 147204 -18045 147248 -18037
rect 147304 -18045 147348 -18037
rect 147404 -18045 147448 -18037
rect 147504 -18045 147548 -18037
rect 147604 -18045 147648 -18037
rect 147704 -18045 147748 -18037
rect 147804 -18045 147848 -18037
rect 147904 -18045 147948 -18037
rect 148004 -18045 148048 -18037
rect 148104 -18045 148148 -18037
rect 148204 -18045 148248 -18037
rect 148304 -18045 148348 -18037
rect 148404 -18045 148448 -18037
rect 148904 -18045 148948 -18037
rect 149004 -18045 149048 -18037
rect 149104 -18045 149148 -18037
rect 149204 -18045 149248 -18037
rect 149304 -18045 149348 -18037
rect 149404 -18045 149448 -18037
rect 149504 -18045 149548 -18037
rect 149604 -18045 149648 -18037
rect 149704 -18045 149748 -18037
rect 149804 -18045 149848 -18037
rect 149904 -18045 149948 -18037
rect 150004 -18045 150048 -18037
rect 150104 -18045 150148 -18037
rect 150204 -18045 150248 -18037
rect 150304 -18045 150348 -18037
rect 150404 -18045 150448 -18037
rect 150904 -18045 150948 -18037
rect 151004 -18045 151048 -18037
rect 151104 -18045 151148 -18037
rect 151204 -18045 151248 -18037
rect 151304 -18045 151348 -18037
rect 151404 -18045 151448 -18037
rect 151504 -18045 151548 -18037
rect 151604 -18045 151648 -18037
rect 151704 -18045 151748 -18037
rect 151804 -18045 151848 -18037
rect 151904 -18045 151948 -18037
rect 152004 -18045 152048 -18037
rect 152104 -18045 152148 -18037
rect 152204 -18045 152248 -18037
rect 152304 -18045 152348 -18037
rect 152404 -18045 152448 -18037
rect 144948 -18089 144956 -18045
rect 145048 -18089 145056 -18045
rect 145148 -18089 145156 -18045
rect 145248 -18089 145256 -18045
rect 145348 -18089 145356 -18045
rect 145448 -18089 145456 -18045
rect 145548 -18089 145556 -18045
rect 145648 -18089 145656 -18045
rect 145748 -18089 145756 -18045
rect 145848 -18089 145856 -18045
rect 145948 -18089 145956 -18045
rect 146048 -18089 146056 -18045
rect 146148 -18089 146156 -18045
rect 146248 -18089 146256 -18045
rect 146348 -18089 146356 -18045
rect 146448 -18089 146456 -18045
rect 146948 -18089 146956 -18045
rect 147048 -18089 147056 -18045
rect 147148 -18089 147156 -18045
rect 147248 -18089 147256 -18045
rect 147348 -18089 147356 -18045
rect 147448 -18089 147456 -18045
rect 147548 -18089 147556 -18045
rect 147648 -18089 147656 -18045
rect 147748 -18089 147756 -18045
rect 147848 -18089 147856 -18045
rect 147948 -18089 147956 -18045
rect 148048 -18089 148056 -18045
rect 148148 -18089 148156 -18045
rect 148248 -18089 148256 -18045
rect 148348 -18089 148356 -18045
rect 148448 -18089 148456 -18045
rect 148948 -18089 148956 -18045
rect 149048 -18089 149056 -18045
rect 149148 -18089 149156 -18045
rect 149248 -18089 149256 -18045
rect 149348 -18089 149356 -18045
rect 149448 -18089 149456 -18045
rect 149548 -18089 149556 -18045
rect 149648 -18089 149656 -18045
rect 149748 -18089 149756 -18045
rect 149848 -18089 149856 -18045
rect 149948 -18089 149956 -18045
rect 150048 -18089 150056 -18045
rect 150148 -18089 150156 -18045
rect 150248 -18089 150256 -18045
rect 150348 -18089 150356 -18045
rect 150448 -18089 150456 -18045
rect 150948 -18089 150956 -18045
rect 151048 -18089 151056 -18045
rect 151148 -18089 151156 -18045
rect 151248 -18089 151256 -18045
rect 151348 -18089 151356 -18045
rect 151448 -18089 151456 -18045
rect 151548 -18089 151556 -18045
rect 151648 -18089 151656 -18045
rect 151748 -18089 151756 -18045
rect 151848 -18089 151856 -18045
rect 151948 -18089 151956 -18045
rect 152048 -18089 152056 -18045
rect 152148 -18089 152156 -18045
rect 152248 -18089 152256 -18045
rect 152348 -18089 152356 -18045
rect 152448 -18089 152456 -18045
rect 144904 -18145 144948 -18137
rect 145004 -18145 145048 -18137
rect 145104 -18145 145148 -18137
rect 145204 -18145 145248 -18137
rect 145304 -18145 145348 -18137
rect 145404 -18145 145448 -18137
rect 145504 -18145 145548 -18137
rect 145604 -18145 145648 -18137
rect 145704 -18145 145748 -18137
rect 145804 -18145 145848 -18137
rect 145904 -18145 145948 -18137
rect 146004 -18145 146048 -18137
rect 146104 -18145 146148 -18137
rect 146204 -18145 146248 -18137
rect 146304 -18145 146348 -18137
rect 146404 -18145 146448 -18137
rect 146904 -18145 146948 -18137
rect 147004 -18145 147048 -18137
rect 147104 -18145 147148 -18137
rect 147204 -18145 147248 -18137
rect 147304 -18145 147348 -18137
rect 147404 -18145 147448 -18137
rect 147504 -18145 147548 -18137
rect 147604 -18145 147648 -18137
rect 147704 -18145 147748 -18137
rect 147804 -18145 147848 -18137
rect 147904 -18145 147948 -18137
rect 148004 -18145 148048 -18137
rect 148104 -18145 148148 -18137
rect 148204 -18145 148248 -18137
rect 148304 -18145 148348 -18137
rect 148404 -18145 148448 -18137
rect 148904 -18145 148948 -18137
rect 149004 -18145 149048 -18137
rect 149104 -18145 149148 -18137
rect 149204 -18145 149248 -18137
rect 149304 -18145 149348 -18137
rect 149404 -18145 149448 -18137
rect 149504 -18145 149548 -18137
rect 149604 -18145 149648 -18137
rect 149704 -18145 149748 -18137
rect 149804 -18145 149848 -18137
rect 149904 -18145 149948 -18137
rect 150004 -18145 150048 -18137
rect 150104 -18145 150148 -18137
rect 150204 -18145 150248 -18137
rect 150304 -18145 150348 -18137
rect 150404 -18145 150448 -18137
rect 150904 -18145 150948 -18137
rect 151004 -18145 151048 -18137
rect 151104 -18145 151148 -18137
rect 151204 -18145 151248 -18137
rect 151304 -18145 151348 -18137
rect 151404 -18145 151448 -18137
rect 151504 -18145 151548 -18137
rect 151604 -18145 151648 -18137
rect 151704 -18145 151748 -18137
rect 151804 -18145 151848 -18137
rect 151904 -18145 151948 -18137
rect 152004 -18145 152048 -18137
rect 152104 -18145 152148 -18137
rect 152204 -18145 152248 -18137
rect 152304 -18145 152348 -18137
rect 152404 -18145 152448 -18137
rect 144948 -18189 144956 -18145
rect 145048 -18189 145056 -18145
rect 145148 -18189 145156 -18145
rect 145248 -18189 145256 -18145
rect 145348 -18189 145356 -18145
rect 145448 -18189 145456 -18145
rect 145548 -18189 145556 -18145
rect 145648 -18189 145656 -18145
rect 145748 -18189 145756 -18145
rect 145848 -18189 145856 -18145
rect 145948 -18189 145956 -18145
rect 146048 -18189 146056 -18145
rect 146148 -18189 146156 -18145
rect 146248 -18189 146256 -18145
rect 146348 -18189 146356 -18145
rect 146448 -18189 146456 -18145
rect 146948 -18189 146956 -18145
rect 147048 -18189 147056 -18145
rect 147148 -18189 147156 -18145
rect 147248 -18189 147256 -18145
rect 147348 -18189 147356 -18145
rect 147448 -18189 147456 -18145
rect 147548 -18189 147556 -18145
rect 147648 -18189 147656 -18145
rect 147748 -18189 147756 -18145
rect 147848 -18189 147856 -18145
rect 147948 -18189 147956 -18145
rect 148048 -18189 148056 -18145
rect 148148 -18189 148156 -18145
rect 148248 -18189 148256 -18145
rect 148348 -18189 148356 -18145
rect 148448 -18189 148456 -18145
rect 148948 -18189 148956 -18145
rect 149048 -18189 149056 -18145
rect 149148 -18189 149156 -18145
rect 149248 -18189 149256 -18145
rect 149348 -18189 149356 -18145
rect 149448 -18189 149456 -18145
rect 149548 -18189 149556 -18145
rect 149648 -18189 149656 -18145
rect 149748 -18189 149756 -18145
rect 149848 -18189 149856 -18145
rect 149948 -18189 149956 -18145
rect 150048 -18189 150056 -18145
rect 150148 -18189 150156 -18145
rect 150248 -18189 150256 -18145
rect 150348 -18189 150356 -18145
rect 150448 -18189 150456 -18145
rect 150948 -18189 150956 -18145
rect 151048 -18189 151056 -18145
rect 151148 -18189 151156 -18145
rect 151248 -18189 151256 -18145
rect 151348 -18189 151356 -18145
rect 151448 -18189 151456 -18145
rect 151548 -18189 151556 -18145
rect 151648 -18189 151656 -18145
rect 151748 -18189 151756 -18145
rect 151848 -18189 151856 -18145
rect 151948 -18189 151956 -18145
rect 152048 -18189 152056 -18145
rect 152148 -18189 152156 -18145
rect 152248 -18189 152256 -18145
rect 152348 -18189 152356 -18145
rect 152448 -18189 152456 -18145
rect 144904 -18245 144948 -18237
rect 145004 -18245 145048 -18237
rect 145104 -18245 145148 -18237
rect 145204 -18245 145248 -18237
rect 145304 -18245 145348 -18237
rect 145404 -18245 145448 -18237
rect 145504 -18245 145548 -18237
rect 145604 -18245 145648 -18237
rect 145704 -18245 145748 -18237
rect 145804 -18245 145848 -18237
rect 145904 -18245 145948 -18237
rect 146004 -18245 146048 -18237
rect 146104 -18245 146148 -18237
rect 146204 -18245 146248 -18237
rect 146304 -18245 146348 -18237
rect 146404 -18245 146448 -18237
rect 146904 -18245 146948 -18237
rect 147004 -18245 147048 -18237
rect 147104 -18245 147148 -18237
rect 147204 -18245 147248 -18237
rect 147304 -18245 147348 -18237
rect 147404 -18245 147448 -18237
rect 147504 -18245 147548 -18237
rect 147604 -18245 147648 -18237
rect 147704 -18245 147748 -18237
rect 147804 -18245 147848 -18237
rect 147904 -18245 147948 -18237
rect 148004 -18245 148048 -18237
rect 148104 -18245 148148 -18237
rect 148204 -18245 148248 -18237
rect 148304 -18245 148348 -18237
rect 148404 -18245 148448 -18237
rect 148904 -18245 148948 -18237
rect 149004 -18245 149048 -18237
rect 149104 -18245 149148 -18237
rect 149204 -18245 149248 -18237
rect 149304 -18245 149348 -18237
rect 149404 -18245 149448 -18237
rect 149504 -18245 149548 -18237
rect 149604 -18245 149648 -18237
rect 149704 -18245 149748 -18237
rect 149804 -18245 149848 -18237
rect 149904 -18245 149948 -18237
rect 150004 -18245 150048 -18237
rect 150104 -18245 150148 -18237
rect 150204 -18245 150248 -18237
rect 150304 -18245 150348 -18237
rect 150404 -18245 150448 -18237
rect 150904 -18245 150948 -18237
rect 151004 -18245 151048 -18237
rect 151104 -18245 151148 -18237
rect 151204 -18245 151248 -18237
rect 151304 -18245 151348 -18237
rect 151404 -18245 151448 -18237
rect 151504 -18245 151548 -18237
rect 151604 -18245 151648 -18237
rect 151704 -18245 151748 -18237
rect 151804 -18245 151848 -18237
rect 151904 -18245 151948 -18237
rect 152004 -18245 152048 -18237
rect 152104 -18245 152148 -18237
rect 152204 -18245 152248 -18237
rect 152304 -18245 152348 -18237
rect 152404 -18245 152448 -18237
rect 144948 -18289 144956 -18245
rect 145048 -18289 145056 -18245
rect 145148 -18289 145156 -18245
rect 145248 -18289 145256 -18245
rect 145348 -18289 145356 -18245
rect 145448 -18289 145456 -18245
rect 145548 -18289 145556 -18245
rect 145648 -18289 145656 -18245
rect 145748 -18289 145756 -18245
rect 145848 -18289 145856 -18245
rect 145948 -18289 145956 -18245
rect 146048 -18289 146056 -18245
rect 146148 -18289 146156 -18245
rect 146248 -18289 146256 -18245
rect 146348 -18289 146356 -18245
rect 146448 -18289 146456 -18245
rect 146948 -18289 146956 -18245
rect 147048 -18289 147056 -18245
rect 147148 -18289 147156 -18245
rect 147248 -18289 147256 -18245
rect 147348 -18289 147356 -18245
rect 147448 -18289 147456 -18245
rect 147548 -18289 147556 -18245
rect 147648 -18289 147656 -18245
rect 147748 -18289 147756 -18245
rect 147848 -18289 147856 -18245
rect 147948 -18289 147956 -18245
rect 148048 -18289 148056 -18245
rect 148148 -18289 148156 -18245
rect 148248 -18289 148256 -18245
rect 148348 -18289 148356 -18245
rect 148448 -18289 148456 -18245
rect 148948 -18289 148956 -18245
rect 149048 -18289 149056 -18245
rect 149148 -18289 149156 -18245
rect 149248 -18289 149256 -18245
rect 149348 -18289 149356 -18245
rect 149448 -18289 149456 -18245
rect 149548 -18289 149556 -18245
rect 149648 -18289 149656 -18245
rect 149748 -18289 149756 -18245
rect 149848 -18289 149856 -18245
rect 149948 -18289 149956 -18245
rect 150048 -18289 150056 -18245
rect 150148 -18289 150156 -18245
rect 150248 -18289 150256 -18245
rect 150348 -18289 150356 -18245
rect 150448 -18289 150456 -18245
rect 150948 -18289 150956 -18245
rect 151048 -18289 151056 -18245
rect 151148 -18289 151156 -18245
rect 151248 -18289 151256 -18245
rect 151348 -18289 151356 -18245
rect 151448 -18289 151456 -18245
rect 151548 -18289 151556 -18245
rect 151648 -18289 151656 -18245
rect 151748 -18289 151756 -18245
rect 151848 -18289 151856 -18245
rect 151948 -18289 151956 -18245
rect 152048 -18289 152056 -18245
rect 152148 -18289 152156 -18245
rect 152248 -18289 152256 -18245
rect 152348 -18289 152356 -18245
rect 152448 -18289 152456 -18245
rect 144904 -18345 144948 -18337
rect 145004 -18345 145048 -18337
rect 145104 -18345 145148 -18337
rect 145204 -18345 145248 -18337
rect 145304 -18345 145348 -18337
rect 145404 -18345 145448 -18337
rect 145504 -18345 145548 -18337
rect 145604 -18345 145648 -18337
rect 145704 -18345 145748 -18337
rect 145804 -18345 145848 -18337
rect 145904 -18345 145948 -18337
rect 146004 -18345 146048 -18337
rect 146104 -18345 146148 -18337
rect 146204 -18345 146248 -18337
rect 146304 -18345 146348 -18337
rect 146404 -18345 146448 -18337
rect 146904 -18345 146948 -18337
rect 147004 -18345 147048 -18337
rect 147104 -18345 147148 -18337
rect 147204 -18345 147248 -18337
rect 147304 -18345 147348 -18337
rect 147404 -18345 147448 -18337
rect 147504 -18345 147548 -18337
rect 147604 -18345 147648 -18337
rect 147704 -18345 147748 -18337
rect 147804 -18345 147848 -18337
rect 147904 -18345 147948 -18337
rect 148004 -18345 148048 -18337
rect 148104 -18345 148148 -18337
rect 148204 -18345 148248 -18337
rect 148304 -18345 148348 -18337
rect 148404 -18345 148448 -18337
rect 148904 -18345 148948 -18337
rect 149004 -18345 149048 -18337
rect 149104 -18345 149148 -18337
rect 149204 -18345 149248 -18337
rect 149304 -18345 149348 -18337
rect 149404 -18345 149448 -18337
rect 149504 -18345 149548 -18337
rect 149604 -18345 149648 -18337
rect 149704 -18345 149748 -18337
rect 149804 -18345 149848 -18337
rect 149904 -18345 149948 -18337
rect 150004 -18345 150048 -18337
rect 150104 -18345 150148 -18337
rect 150204 -18345 150248 -18337
rect 150304 -18345 150348 -18337
rect 150404 -18345 150448 -18337
rect 150904 -18345 150948 -18337
rect 151004 -18345 151048 -18337
rect 151104 -18345 151148 -18337
rect 151204 -18345 151248 -18337
rect 151304 -18345 151348 -18337
rect 151404 -18345 151448 -18337
rect 151504 -18345 151548 -18337
rect 151604 -18345 151648 -18337
rect 151704 -18345 151748 -18337
rect 151804 -18345 151848 -18337
rect 151904 -18345 151948 -18337
rect 152004 -18345 152048 -18337
rect 152104 -18345 152148 -18337
rect 152204 -18345 152248 -18337
rect 152304 -18345 152348 -18337
rect 152404 -18345 152448 -18337
rect 144948 -18389 144956 -18345
rect 145048 -18389 145056 -18345
rect 145148 -18389 145156 -18345
rect 145248 -18389 145256 -18345
rect 145348 -18389 145356 -18345
rect 145448 -18389 145456 -18345
rect 145548 -18389 145556 -18345
rect 145648 -18389 145656 -18345
rect 145748 -18389 145756 -18345
rect 145848 -18389 145856 -18345
rect 145948 -18389 145956 -18345
rect 146048 -18389 146056 -18345
rect 146148 -18389 146156 -18345
rect 146248 -18389 146256 -18345
rect 146348 -18389 146356 -18345
rect 146448 -18389 146456 -18345
rect 146948 -18389 146956 -18345
rect 147048 -18389 147056 -18345
rect 147148 -18389 147156 -18345
rect 147248 -18389 147256 -18345
rect 147348 -18389 147356 -18345
rect 147448 -18389 147456 -18345
rect 147548 -18389 147556 -18345
rect 147648 -18389 147656 -18345
rect 147748 -18389 147756 -18345
rect 147848 -18389 147856 -18345
rect 147948 -18389 147956 -18345
rect 148048 -18389 148056 -18345
rect 148148 -18389 148156 -18345
rect 148248 -18389 148256 -18345
rect 148348 -18389 148356 -18345
rect 148448 -18389 148456 -18345
rect 148948 -18389 148956 -18345
rect 149048 -18389 149056 -18345
rect 149148 -18389 149156 -18345
rect 149248 -18389 149256 -18345
rect 149348 -18389 149356 -18345
rect 149448 -18389 149456 -18345
rect 149548 -18389 149556 -18345
rect 149648 -18389 149656 -18345
rect 149748 -18389 149756 -18345
rect 149848 -18389 149856 -18345
rect 149948 -18389 149956 -18345
rect 150048 -18389 150056 -18345
rect 150148 -18389 150156 -18345
rect 150248 -18389 150256 -18345
rect 150348 -18389 150356 -18345
rect 150448 -18389 150456 -18345
rect 150948 -18389 150956 -18345
rect 151048 -18389 151056 -18345
rect 151148 -18389 151156 -18345
rect 151248 -18389 151256 -18345
rect 151348 -18389 151356 -18345
rect 151448 -18389 151456 -18345
rect 151548 -18389 151556 -18345
rect 151648 -18389 151656 -18345
rect 151748 -18389 151756 -18345
rect 151848 -18389 151856 -18345
rect 151948 -18389 151956 -18345
rect 152048 -18389 152056 -18345
rect 152148 -18389 152156 -18345
rect 152248 -18389 152256 -18345
rect 152348 -18389 152356 -18345
rect 152448 -18389 152456 -18345
rect 144904 -18445 144948 -18437
rect 145004 -18445 145048 -18437
rect 145104 -18445 145148 -18437
rect 145204 -18445 145248 -18437
rect 145304 -18445 145348 -18437
rect 145404 -18445 145448 -18437
rect 145504 -18445 145548 -18437
rect 145604 -18445 145648 -18437
rect 145704 -18445 145748 -18437
rect 145804 -18445 145848 -18437
rect 145904 -18445 145948 -18437
rect 146004 -18445 146048 -18437
rect 146104 -18445 146148 -18437
rect 146204 -18445 146248 -18437
rect 146304 -18445 146348 -18437
rect 146404 -18445 146448 -18437
rect 146904 -18445 146948 -18437
rect 147004 -18445 147048 -18437
rect 147104 -18445 147148 -18437
rect 147204 -18445 147248 -18437
rect 147304 -18445 147348 -18437
rect 147404 -18445 147448 -18437
rect 147504 -18445 147548 -18437
rect 147604 -18445 147648 -18437
rect 147704 -18445 147748 -18437
rect 147804 -18445 147848 -18437
rect 147904 -18445 147948 -18437
rect 148004 -18445 148048 -18437
rect 148104 -18445 148148 -18437
rect 148204 -18445 148248 -18437
rect 148304 -18445 148348 -18437
rect 148404 -18445 148448 -18437
rect 148904 -18445 148948 -18437
rect 149004 -18445 149048 -18437
rect 149104 -18445 149148 -18437
rect 149204 -18445 149248 -18437
rect 149304 -18445 149348 -18437
rect 149404 -18445 149448 -18437
rect 149504 -18445 149548 -18437
rect 149604 -18445 149648 -18437
rect 149704 -18445 149748 -18437
rect 149804 -18445 149848 -18437
rect 149904 -18445 149948 -18437
rect 150004 -18445 150048 -18437
rect 150104 -18445 150148 -18437
rect 150204 -18445 150248 -18437
rect 150304 -18445 150348 -18437
rect 150404 -18445 150448 -18437
rect 150904 -18445 150948 -18437
rect 151004 -18445 151048 -18437
rect 151104 -18445 151148 -18437
rect 151204 -18445 151248 -18437
rect 151304 -18445 151348 -18437
rect 151404 -18445 151448 -18437
rect 151504 -18445 151548 -18437
rect 151604 -18445 151648 -18437
rect 151704 -18445 151748 -18437
rect 151804 -18445 151848 -18437
rect 151904 -18445 151948 -18437
rect 152004 -18445 152048 -18437
rect 152104 -18445 152148 -18437
rect 152204 -18445 152248 -18437
rect 152304 -18445 152348 -18437
rect 152404 -18445 152448 -18437
rect 144948 -18489 144956 -18445
rect 145048 -18489 145056 -18445
rect 145148 -18489 145156 -18445
rect 145248 -18489 145256 -18445
rect 145348 -18489 145356 -18445
rect 145448 -18489 145456 -18445
rect 145548 -18489 145556 -18445
rect 145648 -18489 145656 -18445
rect 145748 -18489 145756 -18445
rect 145848 -18489 145856 -18445
rect 145948 -18489 145956 -18445
rect 146048 -18489 146056 -18445
rect 146148 -18489 146156 -18445
rect 146248 -18489 146256 -18445
rect 146348 -18489 146356 -18445
rect 146448 -18489 146456 -18445
rect 146948 -18489 146956 -18445
rect 147048 -18489 147056 -18445
rect 147148 -18489 147156 -18445
rect 147248 -18489 147256 -18445
rect 147348 -18489 147356 -18445
rect 147448 -18489 147456 -18445
rect 147548 -18489 147556 -18445
rect 147648 -18489 147656 -18445
rect 147748 -18489 147756 -18445
rect 147848 -18489 147856 -18445
rect 147948 -18489 147956 -18445
rect 148048 -18489 148056 -18445
rect 148148 -18489 148156 -18445
rect 148248 -18489 148256 -18445
rect 148348 -18489 148356 -18445
rect 148448 -18489 148456 -18445
rect 148948 -18489 148956 -18445
rect 149048 -18489 149056 -18445
rect 149148 -18489 149156 -18445
rect 149248 -18489 149256 -18445
rect 149348 -18489 149356 -18445
rect 149448 -18489 149456 -18445
rect 149548 -18489 149556 -18445
rect 149648 -18489 149656 -18445
rect 149748 -18489 149756 -18445
rect 149848 -18489 149856 -18445
rect 149948 -18489 149956 -18445
rect 150048 -18489 150056 -18445
rect 150148 -18489 150156 -18445
rect 150248 -18489 150256 -18445
rect 150348 -18489 150356 -18445
rect 150448 -18489 150456 -18445
rect 150948 -18489 150956 -18445
rect 151048 -18489 151056 -18445
rect 151148 -18489 151156 -18445
rect 151248 -18489 151256 -18445
rect 151348 -18489 151356 -18445
rect 151448 -18489 151456 -18445
rect 151548 -18489 151556 -18445
rect 151648 -18489 151656 -18445
rect 151748 -18489 151756 -18445
rect 151848 -18489 151856 -18445
rect 151948 -18489 151956 -18445
rect 152048 -18489 152056 -18445
rect 152148 -18489 152156 -18445
rect 152248 -18489 152256 -18445
rect 152348 -18489 152356 -18445
rect 152448 -18489 152456 -18445
rect 144904 -18545 144948 -18537
rect 145004 -18545 145048 -18537
rect 145104 -18545 145148 -18537
rect 145204 -18545 145248 -18537
rect 145304 -18545 145348 -18537
rect 145404 -18545 145448 -18537
rect 145504 -18545 145548 -18537
rect 145604 -18545 145648 -18537
rect 145704 -18545 145748 -18537
rect 145804 -18545 145848 -18537
rect 145904 -18545 145948 -18537
rect 146004 -18545 146048 -18537
rect 146104 -18545 146148 -18537
rect 146204 -18545 146248 -18537
rect 146304 -18545 146348 -18537
rect 146404 -18545 146448 -18537
rect 146904 -18545 146948 -18537
rect 147004 -18545 147048 -18537
rect 147104 -18545 147148 -18537
rect 147204 -18545 147248 -18537
rect 147304 -18545 147348 -18537
rect 147404 -18545 147448 -18537
rect 147504 -18545 147548 -18537
rect 147604 -18545 147648 -18537
rect 147704 -18545 147748 -18537
rect 147804 -18545 147848 -18537
rect 147904 -18545 147948 -18537
rect 148004 -18545 148048 -18537
rect 148104 -18545 148148 -18537
rect 148204 -18545 148248 -18537
rect 148304 -18545 148348 -18537
rect 148404 -18545 148448 -18537
rect 148904 -18545 148948 -18537
rect 149004 -18545 149048 -18537
rect 149104 -18545 149148 -18537
rect 149204 -18545 149248 -18537
rect 149304 -18545 149348 -18537
rect 149404 -18545 149448 -18537
rect 149504 -18545 149548 -18537
rect 149604 -18545 149648 -18537
rect 149704 -18545 149748 -18537
rect 149804 -18545 149848 -18537
rect 149904 -18545 149948 -18537
rect 150004 -18545 150048 -18537
rect 150104 -18545 150148 -18537
rect 150204 -18545 150248 -18537
rect 150304 -18545 150348 -18537
rect 150404 -18545 150448 -18537
rect 150904 -18545 150948 -18537
rect 151004 -18545 151048 -18537
rect 151104 -18545 151148 -18537
rect 151204 -18545 151248 -18537
rect 151304 -18545 151348 -18537
rect 151404 -18545 151448 -18537
rect 151504 -18545 151548 -18537
rect 151604 -18545 151648 -18537
rect 151704 -18545 151748 -18537
rect 151804 -18545 151848 -18537
rect 151904 -18545 151948 -18537
rect 152004 -18545 152048 -18537
rect 152104 -18545 152148 -18537
rect 152204 -18545 152248 -18537
rect 152304 -18545 152348 -18537
rect 152404 -18545 152448 -18537
rect 144948 -18589 144956 -18545
rect 145048 -18589 145056 -18545
rect 145148 -18589 145156 -18545
rect 145248 -18589 145256 -18545
rect 145348 -18589 145356 -18545
rect 145448 -18589 145456 -18545
rect 145548 -18589 145556 -18545
rect 145648 -18589 145656 -18545
rect 145748 -18589 145756 -18545
rect 145848 -18589 145856 -18545
rect 145948 -18589 145956 -18545
rect 146048 -18589 146056 -18545
rect 146148 -18589 146156 -18545
rect 146248 -18589 146256 -18545
rect 146348 -18589 146356 -18545
rect 146448 -18589 146456 -18545
rect 146948 -18589 146956 -18545
rect 147048 -18589 147056 -18545
rect 147148 -18589 147156 -18545
rect 147248 -18589 147256 -18545
rect 147348 -18589 147356 -18545
rect 147448 -18589 147456 -18545
rect 147548 -18589 147556 -18545
rect 147648 -18589 147656 -18545
rect 147748 -18589 147756 -18545
rect 147848 -18589 147856 -18545
rect 147948 -18589 147956 -18545
rect 148048 -18589 148056 -18545
rect 148148 -18589 148156 -18545
rect 148248 -18589 148256 -18545
rect 148348 -18589 148356 -18545
rect 148448 -18589 148456 -18545
rect 148948 -18589 148956 -18545
rect 149048 -18589 149056 -18545
rect 149148 -18589 149156 -18545
rect 149248 -18589 149256 -18545
rect 149348 -18589 149356 -18545
rect 149448 -18589 149456 -18545
rect 149548 -18589 149556 -18545
rect 149648 -18589 149656 -18545
rect 149748 -18589 149756 -18545
rect 149848 -18589 149856 -18545
rect 149948 -18589 149956 -18545
rect 150048 -18589 150056 -18545
rect 150148 -18589 150156 -18545
rect 150248 -18589 150256 -18545
rect 150348 -18589 150356 -18545
rect 150448 -18589 150456 -18545
rect 150948 -18589 150956 -18545
rect 151048 -18589 151056 -18545
rect 151148 -18589 151156 -18545
rect 151248 -18589 151256 -18545
rect 151348 -18589 151356 -18545
rect 151448 -18589 151456 -18545
rect 151548 -18589 151556 -18545
rect 151648 -18589 151656 -18545
rect 151748 -18589 151756 -18545
rect 151848 -18589 151856 -18545
rect 151948 -18589 151956 -18545
rect 152048 -18589 152056 -18545
rect 152148 -18589 152156 -18545
rect 152248 -18589 152256 -18545
rect 152348 -18589 152356 -18545
rect 152448 -18589 152456 -18545
rect 144904 -18645 144948 -18637
rect 145004 -18645 145048 -18637
rect 145104 -18645 145148 -18637
rect 145204 -18645 145248 -18637
rect 145304 -18645 145348 -18637
rect 145404 -18645 145448 -18637
rect 145504 -18645 145548 -18637
rect 145604 -18645 145648 -18637
rect 145704 -18645 145748 -18637
rect 145804 -18645 145848 -18637
rect 145904 -18645 145948 -18637
rect 146004 -18645 146048 -18637
rect 146104 -18645 146148 -18637
rect 146204 -18645 146248 -18637
rect 146304 -18645 146348 -18637
rect 146404 -18645 146448 -18637
rect 146904 -18645 146948 -18637
rect 147004 -18645 147048 -18637
rect 147104 -18645 147148 -18637
rect 147204 -18645 147248 -18637
rect 147304 -18645 147348 -18637
rect 147404 -18645 147448 -18637
rect 147504 -18645 147548 -18637
rect 147604 -18645 147648 -18637
rect 147704 -18645 147748 -18637
rect 147804 -18645 147848 -18637
rect 147904 -18645 147948 -18637
rect 148004 -18645 148048 -18637
rect 148104 -18645 148148 -18637
rect 148204 -18645 148248 -18637
rect 148304 -18645 148348 -18637
rect 148404 -18645 148448 -18637
rect 148904 -18645 148948 -18637
rect 149004 -18645 149048 -18637
rect 149104 -18645 149148 -18637
rect 149204 -18645 149248 -18637
rect 149304 -18645 149348 -18637
rect 149404 -18645 149448 -18637
rect 149504 -18645 149548 -18637
rect 149604 -18645 149648 -18637
rect 149704 -18645 149748 -18637
rect 149804 -18645 149848 -18637
rect 149904 -18645 149948 -18637
rect 150004 -18645 150048 -18637
rect 150104 -18645 150148 -18637
rect 150204 -18645 150248 -18637
rect 150304 -18645 150348 -18637
rect 150404 -18645 150448 -18637
rect 150904 -18645 150948 -18637
rect 151004 -18645 151048 -18637
rect 151104 -18645 151148 -18637
rect 151204 -18645 151248 -18637
rect 151304 -18645 151348 -18637
rect 151404 -18645 151448 -18637
rect 151504 -18645 151548 -18637
rect 151604 -18645 151648 -18637
rect 151704 -18645 151748 -18637
rect 151804 -18645 151848 -18637
rect 151904 -18645 151948 -18637
rect 152004 -18645 152048 -18637
rect 152104 -18645 152148 -18637
rect 152204 -18645 152248 -18637
rect 152304 -18645 152348 -18637
rect 152404 -18645 152448 -18637
rect 144948 -18689 144956 -18645
rect 145048 -18689 145056 -18645
rect 145148 -18689 145156 -18645
rect 145248 -18689 145256 -18645
rect 145348 -18689 145356 -18645
rect 145448 -18689 145456 -18645
rect 145548 -18689 145556 -18645
rect 145648 -18689 145656 -18645
rect 145748 -18689 145756 -18645
rect 145848 -18689 145856 -18645
rect 145948 -18689 145956 -18645
rect 146048 -18689 146056 -18645
rect 146148 -18689 146156 -18645
rect 146248 -18689 146256 -18645
rect 146348 -18689 146356 -18645
rect 146448 -18689 146456 -18645
rect 146948 -18689 146956 -18645
rect 147048 -18689 147056 -18645
rect 147148 -18689 147156 -18645
rect 147248 -18689 147256 -18645
rect 147348 -18689 147356 -18645
rect 147448 -18689 147456 -18645
rect 147548 -18689 147556 -18645
rect 147648 -18689 147656 -18645
rect 147748 -18689 147756 -18645
rect 147848 -18689 147856 -18645
rect 147948 -18689 147956 -18645
rect 148048 -18689 148056 -18645
rect 148148 -18689 148156 -18645
rect 148248 -18689 148256 -18645
rect 148348 -18689 148356 -18645
rect 148448 -18689 148456 -18645
rect 148948 -18689 148956 -18645
rect 149048 -18689 149056 -18645
rect 149148 -18689 149156 -18645
rect 149248 -18689 149256 -18645
rect 149348 -18689 149356 -18645
rect 149448 -18689 149456 -18645
rect 149548 -18689 149556 -18645
rect 149648 -18689 149656 -18645
rect 149748 -18689 149756 -18645
rect 149848 -18689 149856 -18645
rect 149948 -18689 149956 -18645
rect 150048 -18689 150056 -18645
rect 150148 -18689 150156 -18645
rect 150248 -18689 150256 -18645
rect 150348 -18689 150356 -18645
rect 150448 -18689 150456 -18645
rect 150948 -18689 150956 -18645
rect 151048 -18689 151056 -18645
rect 151148 -18689 151156 -18645
rect 151248 -18689 151256 -18645
rect 151348 -18689 151356 -18645
rect 151448 -18689 151456 -18645
rect 151548 -18689 151556 -18645
rect 151648 -18689 151656 -18645
rect 151748 -18689 151756 -18645
rect 151848 -18689 151856 -18645
rect 151948 -18689 151956 -18645
rect 152048 -18689 152056 -18645
rect 152148 -18689 152156 -18645
rect 152248 -18689 152256 -18645
rect 152348 -18689 152356 -18645
rect 152448 -18689 152456 -18645
rect 144904 -18745 144948 -18737
rect 145004 -18745 145048 -18737
rect 145104 -18745 145148 -18737
rect 145204 -18745 145248 -18737
rect 145304 -18745 145348 -18737
rect 145404 -18745 145448 -18737
rect 145504 -18745 145548 -18737
rect 145604 -18745 145648 -18737
rect 145704 -18745 145748 -18737
rect 145804 -18745 145848 -18737
rect 145904 -18745 145948 -18737
rect 146004 -18745 146048 -18737
rect 146104 -18745 146148 -18737
rect 146204 -18745 146248 -18737
rect 146304 -18745 146348 -18737
rect 146404 -18745 146448 -18737
rect 146904 -18745 146948 -18737
rect 147004 -18745 147048 -18737
rect 147104 -18745 147148 -18737
rect 147204 -18745 147248 -18737
rect 147304 -18745 147348 -18737
rect 147404 -18745 147448 -18737
rect 147504 -18745 147548 -18737
rect 147604 -18745 147648 -18737
rect 147704 -18745 147748 -18737
rect 147804 -18745 147848 -18737
rect 147904 -18745 147948 -18737
rect 148004 -18745 148048 -18737
rect 148104 -18745 148148 -18737
rect 148204 -18745 148248 -18737
rect 148304 -18745 148348 -18737
rect 148404 -18745 148448 -18737
rect 148904 -18745 148948 -18737
rect 149004 -18745 149048 -18737
rect 149104 -18745 149148 -18737
rect 149204 -18745 149248 -18737
rect 149304 -18745 149348 -18737
rect 149404 -18745 149448 -18737
rect 149504 -18745 149548 -18737
rect 149604 -18745 149648 -18737
rect 149704 -18745 149748 -18737
rect 149804 -18745 149848 -18737
rect 149904 -18745 149948 -18737
rect 150004 -18745 150048 -18737
rect 150104 -18745 150148 -18737
rect 150204 -18745 150248 -18737
rect 150304 -18745 150348 -18737
rect 150404 -18745 150448 -18737
rect 150904 -18745 150948 -18737
rect 151004 -18745 151048 -18737
rect 151104 -18745 151148 -18737
rect 151204 -18745 151248 -18737
rect 151304 -18745 151348 -18737
rect 151404 -18745 151448 -18737
rect 151504 -18745 151548 -18737
rect 151604 -18745 151648 -18737
rect 151704 -18745 151748 -18737
rect 151804 -18745 151848 -18737
rect 151904 -18745 151948 -18737
rect 152004 -18745 152048 -18737
rect 152104 -18745 152148 -18737
rect 152204 -18745 152248 -18737
rect 152304 -18745 152348 -18737
rect 152404 -18745 152448 -18737
rect 144948 -18789 144956 -18745
rect 145048 -18789 145056 -18745
rect 145148 -18789 145156 -18745
rect 145248 -18789 145256 -18745
rect 145348 -18789 145356 -18745
rect 145448 -18789 145456 -18745
rect 145548 -18789 145556 -18745
rect 145648 -18789 145656 -18745
rect 145748 -18789 145756 -18745
rect 145848 -18789 145856 -18745
rect 145948 -18789 145956 -18745
rect 146048 -18789 146056 -18745
rect 146148 -18789 146156 -18745
rect 146248 -18789 146256 -18745
rect 146348 -18789 146356 -18745
rect 146448 -18789 146456 -18745
rect 146948 -18789 146956 -18745
rect 147048 -18789 147056 -18745
rect 147148 -18789 147156 -18745
rect 147248 -18789 147256 -18745
rect 147348 -18789 147356 -18745
rect 147448 -18789 147456 -18745
rect 147548 -18789 147556 -18745
rect 147648 -18789 147656 -18745
rect 147748 -18789 147756 -18745
rect 147848 -18789 147856 -18745
rect 147948 -18789 147956 -18745
rect 148048 -18789 148056 -18745
rect 148148 -18789 148156 -18745
rect 148248 -18789 148256 -18745
rect 148348 -18789 148356 -18745
rect 148448 -18789 148456 -18745
rect 148948 -18789 148956 -18745
rect 149048 -18789 149056 -18745
rect 149148 -18789 149156 -18745
rect 149248 -18789 149256 -18745
rect 149348 -18789 149356 -18745
rect 149448 -18789 149456 -18745
rect 149548 -18789 149556 -18745
rect 149648 -18789 149656 -18745
rect 149748 -18789 149756 -18745
rect 149848 -18789 149856 -18745
rect 149948 -18789 149956 -18745
rect 150048 -18789 150056 -18745
rect 150148 -18789 150156 -18745
rect 150248 -18789 150256 -18745
rect 150348 -18789 150356 -18745
rect 150448 -18789 150456 -18745
rect 150948 -18789 150956 -18745
rect 151048 -18789 151056 -18745
rect 151148 -18789 151156 -18745
rect 151248 -18789 151256 -18745
rect 151348 -18789 151356 -18745
rect 151448 -18789 151456 -18745
rect 151548 -18789 151556 -18745
rect 151648 -18789 151656 -18745
rect 151748 -18789 151756 -18745
rect 151848 -18789 151856 -18745
rect 151948 -18789 151956 -18745
rect 152048 -18789 152056 -18745
rect 152148 -18789 152156 -18745
rect 152248 -18789 152256 -18745
rect 152348 -18789 152356 -18745
rect 152448 -18789 152456 -18745
rect 144904 -18845 144948 -18837
rect 145004 -18845 145048 -18837
rect 145104 -18845 145148 -18837
rect 145204 -18845 145248 -18837
rect 145304 -18845 145348 -18837
rect 145404 -18845 145448 -18837
rect 145504 -18845 145548 -18837
rect 145604 -18845 145648 -18837
rect 145704 -18845 145748 -18837
rect 145804 -18845 145848 -18837
rect 145904 -18845 145948 -18837
rect 146004 -18845 146048 -18837
rect 146104 -18845 146148 -18837
rect 146204 -18845 146248 -18837
rect 146304 -18845 146348 -18837
rect 146404 -18845 146448 -18837
rect 146904 -18845 146948 -18837
rect 147004 -18845 147048 -18837
rect 147104 -18845 147148 -18837
rect 147204 -18845 147248 -18837
rect 147304 -18845 147348 -18837
rect 147404 -18845 147448 -18837
rect 147504 -18845 147548 -18837
rect 147604 -18845 147648 -18837
rect 147704 -18845 147748 -18837
rect 147804 -18845 147848 -18837
rect 147904 -18845 147948 -18837
rect 148004 -18845 148048 -18837
rect 148104 -18845 148148 -18837
rect 148204 -18845 148248 -18837
rect 148304 -18845 148348 -18837
rect 148404 -18845 148448 -18837
rect 148904 -18845 148948 -18837
rect 149004 -18845 149048 -18837
rect 149104 -18845 149148 -18837
rect 149204 -18845 149248 -18837
rect 149304 -18845 149348 -18837
rect 149404 -18845 149448 -18837
rect 149504 -18845 149548 -18837
rect 149604 -18845 149648 -18837
rect 149704 -18845 149748 -18837
rect 149804 -18845 149848 -18837
rect 149904 -18845 149948 -18837
rect 150004 -18845 150048 -18837
rect 150104 -18845 150148 -18837
rect 150204 -18845 150248 -18837
rect 150304 -18845 150348 -18837
rect 150404 -18845 150448 -18837
rect 150904 -18845 150948 -18837
rect 151004 -18845 151048 -18837
rect 151104 -18845 151148 -18837
rect 151204 -18845 151248 -18837
rect 151304 -18845 151348 -18837
rect 151404 -18845 151448 -18837
rect 151504 -18845 151548 -18837
rect 151604 -18845 151648 -18837
rect 151704 -18845 151748 -18837
rect 151804 -18845 151848 -18837
rect 151904 -18845 151948 -18837
rect 152004 -18845 152048 -18837
rect 152104 -18845 152148 -18837
rect 152204 -18845 152248 -18837
rect 152304 -18845 152348 -18837
rect 152404 -18845 152448 -18837
rect 144948 -18889 144956 -18845
rect 145048 -18889 145056 -18845
rect 145148 -18889 145156 -18845
rect 145248 -18889 145256 -18845
rect 145348 -18889 145356 -18845
rect 145448 -18889 145456 -18845
rect 145548 -18889 145556 -18845
rect 145648 -18889 145656 -18845
rect 145748 -18889 145756 -18845
rect 145848 -18889 145856 -18845
rect 145948 -18889 145956 -18845
rect 146048 -18889 146056 -18845
rect 146148 -18889 146156 -18845
rect 146248 -18889 146256 -18845
rect 146348 -18889 146356 -18845
rect 146448 -18889 146456 -18845
rect 146948 -18889 146956 -18845
rect 147048 -18889 147056 -18845
rect 147148 -18889 147156 -18845
rect 147248 -18889 147256 -18845
rect 147348 -18889 147356 -18845
rect 147448 -18889 147456 -18845
rect 147548 -18889 147556 -18845
rect 147648 -18889 147656 -18845
rect 147748 -18889 147756 -18845
rect 147848 -18889 147856 -18845
rect 147948 -18889 147956 -18845
rect 148048 -18889 148056 -18845
rect 148148 -18889 148156 -18845
rect 148248 -18889 148256 -18845
rect 148348 -18889 148356 -18845
rect 148448 -18889 148456 -18845
rect 148948 -18889 148956 -18845
rect 149048 -18889 149056 -18845
rect 149148 -18889 149156 -18845
rect 149248 -18889 149256 -18845
rect 149348 -18889 149356 -18845
rect 149448 -18889 149456 -18845
rect 149548 -18889 149556 -18845
rect 149648 -18889 149656 -18845
rect 149748 -18889 149756 -18845
rect 149848 -18889 149856 -18845
rect 149948 -18889 149956 -18845
rect 150048 -18889 150056 -18845
rect 150148 -18889 150156 -18845
rect 150248 -18889 150256 -18845
rect 150348 -18889 150356 -18845
rect 150448 -18889 150456 -18845
rect 150948 -18889 150956 -18845
rect 151048 -18889 151056 -18845
rect 151148 -18889 151156 -18845
rect 151248 -18889 151256 -18845
rect 151348 -18889 151356 -18845
rect 151448 -18889 151456 -18845
rect 151548 -18889 151556 -18845
rect 151648 -18889 151656 -18845
rect 151748 -18889 151756 -18845
rect 151848 -18889 151856 -18845
rect 151948 -18889 151956 -18845
rect 152048 -18889 152056 -18845
rect 152148 -18889 152156 -18845
rect 152248 -18889 152256 -18845
rect 152348 -18889 152356 -18845
rect 152448 -18889 152456 -18845
rect 144904 -18945 144948 -18937
rect 145004 -18945 145048 -18937
rect 145104 -18945 145148 -18937
rect 145204 -18945 145248 -18937
rect 145304 -18945 145348 -18937
rect 145404 -18945 145448 -18937
rect 145504 -18945 145548 -18937
rect 145604 -18945 145648 -18937
rect 145704 -18945 145748 -18937
rect 145804 -18945 145848 -18937
rect 145904 -18945 145948 -18937
rect 146004 -18945 146048 -18937
rect 146104 -18945 146148 -18937
rect 146204 -18945 146248 -18937
rect 146304 -18945 146348 -18937
rect 146404 -18945 146448 -18937
rect 146904 -18945 146948 -18937
rect 147004 -18945 147048 -18937
rect 147104 -18945 147148 -18937
rect 147204 -18945 147248 -18937
rect 147304 -18945 147348 -18937
rect 147404 -18945 147448 -18937
rect 147504 -18945 147548 -18937
rect 147604 -18945 147648 -18937
rect 147704 -18945 147748 -18937
rect 147804 -18945 147848 -18937
rect 147904 -18945 147948 -18937
rect 148004 -18945 148048 -18937
rect 148104 -18945 148148 -18937
rect 148204 -18945 148248 -18937
rect 148304 -18945 148348 -18937
rect 148404 -18945 148448 -18937
rect 148904 -18945 148948 -18937
rect 149004 -18945 149048 -18937
rect 149104 -18945 149148 -18937
rect 149204 -18945 149248 -18937
rect 149304 -18945 149348 -18937
rect 149404 -18945 149448 -18937
rect 149504 -18945 149548 -18937
rect 149604 -18945 149648 -18937
rect 149704 -18945 149748 -18937
rect 149804 -18945 149848 -18937
rect 149904 -18945 149948 -18937
rect 150004 -18945 150048 -18937
rect 150104 -18945 150148 -18937
rect 150204 -18945 150248 -18937
rect 150304 -18945 150348 -18937
rect 150404 -18945 150448 -18937
rect 150904 -18945 150948 -18937
rect 151004 -18945 151048 -18937
rect 151104 -18945 151148 -18937
rect 151204 -18945 151248 -18937
rect 151304 -18945 151348 -18937
rect 151404 -18945 151448 -18937
rect 151504 -18945 151548 -18937
rect 151604 -18945 151648 -18937
rect 151704 -18945 151748 -18937
rect 151804 -18945 151848 -18937
rect 151904 -18945 151948 -18937
rect 152004 -18945 152048 -18937
rect 152104 -18945 152148 -18937
rect 152204 -18945 152248 -18937
rect 152304 -18945 152348 -18937
rect 152404 -18945 152448 -18937
rect 144948 -18989 144956 -18945
rect 145048 -18989 145056 -18945
rect 145148 -18989 145156 -18945
rect 145248 -18989 145256 -18945
rect 145348 -18989 145356 -18945
rect 145448 -18989 145456 -18945
rect 145548 -18989 145556 -18945
rect 145648 -18989 145656 -18945
rect 145748 -18989 145756 -18945
rect 145848 -18989 145856 -18945
rect 145948 -18989 145956 -18945
rect 146048 -18989 146056 -18945
rect 146148 -18989 146156 -18945
rect 146248 -18989 146256 -18945
rect 146348 -18989 146356 -18945
rect 146448 -18989 146456 -18945
rect 146948 -18989 146956 -18945
rect 147048 -18989 147056 -18945
rect 147148 -18989 147156 -18945
rect 147248 -18989 147256 -18945
rect 147348 -18989 147356 -18945
rect 147448 -18989 147456 -18945
rect 147548 -18989 147556 -18945
rect 147648 -18989 147656 -18945
rect 147748 -18989 147756 -18945
rect 147848 -18989 147856 -18945
rect 147948 -18989 147956 -18945
rect 148048 -18989 148056 -18945
rect 148148 -18989 148156 -18945
rect 148248 -18989 148256 -18945
rect 148348 -18989 148356 -18945
rect 148448 -18989 148456 -18945
rect 148948 -18989 148956 -18945
rect 149048 -18989 149056 -18945
rect 149148 -18989 149156 -18945
rect 149248 -18989 149256 -18945
rect 149348 -18989 149356 -18945
rect 149448 -18989 149456 -18945
rect 149548 -18989 149556 -18945
rect 149648 -18989 149656 -18945
rect 149748 -18989 149756 -18945
rect 149848 -18989 149856 -18945
rect 149948 -18989 149956 -18945
rect 150048 -18989 150056 -18945
rect 150148 -18989 150156 -18945
rect 150248 -18989 150256 -18945
rect 150348 -18989 150356 -18945
rect 150448 -18989 150456 -18945
rect 150948 -18989 150956 -18945
rect 151048 -18989 151056 -18945
rect 151148 -18989 151156 -18945
rect 151248 -18989 151256 -18945
rect 151348 -18989 151356 -18945
rect 151448 -18989 151456 -18945
rect 151548 -18989 151556 -18945
rect 151648 -18989 151656 -18945
rect 151748 -18989 151756 -18945
rect 151848 -18989 151856 -18945
rect 151948 -18989 151956 -18945
rect 152048 -18989 152056 -18945
rect 152148 -18989 152156 -18945
rect 152248 -18989 152256 -18945
rect 152348 -18989 152356 -18945
rect 152448 -18989 152456 -18945
rect -82799 -24366 -82755 -24358
rect -82699 -24366 -82655 -24358
rect -82599 -24366 -82555 -24358
rect -82499 -24366 -82455 -24358
rect -82399 -24366 -82355 -24358
rect -82299 -24366 -82255 -24358
rect -82199 -24366 -82155 -24358
rect -82099 -24366 -82055 -24358
rect -81999 -24366 -81955 -24358
rect -81899 -24366 -81855 -24358
rect -81799 -24366 -81755 -24358
rect -81699 -24366 -81655 -24358
rect -81599 -24366 -81555 -24358
rect -81499 -24366 -81455 -24358
rect -81399 -24366 -81355 -24358
rect -81299 -24366 -81255 -24358
rect -80799 -24366 -80755 -24358
rect -80699 -24366 -80655 -24358
rect -80599 -24366 -80555 -24358
rect -80499 -24366 -80455 -24358
rect -80399 -24366 -80355 -24358
rect -80299 -24366 -80255 -24358
rect -80199 -24366 -80155 -24358
rect -80099 -24366 -80055 -24358
rect -79999 -24366 -79955 -24358
rect -79899 -24366 -79855 -24358
rect -79799 -24366 -79755 -24358
rect -79699 -24366 -79655 -24358
rect -79599 -24366 -79555 -24358
rect -79499 -24366 -79455 -24358
rect -79399 -24366 -79355 -24358
rect -79299 -24366 -79255 -24358
rect -78799 -24366 -78755 -24358
rect -78699 -24366 -78655 -24358
rect -78599 -24366 -78555 -24358
rect -78499 -24366 -78455 -24358
rect -78399 -24366 -78355 -24358
rect -78299 -24366 -78255 -24358
rect -78199 -24366 -78155 -24358
rect -78099 -24366 -78055 -24358
rect -77999 -24366 -77955 -24358
rect -77899 -24366 -77855 -24358
rect -77799 -24366 -77755 -24358
rect -77699 -24366 -77655 -24358
rect -77599 -24366 -77555 -24358
rect -77499 -24366 -77455 -24358
rect -77399 -24366 -77355 -24358
rect -77299 -24366 -77255 -24358
rect -76799 -24366 -76755 -24358
rect -76699 -24366 -76655 -24358
rect -76599 -24366 -76555 -24358
rect -76499 -24366 -76455 -24358
rect -76399 -24366 -76355 -24358
rect -76299 -24366 -76255 -24358
rect -76199 -24366 -76155 -24358
rect -76099 -24366 -76055 -24358
rect -75999 -24366 -75955 -24358
rect -75899 -24366 -75855 -24358
rect -75799 -24366 -75755 -24358
rect -75699 -24366 -75655 -24358
rect -75599 -24366 -75555 -24358
rect -75499 -24366 -75455 -24358
rect -75399 -24366 -75355 -24358
rect -75299 -24366 -75255 -24358
rect -82755 -24410 -82747 -24366
rect -82655 -24410 -82647 -24366
rect -82555 -24410 -82547 -24366
rect -82455 -24410 -82447 -24366
rect -82355 -24410 -82347 -24366
rect -82255 -24410 -82247 -24366
rect -82155 -24410 -82147 -24366
rect -82055 -24410 -82047 -24366
rect -81955 -24410 -81947 -24366
rect -81855 -24410 -81847 -24366
rect -81755 -24410 -81747 -24366
rect -81655 -24410 -81647 -24366
rect -81555 -24410 -81547 -24366
rect -81455 -24410 -81447 -24366
rect -81355 -24410 -81347 -24366
rect -81255 -24410 -81247 -24366
rect -80755 -24410 -80747 -24366
rect -80655 -24410 -80647 -24366
rect -80555 -24410 -80547 -24366
rect -80455 -24410 -80447 -24366
rect -80355 -24410 -80347 -24366
rect -80255 -24410 -80247 -24366
rect -80155 -24410 -80147 -24366
rect -80055 -24410 -80047 -24366
rect -79955 -24410 -79947 -24366
rect -79855 -24410 -79847 -24366
rect -79755 -24410 -79747 -24366
rect -79655 -24410 -79647 -24366
rect -79555 -24410 -79547 -24366
rect -79455 -24410 -79447 -24366
rect -79355 -24410 -79347 -24366
rect -79255 -24410 -79247 -24366
rect -78755 -24410 -78747 -24366
rect -78655 -24410 -78647 -24366
rect -78555 -24410 -78547 -24366
rect -78455 -24410 -78447 -24366
rect -78355 -24410 -78347 -24366
rect -78255 -24410 -78247 -24366
rect -78155 -24410 -78147 -24366
rect -78055 -24410 -78047 -24366
rect -77955 -24410 -77947 -24366
rect -77855 -24410 -77847 -24366
rect -77755 -24410 -77747 -24366
rect -77655 -24410 -77647 -24366
rect -77555 -24410 -77547 -24366
rect -77455 -24410 -77447 -24366
rect -77355 -24410 -77347 -24366
rect -77255 -24410 -77247 -24366
rect -76755 -24410 -76747 -24366
rect -76655 -24410 -76647 -24366
rect -76555 -24410 -76547 -24366
rect -76455 -24410 -76447 -24366
rect -76355 -24410 -76347 -24366
rect -76255 -24410 -76247 -24366
rect -76155 -24410 -76147 -24366
rect -76055 -24410 -76047 -24366
rect -75955 -24410 -75947 -24366
rect -75855 -24410 -75847 -24366
rect -75755 -24410 -75747 -24366
rect -75655 -24410 -75647 -24366
rect -75555 -24410 -75547 -24366
rect -75455 -24410 -75447 -24366
rect -75355 -24410 -75347 -24366
rect -75255 -24410 -75247 -24366
rect -82799 -24466 -82755 -24458
rect -82699 -24466 -82655 -24458
rect -82599 -24466 -82555 -24458
rect -82499 -24466 -82455 -24458
rect -82399 -24466 -82355 -24458
rect -82299 -24466 -82255 -24458
rect -82199 -24466 -82155 -24458
rect -82099 -24466 -82055 -24458
rect -81999 -24466 -81955 -24458
rect -81899 -24466 -81855 -24458
rect -81799 -24466 -81755 -24458
rect -81699 -24466 -81655 -24458
rect -81599 -24466 -81555 -24458
rect -81499 -24466 -81455 -24458
rect -81399 -24466 -81355 -24458
rect -81299 -24466 -81255 -24458
rect -80799 -24466 -80755 -24458
rect -80699 -24466 -80655 -24458
rect -80599 -24466 -80555 -24458
rect -80499 -24466 -80455 -24458
rect -80399 -24466 -80355 -24458
rect -80299 -24466 -80255 -24458
rect -80199 -24466 -80155 -24458
rect -80099 -24466 -80055 -24458
rect -79999 -24466 -79955 -24458
rect -79899 -24466 -79855 -24458
rect -79799 -24466 -79755 -24458
rect -79699 -24466 -79655 -24458
rect -79599 -24466 -79555 -24458
rect -79499 -24466 -79455 -24458
rect -79399 -24466 -79355 -24458
rect -79299 -24466 -79255 -24458
rect -78799 -24466 -78755 -24458
rect -78699 -24466 -78655 -24458
rect -78599 -24466 -78555 -24458
rect -78499 -24466 -78455 -24458
rect -78399 -24466 -78355 -24458
rect -78299 -24466 -78255 -24458
rect -78199 -24466 -78155 -24458
rect -78099 -24466 -78055 -24458
rect -77999 -24466 -77955 -24458
rect -77899 -24466 -77855 -24458
rect -77799 -24466 -77755 -24458
rect -77699 -24466 -77655 -24458
rect -77599 -24466 -77555 -24458
rect -77499 -24466 -77455 -24458
rect -77399 -24466 -77355 -24458
rect -77299 -24466 -77255 -24458
rect -76799 -24466 -76755 -24458
rect -76699 -24466 -76655 -24458
rect -76599 -24466 -76555 -24458
rect -76499 -24466 -76455 -24458
rect -76399 -24466 -76355 -24458
rect -76299 -24466 -76255 -24458
rect -76199 -24466 -76155 -24458
rect -76099 -24466 -76055 -24458
rect -75999 -24466 -75955 -24458
rect -75899 -24466 -75855 -24458
rect -75799 -24466 -75755 -24458
rect -75699 -24466 -75655 -24458
rect -75599 -24466 -75555 -24458
rect -75499 -24466 -75455 -24458
rect -75399 -24466 -75355 -24458
rect -75299 -24466 -75255 -24458
rect -82755 -24510 -82747 -24466
rect -82655 -24510 -82647 -24466
rect -82555 -24510 -82547 -24466
rect -82455 -24510 -82447 -24466
rect -82355 -24510 -82347 -24466
rect -82255 -24510 -82247 -24466
rect -82155 -24510 -82147 -24466
rect -82055 -24510 -82047 -24466
rect -81955 -24510 -81947 -24466
rect -81855 -24510 -81847 -24466
rect -81755 -24510 -81747 -24466
rect -81655 -24510 -81647 -24466
rect -81555 -24510 -81547 -24466
rect -81455 -24510 -81447 -24466
rect -81355 -24510 -81347 -24466
rect -81255 -24510 -81247 -24466
rect -80755 -24510 -80747 -24466
rect -80655 -24510 -80647 -24466
rect -80555 -24510 -80547 -24466
rect -80455 -24510 -80447 -24466
rect -80355 -24510 -80347 -24466
rect -80255 -24510 -80247 -24466
rect -80155 -24510 -80147 -24466
rect -80055 -24510 -80047 -24466
rect -79955 -24510 -79947 -24466
rect -79855 -24510 -79847 -24466
rect -79755 -24510 -79747 -24466
rect -79655 -24510 -79647 -24466
rect -79555 -24510 -79547 -24466
rect -79455 -24510 -79447 -24466
rect -79355 -24510 -79347 -24466
rect -79255 -24510 -79247 -24466
rect -78755 -24510 -78747 -24466
rect -78655 -24510 -78647 -24466
rect -78555 -24510 -78547 -24466
rect -78455 -24510 -78447 -24466
rect -78355 -24510 -78347 -24466
rect -78255 -24510 -78247 -24466
rect -78155 -24510 -78147 -24466
rect -78055 -24510 -78047 -24466
rect -77955 -24510 -77947 -24466
rect -77855 -24510 -77847 -24466
rect -77755 -24510 -77747 -24466
rect -77655 -24510 -77647 -24466
rect -77555 -24510 -77547 -24466
rect -77455 -24510 -77447 -24466
rect -77355 -24510 -77347 -24466
rect -77255 -24510 -77247 -24466
rect -76755 -24510 -76747 -24466
rect -76655 -24510 -76647 -24466
rect -76555 -24510 -76547 -24466
rect -76455 -24510 -76447 -24466
rect -76355 -24510 -76347 -24466
rect -76255 -24510 -76247 -24466
rect -76155 -24510 -76147 -24466
rect -76055 -24510 -76047 -24466
rect -75955 -24510 -75947 -24466
rect -75855 -24510 -75847 -24466
rect -75755 -24510 -75747 -24466
rect -75655 -24510 -75647 -24466
rect -75555 -24510 -75547 -24466
rect -75455 -24510 -75447 -24466
rect -75355 -24510 -75347 -24466
rect -75255 -24510 -75247 -24466
rect -82799 -24566 -82755 -24558
rect -82699 -24566 -82655 -24558
rect -82599 -24566 -82555 -24558
rect -82499 -24566 -82455 -24558
rect -82399 -24566 -82355 -24558
rect -82299 -24566 -82255 -24558
rect -82199 -24566 -82155 -24558
rect -82099 -24566 -82055 -24558
rect -81999 -24566 -81955 -24558
rect -81899 -24566 -81855 -24558
rect -81799 -24566 -81755 -24558
rect -81699 -24566 -81655 -24558
rect -81599 -24566 -81555 -24558
rect -81499 -24566 -81455 -24558
rect -81399 -24566 -81355 -24558
rect -81299 -24566 -81255 -24558
rect -80799 -24566 -80755 -24558
rect -80699 -24566 -80655 -24558
rect -80599 -24566 -80555 -24558
rect -80499 -24566 -80455 -24558
rect -80399 -24566 -80355 -24558
rect -80299 -24566 -80255 -24558
rect -80199 -24566 -80155 -24558
rect -80099 -24566 -80055 -24558
rect -79999 -24566 -79955 -24558
rect -79899 -24566 -79855 -24558
rect -79799 -24566 -79755 -24558
rect -79699 -24566 -79655 -24558
rect -79599 -24566 -79555 -24558
rect -79499 -24566 -79455 -24558
rect -79399 -24566 -79355 -24558
rect -79299 -24566 -79255 -24558
rect -78799 -24566 -78755 -24558
rect -78699 -24566 -78655 -24558
rect -78599 -24566 -78555 -24558
rect -78499 -24566 -78455 -24558
rect -78399 -24566 -78355 -24558
rect -78299 -24566 -78255 -24558
rect -78199 -24566 -78155 -24558
rect -78099 -24566 -78055 -24558
rect -77999 -24566 -77955 -24558
rect -77899 -24566 -77855 -24558
rect -77799 -24566 -77755 -24558
rect -77699 -24566 -77655 -24558
rect -77599 -24566 -77555 -24558
rect -77499 -24566 -77455 -24558
rect -77399 -24566 -77355 -24558
rect -77299 -24566 -77255 -24558
rect -76799 -24566 -76755 -24558
rect -76699 -24566 -76655 -24558
rect -76599 -24566 -76555 -24558
rect -76499 -24566 -76455 -24558
rect -76399 -24566 -76355 -24558
rect -76299 -24566 -76255 -24558
rect -76199 -24566 -76155 -24558
rect -76099 -24566 -76055 -24558
rect -75999 -24566 -75955 -24558
rect -75899 -24566 -75855 -24558
rect -75799 -24566 -75755 -24558
rect -75699 -24566 -75655 -24558
rect -75599 -24566 -75555 -24558
rect -75499 -24566 -75455 -24558
rect -75399 -24566 -75355 -24558
rect -75299 -24566 -75255 -24558
rect -82755 -24610 -82747 -24566
rect -82655 -24610 -82647 -24566
rect -82555 -24610 -82547 -24566
rect -82455 -24610 -82447 -24566
rect -82355 -24610 -82347 -24566
rect -82255 -24610 -82247 -24566
rect -82155 -24610 -82147 -24566
rect -82055 -24610 -82047 -24566
rect -81955 -24610 -81947 -24566
rect -81855 -24610 -81847 -24566
rect -81755 -24610 -81747 -24566
rect -81655 -24610 -81647 -24566
rect -81555 -24610 -81547 -24566
rect -81455 -24610 -81447 -24566
rect -81355 -24610 -81347 -24566
rect -81255 -24610 -81247 -24566
rect -80755 -24610 -80747 -24566
rect -80655 -24610 -80647 -24566
rect -80555 -24610 -80547 -24566
rect -80455 -24610 -80447 -24566
rect -80355 -24610 -80347 -24566
rect -80255 -24610 -80247 -24566
rect -80155 -24610 -80147 -24566
rect -80055 -24610 -80047 -24566
rect -79955 -24610 -79947 -24566
rect -79855 -24610 -79847 -24566
rect -79755 -24610 -79747 -24566
rect -79655 -24610 -79647 -24566
rect -79555 -24610 -79547 -24566
rect -79455 -24610 -79447 -24566
rect -79355 -24610 -79347 -24566
rect -79255 -24610 -79247 -24566
rect -78755 -24610 -78747 -24566
rect -78655 -24610 -78647 -24566
rect -78555 -24610 -78547 -24566
rect -78455 -24610 -78447 -24566
rect -78355 -24610 -78347 -24566
rect -78255 -24610 -78247 -24566
rect -78155 -24610 -78147 -24566
rect -78055 -24610 -78047 -24566
rect -77955 -24610 -77947 -24566
rect -77855 -24610 -77847 -24566
rect -77755 -24610 -77747 -24566
rect -77655 -24610 -77647 -24566
rect -77555 -24610 -77547 -24566
rect -77455 -24610 -77447 -24566
rect -77355 -24610 -77347 -24566
rect -77255 -24610 -77247 -24566
rect -76755 -24610 -76747 -24566
rect -76655 -24610 -76647 -24566
rect -76555 -24610 -76547 -24566
rect -76455 -24610 -76447 -24566
rect -76355 -24610 -76347 -24566
rect -76255 -24610 -76247 -24566
rect -76155 -24610 -76147 -24566
rect -76055 -24610 -76047 -24566
rect -75955 -24610 -75947 -24566
rect -75855 -24610 -75847 -24566
rect -75755 -24610 -75747 -24566
rect -75655 -24610 -75647 -24566
rect -75555 -24610 -75547 -24566
rect -75455 -24610 -75447 -24566
rect -75355 -24610 -75347 -24566
rect -75255 -24610 -75247 -24566
rect -82799 -24666 -82755 -24658
rect -82699 -24666 -82655 -24658
rect -82599 -24666 -82555 -24658
rect -82499 -24666 -82455 -24658
rect -82399 -24666 -82355 -24658
rect -82299 -24666 -82255 -24658
rect -82199 -24666 -82155 -24658
rect -82099 -24666 -82055 -24658
rect -81999 -24666 -81955 -24658
rect -81899 -24666 -81855 -24658
rect -81799 -24666 -81755 -24658
rect -81699 -24666 -81655 -24658
rect -81599 -24666 -81555 -24658
rect -81499 -24666 -81455 -24658
rect -81399 -24666 -81355 -24658
rect -81299 -24666 -81255 -24658
rect -80799 -24666 -80755 -24658
rect -80699 -24666 -80655 -24658
rect -80599 -24666 -80555 -24658
rect -80499 -24666 -80455 -24658
rect -80399 -24666 -80355 -24658
rect -80299 -24666 -80255 -24658
rect -80199 -24666 -80155 -24658
rect -80099 -24666 -80055 -24658
rect -79999 -24666 -79955 -24658
rect -79899 -24666 -79855 -24658
rect -79799 -24666 -79755 -24658
rect -79699 -24666 -79655 -24658
rect -79599 -24666 -79555 -24658
rect -79499 -24666 -79455 -24658
rect -79399 -24666 -79355 -24658
rect -79299 -24666 -79255 -24658
rect -78799 -24666 -78755 -24658
rect -78699 -24666 -78655 -24658
rect -78599 -24666 -78555 -24658
rect -78499 -24666 -78455 -24658
rect -78399 -24666 -78355 -24658
rect -78299 -24666 -78255 -24658
rect -78199 -24666 -78155 -24658
rect -78099 -24666 -78055 -24658
rect -77999 -24666 -77955 -24658
rect -77899 -24666 -77855 -24658
rect -77799 -24666 -77755 -24658
rect -77699 -24666 -77655 -24658
rect -77599 -24666 -77555 -24658
rect -77499 -24666 -77455 -24658
rect -77399 -24666 -77355 -24658
rect -77299 -24666 -77255 -24658
rect -76799 -24666 -76755 -24658
rect -76699 -24666 -76655 -24658
rect -76599 -24666 -76555 -24658
rect -76499 -24666 -76455 -24658
rect -76399 -24666 -76355 -24658
rect -76299 -24666 -76255 -24658
rect -76199 -24666 -76155 -24658
rect -76099 -24666 -76055 -24658
rect -75999 -24666 -75955 -24658
rect -75899 -24666 -75855 -24658
rect -75799 -24666 -75755 -24658
rect -75699 -24666 -75655 -24658
rect -75599 -24666 -75555 -24658
rect -75499 -24666 -75455 -24658
rect -75399 -24666 -75355 -24658
rect -75299 -24666 -75255 -24658
rect -82755 -24710 -82747 -24666
rect -82655 -24710 -82647 -24666
rect -82555 -24710 -82547 -24666
rect -82455 -24710 -82447 -24666
rect -82355 -24710 -82347 -24666
rect -82255 -24710 -82247 -24666
rect -82155 -24710 -82147 -24666
rect -82055 -24710 -82047 -24666
rect -81955 -24710 -81947 -24666
rect -81855 -24710 -81847 -24666
rect -81755 -24710 -81747 -24666
rect -81655 -24710 -81647 -24666
rect -81555 -24710 -81547 -24666
rect -81455 -24710 -81447 -24666
rect -81355 -24710 -81347 -24666
rect -81255 -24710 -81247 -24666
rect -80755 -24710 -80747 -24666
rect -80655 -24710 -80647 -24666
rect -80555 -24710 -80547 -24666
rect -80455 -24710 -80447 -24666
rect -80355 -24710 -80347 -24666
rect -80255 -24710 -80247 -24666
rect -80155 -24710 -80147 -24666
rect -80055 -24710 -80047 -24666
rect -79955 -24710 -79947 -24666
rect -79855 -24710 -79847 -24666
rect -79755 -24710 -79747 -24666
rect -79655 -24710 -79647 -24666
rect -79555 -24710 -79547 -24666
rect -79455 -24710 -79447 -24666
rect -79355 -24710 -79347 -24666
rect -79255 -24710 -79247 -24666
rect -78755 -24710 -78747 -24666
rect -78655 -24710 -78647 -24666
rect -78555 -24710 -78547 -24666
rect -78455 -24710 -78447 -24666
rect -78355 -24710 -78347 -24666
rect -78255 -24710 -78247 -24666
rect -78155 -24710 -78147 -24666
rect -78055 -24710 -78047 -24666
rect -77955 -24710 -77947 -24666
rect -77855 -24710 -77847 -24666
rect -77755 -24710 -77747 -24666
rect -77655 -24710 -77647 -24666
rect -77555 -24710 -77547 -24666
rect -77455 -24710 -77447 -24666
rect -77355 -24710 -77347 -24666
rect -77255 -24710 -77247 -24666
rect -76755 -24710 -76747 -24666
rect -76655 -24710 -76647 -24666
rect -76555 -24710 -76547 -24666
rect -76455 -24710 -76447 -24666
rect -76355 -24710 -76347 -24666
rect -76255 -24710 -76247 -24666
rect -76155 -24710 -76147 -24666
rect -76055 -24710 -76047 -24666
rect -75955 -24710 -75947 -24666
rect -75855 -24710 -75847 -24666
rect -75755 -24710 -75747 -24666
rect -75655 -24710 -75647 -24666
rect -75555 -24710 -75547 -24666
rect -75455 -24710 -75447 -24666
rect -75355 -24710 -75347 -24666
rect -75255 -24710 -75247 -24666
rect -82799 -24766 -82755 -24758
rect -82699 -24766 -82655 -24758
rect -82599 -24766 -82555 -24758
rect -82499 -24766 -82455 -24758
rect -82399 -24766 -82355 -24758
rect -82299 -24766 -82255 -24758
rect -82199 -24766 -82155 -24758
rect -82099 -24766 -82055 -24758
rect -81999 -24766 -81955 -24758
rect -81899 -24766 -81855 -24758
rect -81799 -24766 -81755 -24758
rect -81699 -24766 -81655 -24758
rect -81599 -24766 -81555 -24758
rect -81499 -24766 -81455 -24758
rect -81399 -24766 -81355 -24758
rect -81299 -24766 -81255 -24758
rect -80799 -24766 -80755 -24758
rect -80699 -24766 -80655 -24758
rect -80599 -24766 -80555 -24758
rect -80499 -24766 -80455 -24758
rect -80399 -24766 -80355 -24758
rect -80299 -24766 -80255 -24758
rect -80199 -24766 -80155 -24758
rect -80099 -24766 -80055 -24758
rect -79999 -24766 -79955 -24758
rect -79899 -24766 -79855 -24758
rect -79799 -24766 -79755 -24758
rect -79699 -24766 -79655 -24758
rect -79599 -24766 -79555 -24758
rect -79499 -24766 -79455 -24758
rect -79399 -24766 -79355 -24758
rect -79299 -24766 -79255 -24758
rect -78799 -24766 -78755 -24758
rect -78699 -24766 -78655 -24758
rect -78599 -24766 -78555 -24758
rect -78499 -24766 -78455 -24758
rect -78399 -24766 -78355 -24758
rect -78299 -24766 -78255 -24758
rect -78199 -24766 -78155 -24758
rect -78099 -24766 -78055 -24758
rect -77999 -24766 -77955 -24758
rect -77899 -24766 -77855 -24758
rect -77799 -24766 -77755 -24758
rect -77699 -24766 -77655 -24758
rect -77599 -24766 -77555 -24758
rect -77499 -24766 -77455 -24758
rect -77399 -24766 -77355 -24758
rect -77299 -24766 -77255 -24758
rect -76799 -24766 -76755 -24758
rect -76699 -24766 -76655 -24758
rect -76599 -24766 -76555 -24758
rect -76499 -24766 -76455 -24758
rect -76399 -24766 -76355 -24758
rect -76299 -24766 -76255 -24758
rect -76199 -24766 -76155 -24758
rect -76099 -24766 -76055 -24758
rect -75999 -24766 -75955 -24758
rect -75899 -24766 -75855 -24758
rect -75799 -24766 -75755 -24758
rect -75699 -24766 -75655 -24758
rect -75599 -24766 -75555 -24758
rect -75499 -24766 -75455 -24758
rect -75399 -24766 -75355 -24758
rect -75299 -24766 -75255 -24758
rect -82755 -24810 -82747 -24766
rect -82655 -24810 -82647 -24766
rect -82555 -24810 -82547 -24766
rect -82455 -24810 -82447 -24766
rect -82355 -24810 -82347 -24766
rect -82255 -24810 -82247 -24766
rect -82155 -24810 -82147 -24766
rect -82055 -24810 -82047 -24766
rect -81955 -24810 -81947 -24766
rect -81855 -24810 -81847 -24766
rect -81755 -24810 -81747 -24766
rect -81655 -24810 -81647 -24766
rect -81555 -24810 -81547 -24766
rect -81455 -24810 -81447 -24766
rect -81355 -24810 -81347 -24766
rect -81255 -24810 -81247 -24766
rect -80755 -24810 -80747 -24766
rect -80655 -24810 -80647 -24766
rect -80555 -24810 -80547 -24766
rect -80455 -24810 -80447 -24766
rect -80355 -24810 -80347 -24766
rect -80255 -24810 -80247 -24766
rect -80155 -24810 -80147 -24766
rect -80055 -24810 -80047 -24766
rect -79955 -24810 -79947 -24766
rect -79855 -24810 -79847 -24766
rect -79755 -24810 -79747 -24766
rect -79655 -24810 -79647 -24766
rect -79555 -24810 -79547 -24766
rect -79455 -24810 -79447 -24766
rect -79355 -24810 -79347 -24766
rect -79255 -24810 -79247 -24766
rect -78755 -24810 -78747 -24766
rect -78655 -24810 -78647 -24766
rect -78555 -24810 -78547 -24766
rect -78455 -24810 -78447 -24766
rect -78355 -24810 -78347 -24766
rect -78255 -24810 -78247 -24766
rect -78155 -24810 -78147 -24766
rect -78055 -24810 -78047 -24766
rect -77955 -24810 -77947 -24766
rect -77855 -24810 -77847 -24766
rect -77755 -24810 -77747 -24766
rect -77655 -24810 -77647 -24766
rect -77555 -24810 -77547 -24766
rect -77455 -24810 -77447 -24766
rect -77355 -24810 -77347 -24766
rect -77255 -24810 -77247 -24766
rect -76755 -24810 -76747 -24766
rect -76655 -24810 -76647 -24766
rect -76555 -24810 -76547 -24766
rect -76455 -24810 -76447 -24766
rect -76355 -24810 -76347 -24766
rect -76255 -24810 -76247 -24766
rect -76155 -24810 -76147 -24766
rect -76055 -24810 -76047 -24766
rect -75955 -24810 -75947 -24766
rect -75855 -24810 -75847 -24766
rect -75755 -24810 -75747 -24766
rect -75655 -24810 -75647 -24766
rect -75555 -24810 -75547 -24766
rect -75455 -24810 -75447 -24766
rect -75355 -24810 -75347 -24766
rect -75255 -24810 -75247 -24766
rect -82799 -24866 -82755 -24858
rect -82699 -24866 -82655 -24858
rect -82599 -24866 -82555 -24858
rect -82499 -24866 -82455 -24858
rect -82399 -24866 -82355 -24858
rect -82299 -24866 -82255 -24858
rect -82199 -24866 -82155 -24858
rect -82099 -24866 -82055 -24858
rect -81999 -24866 -81955 -24858
rect -81899 -24866 -81855 -24858
rect -81799 -24866 -81755 -24858
rect -81699 -24866 -81655 -24858
rect -81599 -24866 -81555 -24858
rect -81499 -24866 -81455 -24858
rect -81399 -24866 -81355 -24858
rect -81299 -24866 -81255 -24858
rect -80799 -24866 -80755 -24858
rect -80699 -24866 -80655 -24858
rect -80599 -24866 -80555 -24858
rect -80499 -24866 -80455 -24858
rect -80399 -24866 -80355 -24858
rect -80299 -24866 -80255 -24858
rect -80199 -24866 -80155 -24858
rect -80099 -24866 -80055 -24858
rect -79999 -24866 -79955 -24858
rect -79899 -24866 -79855 -24858
rect -79799 -24866 -79755 -24858
rect -79699 -24866 -79655 -24858
rect -79599 -24866 -79555 -24858
rect -79499 -24866 -79455 -24858
rect -79399 -24866 -79355 -24858
rect -79299 -24866 -79255 -24858
rect -78799 -24866 -78755 -24858
rect -78699 -24866 -78655 -24858
rect -78599 -24866 -78555 -24858
rect -78499 -24866 -78455 -24858
rect -78399 -24866 -78355 -24858
rect -78299 -24866 -78255 -24858
rect -78199 -24866 -78155 -24858
rect -78099 -24866 -78055 -24858
rect -77999 -24866 -77955 -24858
rect -77899 -24866 -77855 -24858
rect -77799 -24866 -77755 -24858
rect -77699 -24866 -77655 -24858
rect -77599 -24866 -77555 -24858
rect -77499 -24866 -77455 -24858
rect -77399 -24866 -77355 -24858
rect -77299 -24866 -77255 -24858
rect -76799 -24866 -76755 -24858
rect -76699 -24866 -76655 -24858
rect -76599 -24866 -76555 -24858
rect -76499 -24866 -76455 -24858
rect -76399 -24866 -76355 -24858
rect -76299 -24866 -76255 -24858
rect -76199 -24866 -76155 -24858
rect -76099 -24866 -76055 -24858
rect -75999 -24866 -75955 -24858
rect -75899 -24866 -75855 -24858
rect -75799 -24866 -75755 -24858
rect -75699 -24866 -75655 -24858
rect -75599 -24866 -75555 -24858
rect -75499 -24866 -75455 -24858
rect -75399 -24866 -75355 -24858
rect -75299 -24866 -75255 -24858
rect -82755 -24910 -82747 -24866
rect -82655 -24910 -82647 -24866
rect -82555 -24910 -82547 -24866
rect -82455 -24910 -82447 -24866
rect -82355 -24910 -82347 -24866
rect -82255 -24910 -82247 -24866
rect -82155 -24910 -82147 -24866
rect -82055 -24910 -82047 -24866
rect -81955 -24910 -81947 -24866
rect -81855 -24910 -81847 -24866
rect -81755 -24910 -81747 -24866
rect -81655 -24910 -81647 -24866
rect -81555 -24910 -81547 -24866
rect -81455 -24910 -81447 -24866
rect -81355 -24910 -81347 -24866
rect -81255 -24910 -81247 -24866
rect -80755 -24910 -80747 -24866
rect -80655 -24910 -80647 -24866
rect -80555 -24910 -80547 -24866
rect -80455 -24910 -80447 -24866
rect -80355 -24910 -80347 -24866
rect -80255 -24910 -80247 -24866
rect -80155 -24910 -80147 -24866
rect -80055 -24910 -80047 -24866
rect -79955 -24910 -79947 -24866
rect -79855 -24910 -79847 -24866
rect -79755 -24910 -79747 -24866
rect -79655 -24910 -79647 -24866
rect -79555 -24910 -79547 -24866
rect -79455 -24910 -79447 -24866
rect -79355 -24910 -79347 -24866
rect -79255 -24910 -79247 -24866
rect -78755 -24910 -78747 -24866
rect -78655 -24910 -78647 -24866
rect -78555 -24910 -78547 -24866
rect -78455 -24910 -78447 -24866
rect -78355 -24910 -78347 -24866
rect -78255 -24910 -78247 -24866
rect -78155 -24910 -78147 -24866
rect -78055 -24910 -78047 -24866
rect -77955 -24910 -77947 -24866
rect -77855 -24910 -77847 -24866
rect -77755 -24910 -77747 -24866
rect -77655 -24910 -77647 -24866
rect -77555 -24910 -77547 -24866
rect -77455 -24910 -77447 -24866
rect -77355 -24910 -77347 -24866
rect -77255 -24910 -77247 -24866
rect -76755 -24910 -76747 -24866
rect -76655 -24910 -76647 -24866
rect -76555 -24910 -76547 -24866
rect -76455 -24910 -76447 -24866
rect -76355 -24910 -76347 -24866
rect -76255 -24910 -76247 -24866
rect -76155 -24910 -76147 -24866
rect -76055 -24910 -76047 -24866
rect -75955 -24910 -75947 -24866
rect -75855 -24910 -75847 -24866
rect -75755 -24910 -75747 -24866
rect -75655 -24910 -75647 -24866
rect -75555 -24910 -75547 -24866
rect -75455 -24910 -75447 -24866
rect -75355 -24910 -75347 -24866
rect -75255 -24910 -75247 -24866
rect -82799 -24966 -82755 -24958
rect -82699 -24966 -82655 -24958
rect -82599 -24966 -82555 -24958
rect -82499 -24966 -82455 -24958
rect -82399 -24966 -82355 -24958
rect -82299 -24966 -82255 -24958
rect -82199 -24966 -82155 -24958
rect -82099 -24966 -82055 -24958
rect -81999 -24966 -81955 -24958
rect -81899 -24966 -81855 -24958
rect -81799 -24966 -81755 -24958
rect -81699 -24966 -81655 -24958
rect -81599 -24966 -81555 -24958
rect -81499 -24966 -81455 -24958
rect -81399 -24966 -81355 -24958
rect -81299 -24966 -81255 -24958
rect -80799 -24966 -80755 -24958
rect -80699 -24966 -80655 -24958
rect -80599 -24966 -80555 -24958
rect -80499 -24966 -80455 -24958
rect -80399 -24966 -80355 -24958
rect -80299 -24966 -80255 -24958
rect -80199 -24966 -80155 -24958
rect -80099 -24966 -80055 -24958
rect -79999 -24966 -79955 -24958
rect -79899 -24966 -79855 -24958
rect -79799 -24966 -79755 -24958
rect -79699 -24966 -79655 -24958
rect -79599 -24966 -79555 -24958
rect -79499 -24966 -79455 -24958
rect -79399 -24966 -79355 -24958
rect -79299 -24966 -79255 -24958
rect -78799 -24966 -78755 -24958
rect -78699 -24966 -78655 -24958
rect -78599 -24966 -78555 -24958
rect -78499 -24966 -78455 -24958
rect -78399 -24966 -78355 -24958
rect -78299 -24966 -78255 -24958
rect -78199 -24966 -78155 -24958
rect -78099 -24966 -78055 -24958
rect -77999 -24966 -77955 -24958
rect -77899 -24966 -77855 -24958
rect -77799 -24966 -77755 -24958
rect -77699 -24966 -77655 -24958
rect -77599 -24966 -77555 -24958
rect -77499 -24966 -77455 -24958
rect -77399 -24966 -77355 -24958
rect -77299 -24966 -77255 -24958
rect -76799 -24966 -76755 -24958
rect -76699 -24966 -76655 -24958
rect -76599 -24966 -76555 -24958
rect -76499 -24966 -76455 -24958
rect -76399 -24966 -76355 -24958
rect -76299 -24966 -76255 -24958
rect -76199 -24966 -76155 -24958
rect -76099 -24966 -76055 -24958
rect -75999 -24966 -75955 -24958
rect -75899 -24966 -75855 -24958
rect -75799 -24966 -75755 -24958
rect -75699 -24966 -75655 -24958
rect -75599 -24966 -75555 -24958
rect -75499 -24966 -75455 -24958
rect -75399 -24966 -75355 -24958
rect -75299 -24966 -75255 -24958
rect -82755 -25010 -82747 -24966
rect -82655 -25010 -82647 -24966
rect -82555 -25010 -82547 -24966
rect -82455 -25010 -82447 -24966
rect -82355 -25010 -82347 -24966
rect -82255 -25010 -82247 -24966
rect -82155 -25010 -82147 -24966
rect -82055 -25010 -82047 -24966
rect -81955 -25010 -81947 -24966
rect -81855 -25010 -81847 -24966
rect -81755 -25010 -81747 -24966
rect -81655 -25010 -81647 -24966
rect -81555 -25010 -81547 -24966
rect -81455 -25010 -81447 -24966
rect -81355 -25010 -81347 -24966
rect -81255 -25010 -81247 -24966
rect -80755 -25010 -80747 -24966
rect -80655 -25010 -80647 -24966
rect -80555 -25010 -80547 -24966
rect -80455 -25010 -80447 -24966
rect -80355 -25010 -80347 -24966
rect -80255 -25010 -80247 -24966
rect -80155 -25010 -80147 -24966
rect -80055 -25010 -80047 -24966
rect -79955 -25010 -79947 -24966
rect -79855 -25010 -79847 -24966
rect -79755 -25010 -79747 -24966
rect -79655 -25010 -79647 -24966
rect -79555 -25010 -79547 -24966
rect -79455 -25010 -79447 -24966
rect -79355 -25010 -79347 -24966
rect -79255 -25010 -79247 -24966
rect -78755 -25010 -78747 -24966
rect -78655 -25010 -78647 -24966
rect -78555 -25010 -78547 -24966
rect -78455 -25010 -78447 -24966
rect -78355 -25010 -78347 -24966
rect -78255 -25010 -78247 -24966
rect -78155 -25010 -78147 -24966
rect -78055 -25010 -78047 -24966
rect -77955 -25010 -77947 -24966
rect -77855 -25010 -77847 -24966
rect -77755 -25010 -77747 -24966
rect -77655 -25010 -77647 -24966
rect -77555 -25010 -77547 -24966
rect -77455 -25010 -77447 -24966
rect -77355 -25010 -77347 -24966
rect -77255 -25010 -77247 -24966
rect -76755 -25010 -76747 -24966
rect -76655 -25010 -76647 -24966
rect -76555 -25010 -76547 -24966
rect -76455 -25010 -76447 -24966
rect -76355 -25010 -76347 -24966
rect -76255 -25010 -76247 -24966
rect -76155 -25010 -76147 -24966
rect -76055 -25010 -76047 -24966
rect -75955 -25010 -75947 -24966
rect -75855 -25010 -75847 -24966
rect -75755 -25010 -75747 -24966
rect -75655 -25010 -75647 -24966
rect -75555 -25010 -75547 -24966
rect -75455 -25010 -75447 -24966
rect -75355 -25010 -75347 -24966
rect -75255 -25010 -75247 -24966
rect -82799 -25066 -82755 -25058
rect -82699 -25066 -82655 -25058
rect -82599 -25066 -82555 -25058
rect -82499 -25066 -82455 -25058
rect -82399 -25066 -82355 -25058
rect -82299 -25066 -82255 -25058
rect -82199 -25066 -82155 -25058
rect -82099 -25066 -82055 -25058
rect -81999 -25066 -81955 -25058
rect -81899 -25066 -81855 -25058
rect -81799 -25066 -81755 -25058
rect -81699 -25066 -81655 -25058
rect -81599 -25066 -81555 -25058
rect -81499 -25066 -81455 -25058
rect -81399 -25066 -81355 -25058
rect -81299 -25066 -81255 -25058
rect -80799 -25066 -80755 -25058
rect -80699 -25066 -80655 -25058
rect -80599 -25066 -80555 -25058
rect -80499 -25066 -80455 -25058
rect -80399 -25066 -80355 -25058
rect -80299 -25066 -80255 -25058
rect -80199 -25066 -80155 -25058
rect -80099 -25066 -80055 -25058
rect -79999 -25066 -79955 -25058
rect -79899 -25066 -79855 -25058
rect -79799 -25066 -79755 -25058
rect -79699 -25066 -79655 -25058
rect -79599 -25066 -79555 -25058
rect -79499 -25066 -79455 -25058
rect -79399 -25066 -79355 -25058
rect -79299 -25066 -79255 -25058
rect -78799 -25066 -78755 -25058
rect -78699 -25066 -78655 -25058
rect -78599 -25066 -78555 -25058
rect -78499 -25066 -78455 -25058
rect -78399 -25066 -78355 -25058
rect -78299 -25066 -78255 -25058
rect -78199 -25066 -78155 -25058
rect -78099 -25066 -78055 -25058
rect -77999 -25066 -77955 -25058
rect -77899 -25066 -77855 -25058
rect -77799 -25066 -77755 -25058
rect -77699 -25066 -77655 -25058
rect -77599 -25066 -77555 -25058
rect -77499 -25066 -77455 -25058
rect -77399 -25066 -77355 -25058
rect -77299 -25066 -77255 -25058
rect -76799 -25066 -76755 -25058
rect -76699 -25066 -76655 -25058
rect -76599 -25066 -76555 -25058
rect -76499 -25066 -76455 -25058
rect -76399 -25066 -76355 -25058
rect -76299 -25066 -76255 -25058
rect -76199 -25066 -76155 -25058
rect -76099 -25066 -76055 -25058
rect -75999 -25066 -75955 -25058
rect -75899 -25066 -75855 -25058
rect -75799 -25066 -75755 -25058
rect -75699 -25066 -75655 -25058
rect -75599 -25066 -75555 -25058
rect -75499 -25066 -75455 -25058
rect -75399 -25066 -75355 -25058
rect -75299 -25066 -75255 -25058
rect -82755 -25110 -82747 -25066
rect -82655 -25110 -82647 -25066
rect -82555 -25110 -82547 -25066
rect -82455 -25110 -82447 -25066
rect -82355 -25110 -82347 -25066
rect -82255 -25110 -82247 -25066
rect -82155 -25110 -82147 -25066
rect -82055 -25110 -82047 -25066
rect -81955 -25110 -81947 -25066
rect -81855 -25110 -81847 -25066
rect -81755 -25110 -81747 -25066
rect -81655 -25110 -81647 -25066
rect -81555 -25110 -81547 -25066
rect -81455 -25110 -81447 -25066
rect -81355 -25110 -81347 -25066
rect -81255 -25110 -81247 -25066
rect -80755 -25110 -80747 -25066
rect -80655 -25110 -80647 -25066
rect -80555 -25110 -80547 -25066
rect -80455 -25110 -80447 -25066
rect -80355 -25110 -80347 -25066
rect -80255 -25110 -80247 -25066
rect -80155 -25110 -80147 -25066
rect -80055 -25110 -80047 -25066
rect -79955 -25110 -79947 -25066
rect -79855 -25110 -79847 -25066
rect -79755 -25110 -79747 -25066
rect -79655 -25110 -79647 -25066
rect -79555 -25110 -79547 -25066
rect -79455 -25110 -79447 -25066
rect -79355 -25110 -79347 -25066
rect -79255 -25110 -79247 -25066
rect -78755 -25110 -78747 -25066
rect -78655 -25110 -78647 -25066
rect -78555 -25110 -78547 -25066
rect -78455 -25110 -78447 -25066
rect -78355 -25110 -78347 -25066
rect -78255 -25110 -78247 -25066
rect -78155 -25110 -78147 -25066
rect -78055 -25110 -78047 -25066
rect -77955 -25110 -77947 -25066
rect -77855 -25110 -77847 -25066
rect -77755 -25110 -77747 -25066
rect -77655 -25110 -77647 -25066
rect -77555 -25110 -77547 -25066
rect -77455 -25110 -77447 -25066
rect -77355 -25110 -77347 -25066
rect -77255 -25110 -77247 -25066
rect -76755 -25110 -76747 -25066
rect -76655 -25110 -76647 -25066
rect -76555 -25110 -76547 -25066
rect -76455 -25110 -76447 -25066
rect -76355 -25110 -76347 -25066
rect -76255 -25110 -76247 -25066
rect -76155 -25110 -76147 -25066
rect -76055 -25110 -76047 -25066
rect -75955 -25110 -75947 -25066
rect -75855 -25110 -75847 -25066
rect -75755 -25110 -75747 -25066
rect -75655 -25110 -75647 -25066
rect -75555 -25110 -75547 -25066
rect -75455 -25110 -75447 -25066
rect -75355 -25110 -75347 -25066
rect -75255 -25110 -75247 -25066
rect -82799 -25166 -82755 -25158
rect -82699 -25166 -82655 -25158
rect -82599 -25166 -82555 -25158
rect -82499 -25166 -82455 -25158
rect -82399 -25166 -82355 -25158
rect -82299 -25166 -82255 -25158
rect -82199 -25166 -82155 -25158
rect -82099 -25166 -82055 -25158
rect -81999 -25166 -81955 -25158
rect -81899 -25166 -81855 -25158
rect -81799 -25166 -81755 -25158
rect -81699 -25166 -81655 -25158
rect -81599 -25166 -81555 -25158
rect -81499 -25166 -81455 -25158
rect -81399 -25166 -81355 -25158
rect -81299 -25166 -81255 -25158
rect -80799 -25166 -80755 -25158
rect -80699 -25166 -80655 -25158
rect -80599 -25166 -80555 -25158
rect -80499 -25166 -80455 -25158
rect -80399 -25166 -80355 -25158
rect -80299 -25166 -80255 -25158
rect -80199 -25166 -80155 -25158
rect -80099 -25166 -80055 -25158
rect -79999 -25166 -79955 -25158
rect -79899 -25166 -79855 -25158
rect -79799 -25166 -79755 -25158
rect -79699 -25166 -79655 -25158
rect -79599 -25166 -79555 -25158
rect -79499 -25166 -79455 -25158
rect -79399 -25166 -79355 -25158
rect -79299 -25166 -79255 -25158
rect -78799 -25166 -78755 -25158
rect -78699 -25166 -78655 -25158
rect -78599 -25166 -78555 -25158
rect -78499 -25166 -78455 -25158
rect -78399 -25166 -78355 -25158
rect -78299 -25166 -78255 -25158
rect -78199 -25166 -78155 -25158
rect -78099 -25166 -78055 -25158
rect -77999 -25166 -77955 -25158
rect -77899 -25166 -77855 -25158
rect -77799 -25166 -77755 -25158
rect -77699 -25166 -77655 -25158
rect -77599 -25166 -77555 -25158
rect -77499 -25166 -77455 -25158
rect -77399 -25166 -77355 -25158
rect -77299 -25166 -77255 -25158
rect -76799 -25166 -76755 -25158
rect -76699 -25166 -76655 -25158
rect -76599 -25166 -76555 -25158
rect -76499 -25166 -76455 -25158
rect -76399 -25166 -76355 -25158
rect -76299 -25166 -76255 -25158
rect -76199 -25166 -76155 -25158
rect -76099 -25166 -76055 -25158
rect -75999 -25166 -75955 -25158
rect -75899 -25166 -75855 -25158
rect -75799 -25166 -75755 -25158
rect -75699 -25166 -75655 -25158
rect -75599 -25166 -75555 -25158
rect -75499 -25166 -75455 -25158
rect -75399 -25166 -75355 -25158
rect -75299 -25166 -75255 -25158
rect -82755 -25210 -82747 -25166
rect -82655 -25210 -82647 -25166
rect -82555 -25210 -82547 -25166
rect -82455 -25210 -82447 -25166
rect -82355 -25210 -82347 -25166
rect -82255 -25210 -82247 -25166
rect -82155 -25210 -82147 -25166
rect -82055 -25210 -82047 -25166
rect -81955 -25210 -81947 -25166
rect -81855 -25210 -81847 -25166
rect -81755 -25210 -81747 -25166
rect -81655 -25210 -81647 -25166
rect -81555 -25210 -81547 -25166
rect -81455 -25210 -81447 -25166
rect -81355 -25210 -81347 -25166
rect -81255 -25210 -81247 -25166
rect -80755 -25210 -80747 -25166
rect -80655 -25210 -80647 -25166
rect -80555 -25210 -80547 -25166
rect -80455 -25210 -80447 -25166
rect -80355 -25210 -80347 -25166
rect -80255 -25210 -80247 -25166
rect -80155 -25210 -80147 -25166
rect -80055 -25210 -80047 -25166
rect -79955 -25210 -79947 -25166
rect -79855 -25210 -79847 -25166
rect -79755 -25210 -79747 -25166
rect -79655 -25210 -79647 -25166
rect -79555 -25210 -79547 -25166
rect -79455 -25210 -79447 -25166
rect -79355 -25210 -79347 -25166
rect -79255 -25210 -79247 -25166
rect -78755 -25210 -78747 -25166
rect -78655 -25210 -78647 -25166
rect -78555 -25210 -78547 -25166
rect -78455 -25210 -78447 -25166
rect -78355 -25210 -78347 -25166
rect -78255 -25210 -78247 -25166
rect -78155 -25210 -78147 -25166
rect -78055 -25210 -78047 -25166
rect -77955 -25210 -77947 -25166
rect -77855 -25210 -77847 -25166
rect -77755 -25210 -77747 -25166
rect -77655 -25210 -77647 -25166
rect -77555 -25210 -77547 -25166
rect -77455 -25210 -77447 -25166
rect -77355 -25210 -77347 -25166
rect -77255 -25210 -77247 -25166
rect -76755 -25210 -76747 -25166
rect -76655 -25210 -76647 -25166
rect -76555 -25210 -76547 -25166
rect -76455 -25210 -76447 -25166
rect -76355 -25210 -76347 -25166
rect -76255 -25210 -76247 -25166
rect -76155 -25210 -76147 -25166
rect -76055 -25210 -76047 -25166
rect -75955 -25210 -75947 -25166
rect -75855 -25210 -75847 -25166
rect -75755 -25210 -75747 -25166
rect -75655 -25210 -75647 -25166
rect -75555 -25210 -75547 -25166
rect -75455 -25210 -75447 -25166
rect -75355 -25210 -75347 -25166
rect -75255 -25210 -75247 -25166
rect -82799 -25266 -82755 -25258
rect -82699 -25266 -82655 -25258
rect -82599 -25266 -82555 -25258
rect -82499 -25266 -82455 -25258
rect -82399 -25266 -82355 -25258
rect -82299 -25266 -82255 -25258
rect -82199 -25266 -82155 -25258
rect -82099 -25266 -82055 -25258
rect -81999 -25266 -81955 -25258
rect -81899 -25266 -81855 -25258
rect -81799 -25266 -81755 -25258
rect -81699 -25266 -81655 -25258
rect -81599 -25266 -81555 -25258
rect -81499 -25266 -81455 -25258
rect -81399 -25266 -81355 -25258
rect -81299 -25266 -81255 -25258
rect -80799 -25266 -80755 -25258
rect -80699 -25266 -80655 -25258
rect -80599 -25266 -80555 -25258
rect -80499 -25266 -80455 -25258
rect -80399 -25266 -80355 -25258
rect -80299 -25266 -80255 -25258
rect -80199 -25266 -80155 -25258
rect -80099 -25266 -80055 -25258
rect -79999 -25266 -79955 -25258
rect -79899 -25266 -79855 -25258
rect -79799 -25266 -79755 -25258
rect -79699 -25266 -79655 -25258
rect -79599 -25266 -79555 -25258
rect -79499 -25266 -79455 -25258
rect -79399 -25266 -79355 -25258
rect -79299 -25266 -79255 -25258
rect -78799 -25266 -78755 -25258
rect -78699 -25266 -78655 -25258
rect -78599 -25266 -78555 -25258
rect -78499 -25266 -78455 -25258
rect -78399 -25266 -78355 -25258
rect -78299 -25266 -78255 -25258
rect -78199 -25266 -78155 -25258
rect -78099 -25266 -78055 -25258
rect -77999 -25266 -77955 -25258
rect -77899 -25266 -77855 -25258
rect -77799 -25266 -77755 -25258
rect -77699 -25266 -77655 -25258
rect -77599 -25266 -77555 -25258
rect -77499 -25266 -77455 -25258
rect -77399 -25266 -77355 -25258
rect -77299 -25266 -77255 -25258
rect -76799 -25266 -76755 -25258
rect -76699 -25266 -76655 -25258
rect -76599 -25266 -76555 -25258
rect -76499 -25266 -76455 -25258
rect -76399 -25266 -76355 -25258
rect -76299 -25266 -76255 -25258
rect -76199 -25266 -76155 -25258
rect -76099 -25266 -76055 -25258
rect -75999 -25266 -75955 -25258
rect -75899 -25266 -75855 -25258
rect -75799 -25266 -75755 -25258
rect -75699 -25266 -75655 -25258
rect -75599 -25266 -75555 -25258
rect -75499 -25266 -75455 -25258
rect -75399 -25266 -75355 -25258
rect -75299 -25266 -75255 -25258
rect -82755 -25310 -82747 -25266
rect -82655 -25310 -82647 -25266
rect -82555 -25310 -82547 -25266
rect -82455 -25310 -82447 -25266
rect -82355 -25310 -82347 -25266
rect -82255 -25310 -82247 -25266
rect -82155 -25310 -82147 -25266
rect -82055 -25310 -82047 -25266
rect -81955 -25310 -81947 -25266
rect -81855 -25310 -81847 -25266
rect -81755 -25310 -81747 -25266
rect -81655 -25310 -81647 -25266
rect -81555 -25310 -81547 -25266
rect -81455 -25310 -81447 -25266
rect -81355 -25310 -81347 -25266
rect -81255 -25310 -81247 -25266
rect -80755 -25310 -80747 -25266
rect -80655 -25310 -80647 -25266
rect -80555 -25310 -80547 -25266
rect -80455 -25310 -80447 -25266
rect -80355 -25310 -80347 -25266
rect -80255 -25310 -80247 -25266
rect -80155 -25310 -80147 -25266
rect -80055 -25310 -80047 -25266
rect -79955 -25310 -79947 -25266
rect -79855 -25310 -79847 -25266
rect -79755 -25310 -79747 -25266
rect -79655 -25310 -79647 -25266
rect -79555 -25310 -79547 -25266
rect -79455 -25310 -79447 -25266
rect -79355 -25310 -79347 -25266
rect -79255 -25310 -79247 -25266
rect -78755 -25310 -78747 -25266
rect -78655 -25310 -78647 -25266
rect -78555 -25310 -78547 -25266
rect -78455 -25310 -78447 -25266
rect -78355 -25310 -78347 -25266
rect -78255 -25310 -78247 -25266
rect -78155 -25310 -78147 -25266
rect -78055 -25310 -78047 -25266
rect -77955 -25310 -77947 -25266
rect -77855 -25310 -77847 -25266
rect -77755 -25310 -77747 -25266
rect -77655 -25310 -77647 -25266
rect -77555 -25310 -77547 -25266
rect -77455 -25310 -77447 -25266
rect -77355 -25310 -77347 -25266
rect -77255 -25310 -77247 -25266
rect -76755 -25310 -76747 -25266
rect -76655 -25310 -76647 -25266
rect -76555 -25310 -76547 -25266
rect -76455 -25310 -76447 -25266
rect -76355 -25310 -76347 -25266
rect -76255 -25310 -76247 -25266
rect -76155 -25310 -76147 -25266
rect -76055 -25310 -76047 -25266
rect -75955 -25310 -75947 -25266
rect -75855 -25310 -75847 -25266
rect -75755 -25310 -75747 -25266
rect -75655 -25310 -75647 -25266
rect -75555 -25310 -75547 -25266
rect -75455 -25310 -75447 -25266
rect -75355 -25310 -75347 -25266
rect -75255 -25310 -75247 -25266
rect -82799 -25366 -82755 -25358
rect -82699 -25366 -82655 -25358
rect -82599 -25366 -82555 -25358
rect -82499 -25366 -82455 -25358
rect -82399 -25366 -82355 -25358
rect -82299 -25366 -82255 -25358
rect -82199 -25366 -82155 -25358
rect -82099 -25366 -82055 -25358
rect -81999 -25366 -81955 -25358
rect -81899 -25366 -81855 -25358
rect -81799 -25366 -81755 -25358
rect -81699 -25366 -81655 -25358
rect -81599 -25366 -81555 -25358
rect -81499 -25366 -81455 -25358
rect -81399 -25366 -81355 -25358
rect -81299 -25366 -81255 -25358
rect -80799 -25366 -80755 -25358
rect -80699 -25366 -80655 -25358
rect -80599 -25366 -80555 -25358
rect -80499 -25366 -80455 -25358
rect -80399 -25366 -80355 -25358
rect -80299 -25366 -80255 -25358
rect -80199 -25366 -80155 -25358
rect -80099 -25366 -80055 -25358
rect -79999 -25366 -79955 -25358
rect -79899 -25366 -79855 -25358
rect -79799 -25366 -79755 -25358
rect -79699 -25366 -79655 -25358
rect -79599 -25366 -79555 -25358
rect -79499 -25366 -79455 -25358
rect -79399 -25366 -79355 -25358
rect -79299 -25366 -79255 -25358
rect -78799 -25366 -78755 -25358
rect -78699 -25366 -78655 -25358
rect -78599 -25366 -78555 -25358
rect -78499 -25366 -78455 -25358
rect -78399 -25366 -78355 -25358
rect -78299 -25366 -78255 -25358
rect -78199 -25366 -78155 -25358
rect -78099 -25366 -78055 -25358
rect -77999 -25366 -77955 -25358
rect -77899 -25366 -77855 -25358
rect -77799 -25366 -77755 -25358
rect -77699 -25366 -77655 -25358
rect -77599 -25366 -77555 -25358
rect -77499 -25366 -77455 -25358
rect -77399 -25366 -77355 -25358
rect -77299 -25366 -77255 -25358
rect -76799 -25366 -76755 -25358
rect -76699 -25366 -76655 -25358
rect -76599 -25366 -76555 -25358
rect -76499 -25366 -76455 -25358
rect -76399 -25366 -76355 -25358
rect -76299 -25366 -76255 -25358
rect -76199 -25366 -76155 -25358
rect -76099 -25366 -76055 -25358
rect -75999 -25366 -75955 -25358
rect -75899 -25366 -75855 -25358
rect -75799 -25366 -75755 -25358
rect -75699 -25366 -75655 -25358
rect -75599 -25366 -75555 -25358
rect -75499 -25366 -75455 -25358
rect -75399 -25366 -75355 -25358
rect -75299 -25366 -75255 -25358
rect -82755 -25410 -82747 -25366
rect -82655 -25410 -82647 -25366
rect -82555 -25410 -82547 -25366
rect -82455 -25410 -82447 -25366
rect -82355 -25410 -82347 -25366
rect -82255 -25410 -82247 -25366
rect -82155 -25410 -82147 -25366
rect -82055 -25410 -82047 -25366
rect -81955 -25410 -81947 -25366
rect -81855 -25410 -81847 -25366
rect -81755 -25410 -81747 -25366
rect -81655 -25410 -81647 -25366
rect -81555 -25410 -81547 -25366
rect -81455 -25410 -81447 -25366
rect -81355 -25410 -81347 -25366
rect -81255 -25410 -81247 -25366
rect -80755 -25410 -80747 -25366
rect -80655 -25410 -80647 -25366
rect -80555 -25410 -80547 -25366
rect -80455 -25410 -80447 -25366
rect -80355 -25410 -80347 -25366
rect -80255 -25410 -80247 -25366
rect -80155 -25410 -80147 -25366
rect -80055 -25410 -80047 -25366
rect -79955 -25410 -79947 -25366
rect -79855 -25410 -79847 -25366
rect -79755 -25410 -79747 -25366
rect -79655 -25410 -79647 -25366
rect -79555 -25410 -79547 -25366
rect -79455 -25410 -79447 -25366
rect -79355 -25410 -79347 -25366
rect -79255 -25410 -79247 -25366
rect -78755 -25410 -78747 -25366
rect -78655 -25410 -78647 -25366
rect -78555 -25410 -78547 -25366
rect -78455 -25410 -78447 -25366
rect -78355 -25410 -78347 -25366
rect -78255 -25410 -78247 -25366
rect -78155 -25410 -78147 -25366
rect -78055 -25410 -78047 -25366
rect -77955 -25410 -77947 -25366
rect -77855 -25410 -77847 -25366
rect -77755 -25410 -77747 -25366
rect -77655 -25410 -77647 -25366
rect -77555 -25410 -77547 -25366
rect -77455 -25410 -77447 -25366
rect -77355 -25410 -77347 -25366
rect -77255 -25410 -77247 -25366
rect -76755 -25410 -76747 -25366
rect -76655 -25410 -76647 -25366
rect -76555 -25410 -76547 -25366
rect -76455 -25410 -76447 -25366
rect -76355 -25410 -76347 -25366
rect -76255 -25410 -76247 -25366
rect -76155 -25410 -76147 -25366
rect -76055 -25410 -76047 -25366
rect -75955 -25410 -75947 -25366
rect -75855 -25410 -75847 -25366
rect -75755 -25410 -75747 -25366
rect -75655 -25410 -75647 -25366
rect -75555 -25410 -75547 -25366
rect -75455 -25410 -75447 -25366
rect -75355 -25410 -75347 -25366
rect -75255 -25410 -75247 -25366
rect -82799 -25466 -82755 -25458
rect -82699 -25466 -82655 -25458
rect -82599 -25466 -82555 -25458
rect -82499 -25466 -82455 -25458
rect -82399 -25466 -82355 -25458
rect -82299 -25466 -82255 -25458
rect -82199 -25466 -82155 -25458
rect -82099 -25466 -82055 -25458
rect -81999 -25466 -81955 -25458
rect -81899 -25466 -81855 -25458
rect -81799 -25466 -81755 -25458
rect -81699 -25466 -81655 -25458
rect -81599 -25466 -81555 -25458
rect -81499 -25466 -81455 -25458
rect -81399 -25466 -81355 -25458
rect -81299 -25466 -81255 -25458
rect -80799 -25466 -80755 -25458
rect -80699 -25466 -80655 -25458
rect -80599 -25466 -80555 -25458
rect -80499 -25466 -80455 -25458
rect -80399 -25466 -80355 -25458
rect -80299 -25466 -80255 -25458
rect -80199 -25466 -80155 -25458
rect -80099 -25466 -80055 -25458
rect -79999 -25466 -79955 -25458
rect -79899 -25466 -79855 -25458
rect -79799 -25466 -79755 -25458
rect -79699 -25466 -79655 -25458
rect -79599 -25466 -79555 -25458
rect -79499 -25466 -79455 -25458
rect -79399 -25466 -79355 -25458
rect -79299 -25466 -79255 -25458
rect -78799 -25466 -78755 -25458
rect -78699 -25466 -78655 -25458
rect -78599 -25466 -78555 -25458
rect -78499 -25466 -78455 -25458
rect -78399 -25466 -78355 -25458
rect -78299 -25466 -78255 -25458
rect -78199 -25466 -78155 -25458
rect -78099 -25466 -78055 -25458
rect -77999 -25466 -77955 -25458
rect -77899 -25466 -77855 -25458
rect -77799 -25466 -77755 -25458
rect -77699 -25466 -77655 -25458
rect -77599 -25466 -77555 -25458
rect -77499 -25466 -77455 -25458
rect -77399 -25466 -77355 -25458
rect -77299 -25466 -77255 -25458
rect -76799 -25466 -76755 -25458
rect -76699 -25466 -76655 -25458
rect -76599 -25466 -76555 -25458
rect -76499 -25466 -76455 -25458
rect -76399 -25466 -76355 -25458
rect -76299 -25466 -76255 -25458
rect -76199 -25466 -76155 -25458
rect -76099 -25466 -76055 -25458
rect -75999 -25466 -75955 -25458
rect -75899 -25466 -75855 -25458
rect -75799 -25466 -75755 -25458
rect -75699 -25466 -75655 -25458
rect -75599 -25466 -75555 -25458
rect -75499 -25466 -75455 -25458
rect -75399 -25466 -75355 -25458
rect -75299 -25466 -75255 -25458
rect -82755 -25510 -82747 -25466
rect -82655 -25510 -82647 -25466
rect -82555 -25510 -82547 -25466
rect -82455 -25510 -82447 -25466
rect -82355 -25510 -82347 -25466
rect -82255 -25510 -82247 -25466
rect -82155 -25510 -82147 -25466
rect -82055 -25510 -82047 -25466
rect -81955 -25510 -81947 -25466
rect -81855 -25510 -81847 -25466
rect -81755 -25510 -81747 -25466
rect -81655 -25510 -81647 -25466
rect -81555 -25510 -81547 -25466
rect -81455 -25510 -81447 -25466
rect -81355 -25510 -81347 -25466
rect -81255 -25510 -81247 -25466
rect -80755 -25510 -80747 -25466
rect -80655 -25510 -80647 -25466
rect -80555 -25510 -80547 -25466
rect -80455 -25510 -80447 -25466
rect -80355 -25510 -80347 -25466
rect -80255 -25510 -80247 -25466
rect -80155 -25510 -80147 -25466
rect -80055 -25510 -80047 -25466
rect -79955 -25510 -79947 -25466
rect -79855 -25510 -79847 -25466
rect -79755 -25510 -79747 -25466
rect -79655 -25510 -79647 -25466
rect -79555 -25510 -79547 -25466
rect -79455 -25510 -79447 -25466
rect -79355 -25510 -79347 -25466
rect -79255 -25510 -79247 -25466
rect -78755 -25510 -78747 -25466
rect -78655 -25510 -78647 -25466
rect -78555 -25510 -78547 -25466
rect -78455 -25510 -78447 -25466
rect -78355 -25510 -78347 -25466
rect -78255 -25510 -78247 -25466
rect -78155 -25510 -78147 -25466
rect -78055 -25510 -78047 -25466
rect -77955 -25510 -77947 -25466
rect -77855 -25510 -77847 -25466
rect -77755 -25510 -77747 -25466
rect -77655 -25510 -77647 -25466
rect -77555 -25510 -77547 -25466
rect -77455 -25510 -77447 -25466
rect -77355 -25510 -77347 -25466
rect -77255 -25510 -77247 -25466
rect -76755 -25510 -76747 -25466
rect -76655 -25510 -76647 -25466
rect -76555 -25510 -76547 -25466
rect -76455 -25510 -76447 -25466
rect -76355 -25510 -76347 -25466
rect -76255 -25510 -76247 -25466
rect -76155 -25510 -76147 -25466
rect -76055 -25510 -76047 -25466
rect -75955 -25510 -75947 -25466
rect -75855 -25510 -75847 -25466
rect -75755 -25510 -75747 -25466
rect -75655 -25510 -75647 -25466
rect -75555 -25510 -75547 -25466
rect -75455 -25510 -75447 -25466
rect -75355 -25510 -75347 -25466
rect -75255 -25510 -75247 -25466
rect -82799 -25566 -82755 -25558
rect -82699 -25566 -82655 -25558
rect -82599 -25566 -82555 -25558
rect -82499 -25566 -82455 -25558
rect -82399 -25566 -82355 -25558
rect -82299 -25566 -82255 -25558
rect -82199 -25566 -82155 -25558
rect -82099 -25566 -82055 -25558
rect -81999 -25566 -81955 -25558
rect -81899 -25566 -81855 -25558
rect -81799 -25566 -81755 -25558
rect -81699 -25566 -81655 -25558
rect -81599 -25566 -81555 -25558
rect -81499 -25566 -81455 -25558
rect -81399 -25566 -81355 -25558
rect -81299 -25566 -81255 -25558
rect -80799 -25566 -80755 -25558
rect -80699 -25566 -80655 -25558
rect -80599 -25566 -80555 -25558
rect -80499 -25566 -80455 -25558
rect -80399 -25566 -80355 -25558
rect -80299 -25566 -80255 -25558
rect -80199 -25566 -80155 -25558
rect -80099 -25566 -80055 -25558
rect -79999 -25566 -79955 -25558
rect -79899 -25566 -79855 -25558
rect -79799 -25566 -79755 -25558
rect -79699 -25566 -79655 -25558
rect -79599 -25566 -79555 -25558
rect -79499 -25566 -79455 -25558
rect -79399 -25566 -79355 -25558
rect -79299 -25566 -79255 -25558
rect -78799 -25566 -78755 -25558
rect -78699 -25566 -78655 -25558
rect -78599 -25566 -78555 -25558
rect -78499 -25566 -78455 -25558
rect -78399 -25566 -78355 -25558
rect -78299 -25566 -78255 -25558
rect -78199 -25566 -78155 -25558
rect -78099 -25566 -78055 -25558
rect -77999 -25566 -77955 -25558
rect -77899 -25566 -77855 -25558
rect -77799 -25566 -77755 -25558
rect -77699 -25566 -77655 -25558
rect -77599 -25566 -77555 -25558
rect -77499 -25566 -77455 -25558
rect -77399 -25566 -77355 -25558
rect -77299 -25566 -77255 -25558
rect -76799 -25566 -76755 -25558
rect -76699 -25566 -76655 -25558
rect -76599 -25566 -76555 -25558
rect -76499 -25566 -76455 -25558
rect -76399 -25566 -76355 -25558
rect -76299 -25566 -76255 -25558
rect -76199 -25566 -76155 -25558
rect -76099 -25566 -76055 -25558
rect -75999 -25566 -75955 -25558
rect -75899 -25566 -75855 -25558
rect -75799 -25566 -75755 -25558
rect -75699 -25566 -75655 -25558
rect -75599 -25566 -75555 -25558
rect -75499 -25566 -75455 -25558
rect -75399 -25566 -75355 -25558
rect -75299 -25566 -75255 -25558
rect -82755 -25610 -82747 -25566
rect -82655 -25610 -82647 -25566
rect -82555 -25610 -82547 -25566
rect -82455 -25610 -82447 -25566
rect -82355 -25610 -82347 -25566
rect -82255 -25610 -82247 -25566
rect -82155 -25610 -82147 -25566
rect -82055 -25610 -82047 -25566
rect -81955 -25610 -81947 -25566
rect -81855 -25610 -81847 -25566
rect -81755 -25610 -81747 -25566
rect -81655 -25610 -81647 -25566
rect -81555 -25610 -81547 -25566
rect -81455 -25610 -81447 -25566
rect -81355 -25610 -81347 -25566
rect -81255 -25610 -81247 -25566
rect -80755 -25610 -80747 -25566
rect -80655 -25610 -80647 -25566
rect -80555 -25610 -80547 -25566
rect -80455 -25610 -80447 -25566
rect -80355 -25610 -80347 -25566
rect -80255 -25610 -80247 -25566
rect -80155 -25610 -80147 -25566
rect -80055 -25610 -80047 -25566
rect -79955 -25610 -79947 -25566
rect -79855 -25610 -79847 -25566
rect -79755 -25610 -79747 -25566
rect -79655 -25610 -79647 -25566
rect -79555 -25610 -79547 -25566
rect -79455 -25610 -79447 -25566
rect -79355 -25610 -79347 -25566
rect -79255 -25610 -79247 -25566
rect -78755 -25610 -78747 -25566
rect -78655 -25610 -78647 -25566
rect -78555 -25610 -78547 -25566
rect -78455 -25610 -78447 -25566
rect -78355 -25610 -78347 -25566
rect -78255 -25610 -78247 -25566
rect -78155 -25610 -78147 -25566
rect -78055 -25610 -78047 -25566
rect -77955 -25610 -77947 -25566
rect -77855 -25610 -77847 -25566
rect -77755 -25610 -77747 -25566
rect -77655 -25610 -77647 -25566
rect -77555 -25610 -77547 -25566
rect -77455 -25610 -77447 -25566
rect -77355 -25610 -77347 -25566
rect -77255 -25610 -77247 -25566
rect -76755 -25610 -76747 -25566
rect -76655 -25610 -76647 -25566
rect -76555 -25610 -76547 -25566
rect -76455 -25610 -76447 -25566
rect -76355 -25610 -76347 -25566
rect -76255 -25610 -76247 -25566
rect -76155 -25610 -76147 -25566
rect -76055 -25610 -76047 -25566
rect -75955 -25610 -75947 -25566
rect -75855 -25610 -75847 -25566
rect -75755 -25610 -75747 -25566
rect -75655 -25610 -75647 -25566
rect -75555 -25610 -75547 -25566
rect -75455 -25610 -75447 -25566
rect -75355 -25610 -75347 -25566
rect -75255 -25610 -75247 -25566
rect -82799 -25666 -82755 -25658
rect -82699 -25666 -82655 -25658
rect -82599 -25666 -82555 -25658
rect -82499 -25666 -82455 -25658
rect -82399 -25666 -82355 -25658
rect -82299 -25666 -82255 -25658
rect -82199 -25666 -82155 -25658
rect -82099 -25666 -82055 -25658
rect -81999 -25666 -81955 -25658
rect -81899 -25666 -81855 -25658
rect -81799 -25666 -81755 -25658
rect -81699 -25666 -81655 -25658
rect -81599 -25666 -81555 -25658
rect -81499 -25666 -81455 -25658
rect -81399 -25666 -81355 -25658
rect -81299 -25666 -81255 -25658
rect -80799 -25666 -80755 -25658
rect -80699 -25666 -80655 -25658
rect -80599 -25666 -80555 -25658
rect -80499 -25666 -80455 -25658
rect -80399 -25666 -80355 -25658
rect -80299 -25666 -80255 -25658
rect -80199 -25666 -80155 -25658
rect -80099 -25666 -80055 -25658
rect -79999 -25666 -79955 -25658
rect -79899 -25666 -79855 -25658
rect -79799 -25666 -79755 -25658
rect -79699 -25666 -79655 -25658
rect -79599 -25666 -79555 -25658
rect -79499 -25666 -79455 -25658
rect -79399 -25666 -79355 -25658
rect -79299 -25666 -79255 -25658
rect -78799 -25666 -78755 -25658
rect -78699 -25666 -78655 -25658
rect -78599 -25666 -78555 -25658
rect -78499 -25666 -78455 -25658
rect -78399 -25666 -78355 -25658
rect -78299 -25666 -78255 -25658
rect -78199 -25666 -78155 -25658
rect -78099 -25666 -78055 -25658
rect -77999 -25666 -77955 -25658
rect -77899 -25666 -77855 -25658
rect -77799 -25666 -77755 -25658
rect -77699 -25666 -77655 -25658
rect -77599 -25666 -77555 -25658
rect -77499 -25666 -77455 -25658
rect -77399 -25666 -77355 -25658
rect -77299 -25666 -77255 -25658
rect -76799 -25666 -76755 -25658
rect -76699 -25666 -76655 -25658
rect -76599 -25666 -76555 -25658
rect -76499 -25666 -76455 -25658
rect -76399 -25666 -76355 -25658
rect -76299 -25666 -76255 -25658
rect -76199 -25666 -76155 -25658
rect -76099 -25666 -76055 -25658
rect -75999 -25666 -75955 -25658
rect -75899 -25666 -75855 -25658
rect -75799 -25666 -75755 -25658
rect -75699 -25666 -75655 -25658
rect -75599 -25666 -75555 -25658
rect -75499 -25666 -75455 -25658
rect -75399 -25666 -75355 -25658
rect -75299 -25666 -75255 -25658
rect -82755 -25710 -82747 -25666
rect -82655 -25710 -82647 -25666
rect -82555 -25710 -82547 -25666
rect -82455 -25710 -82447 -25666
rect -82355 -25710 -82347 -25666
rect -82255 -25710 -82247 -25666
rect -82155 -25710 -82147 -25666
rect -82055 -25710 -82047 -25666
rect -81955 -25710 -81947 -25666
rect -81855 -25710 -81847 -25666
rect -81755 -25710 -81747 -25666
rect -81655 -25710 -81647 -25666
rect -81555 -25710 -81547 -25666
rect -81455 -25710 -81447 -25666
rect -81355 -25710 -81347 -25666
rect -81255 -25710 -81247 -25666
rect -80755 -25710 -80747 -25666
rect -80655 -25710 -80647 -25666
rect -80555 -25710 -80547 -25666
rect -80455 -25710 -80447 -25666
rect -80355 -25710 -80347 -25666
rect -80255 -25710 -80247 -25666
rect -80155 -25710 -80147 -25666
rect -80055 -25710 -80047 -25666
rect -79955 -25710 -79947 -25666
rect -79855 -25710 -79847 -25666
rect -79755 -25710 -79747 -25666
rect -79655 -25710 -79647 -25666
rect -79555 -25710 -79547 -25666
rect -79455 -25710 -79447 -25666
rect -79355 -25710 -79347 -25666
rect -79255 -25710 -79247 -25666
rect -78755 -25710 -78747 -25666
rect -78655 -25710 -78647 -25666
rect -78555 -25710 -78547 -25666
rect -78455 -25710 -78447 -25666
rect -78355 -25710 -78347 -25666
rect -78255 -25710 -78247 -25666
rect -78155 -25710 -78147 -25666
rect -78055 -25710 -78047 -25666
rect -77955 -25710 -77947 -25666
rect -77855 -25710 -77847 -25666
rect -77755 -25710 -77747 -25666
rect -77655 -25710 -77647 -25666
rect -77555 -25710 -77547 -25666
rect -77455 -25710 -77447 -25666
rect -77355 -25710 -77347 -25666
rect -77255 -25710 -77247 -25666
rect -76755 -25710 -76747 -25666
rect -76655 -25710 -76647 -25666
rect -76555 -25710 -76547 -25666
rect -76455 -25710 -76447 -25666
rect -76355 -25710 -76347 -25666
rect -76255 -25710 -76247 -25666
rect -76155 -25710 -76147 -25666
rect -76055 -25710 -76047 -25666
rect -75955 -25710 -75947 -25666
rect -75855 -25710 -75847 -25666
rect -75755 -25710 -75747 -25666
rect -75655 -25710 -75647 -25666
rect -75555 -25710 -75547 -25666
rect -75455 -25710 -75447 -25666
rect -75355 -25710 -75347 -25666
rect -75255 -25710 -75247 -25666
rect -82799 -25766 -82755 -25758
rect -82699 -25766 -82655 -25758
rect -82599 -25766 -82555 -25758
rect -82499 -25766 -82455 -25758
rect -82399 -25766 -82355 -25758
rect -82299 -25766 -82255 -25758
rect -82199 -25766 -82155 -25758
rect -82099 -25766 -82055 -25758
rect -81999 -25766 -81955 -25758
rect -81899 -25766 -81855 -25758
rect -81799 -25766 -81755 -25758
rect -81699 -25766 -81655 -25758
rect -81599 -25766 -81555 -25758
rect -81499 -25766 -81455 -25758
rect -81399 -25766 -81355 -25758
rect -81299 -25766 -81255 -25758
rect -80799 -25766 -80755 -25758
rect -80699 -25766 -80655 -25758
rect -80599 -25766 -80555 -25758
rect -80499 -25766 -80455 -25758
rect -80399 -25766 -80355 -25758
rect -80299 -25766 -80255 -25758
rect -80199 -25766 -80155 -25758
rect -80099 -25766 -80055 -25758
rect -79999 -25766 -79955 -25758
rect -79899 -25766 -79855 -25758
rect -79799 -25766 -79755 -25758
rect -79699 -25766 -79655 -25758
rect -79599 -25766 -79555 -25758
rect -79499 -25766 -79455 -25758
rect -79399 -25766 -79355 -25758
rect -79299 -25766 -79255 -25758
rect -78799 -25766 -78755 -25758
rect -78699 -25766 -78655 -25758
rect -78599 -25766 -78555 -25758
rect -78499 -25766 -78455 -25758
rect -78399 -25766 -78355 -25758
rect -78299 -25766 -78255 -25758
rect -78199 -25766 -78155 -25758
rect -78099 -25766 -78055 -25758
rect -77999 -25766 -77955 -25758
rect -77899 -25766 -77855 -25758
rect -77799 -25766 -77755 -25758
rect -77699 -25766 -77655 -25758
rect -77599 -25766 -77555 -25758
rect -77499 -25766 -77455 -25758
rect -77399 -25766 -77355 -25758
rect -77299 -25766 -77255 -25758
rect -76799 -25766 -76755 -25758
rect -76699 -25766 -76655 -25758
rect -76599 -25766 -76555 -25758
rect -76499 -25766 -76455 -25758
rect -76399 -25766 -76355 -25758
rect -76299 -25766 -76255 -25758
rect -76199 -25766 -76155 -25758
rect -76099 -25766 -76055 -25758
rect -75999 -25766 -75955 -25758
rect -75899 -25766 -75855 -25758
rect -75799 -25766 -75755 -25758
rect -75699 -25766 -75655 -25758
rect -75599 -25766 -75555 -25758
rect -75499 -25766 -75455 -25758
rect -75399 -25766 -75355 -25758
rect -75299 -25766 -75255 -25758
rect -82755 -25810 -82747 -25766
rect -82655 -25810 -82647 -25766
rect -82555 -25810 -82547 -25766
rect -82455 -25810 -82447 -25766
rect -82355 -25810 -82347 -25766
rect -82255 -25810 -82247 -25766
rect -82155 -25810 -82147 -25766
rect -82055 -25810 -82047 -25766
rect -81955 -25810 -81947 -25766
rect -81855 -25810 -81847 -25766
rect -81755 -25810 -81747 -25766
rect -81655 -25810 -81647 -25766
rect -81555 -25810 -81547 -25766
rect -81455 -25810 -81447 -25766
rect -81355 -25810 -81347 -25766
rect -81255 -25810 -81247 -25766
rect -80755 -25810 -80747 -25766
rect -80655 -25810 -80647 -25766
rect -80555 -25810 -80547 -25766
rect -80455 -25810 -80447 -25766
rect -80355 -25810 -80347 -25766
rect -80255 -25810 -80247 -25766
rect -80155 -25810 -80147 -25766
rect -80055 -25810 -80047 -25766
rect -79955 -25810 -79947 -25766
rect -79855 -25810 -79847 -25766
rect -79755 -25810 -79747 -25766
rect -79655 -25810 -79647 -25766
rect -79555 -25810 -79547 -25766
rect -79455 -25810 -79447 -25766
rect -79355 -25810 -79347 -25766
rect -79255 -25810 -79247 -25766
rect -78755 -25810 -78747 -25766
rect -78655 -25810 -78647 -25766
rect -78555 -25810 -78547 -25766
rect -78455 -25810 -78447 -25766
rect -78355 -25810 -78347 -25766
rect -78255 -25810 -78247 -25766
rect -78155 -25810 -78147 -25766
rect -78055 -25810 -78047 -25766
rect -77955 -25810 -77947 -25766
rect -77855 -25810 -77847 -25766
rect -77755 -25810 -77747 -25766
rect -77655 -25810 -77647 -25766
rect -77555 -25810 -77547 -25766
rect -77455 -25810 -77447 -25766
rect -77355 -25810 -77347 -25766
rect -77255 -25810 -77247 -25766
rect -76755 -25810 -76747 -25766
rect -76655 -25810 -76647 -25766
rect -76555 -25810 -76547 -25766
rect -76455 -25810 -76447 -25766
rect -76355 -25810 -76347 -25766
rect -76255 -25810 -76247 -25766
rect -76155 -25810 -76147 -25766
rect -76055 -25810 -76047 -25766
rect -75955 -25810 -75947 -25766
rect -75855 -25810 -75847 -25766
rect -75755 -25810 -75747 -25766
rect -75655 -25810 -75647 -25766
rect -75555 -25810 -75547 -25766
rect -75455 -25810 -75447 -25766
rect -75355 -25810 -75347 -25766
rect -75255 -25810 -75247 -25766
rect -82799 -25866 -82755 -25858
rect -82699 -25866 -82655 -25858
rect -82599 -25866 -82555 -25858
rect -82499 -25866 -82455 -25858
rect -82399 -25866 -82355 -25858
rect -82299 -25866 -82255 -25858
rect -82199 -25866 -82155 -25858
rect -82099 -25866 -82055 -25858
rect -81999 -25866 -81955 -25858
rect -81899 -25866 -81855 -25858
rect -81799 -25866 -81755 -25858
rect -81699 -25866 -81655 -25858
rect -81599 -25866 -81555 -25858
rect -81499 -25866 -81455 -25858
rect -81399 -25866 -81355 -25858
rect -81299 -25866 -81255 -25858
rect -80799 -25866 -80755 -25858
rect -80699 -25866 -80655 -25858
rect -80599 -25866 -80555 -25858
rect -80499 -25866 -80455 -25858
rect -80399 -25866 -80355 -25858
rect -80299 -25866 -80255 -25858
rect -80199 -25866 -80155 -25858
rect -80099 -25866 -80055 -25858
rect -79999 -25866 -79955 -25858
rect -79899 -25866 -79855 -25858
rect -79799 -25866 -79755 -25858
rect -79699 -25866 -79655 -25858
rect -79599 -25866 -79555 -25858
rect -79499 -25866 -79455 -25858
rect -79399 -25866 -79355 -25858
rect -79299 -25866 -79255 -25858
rect -78799 -25866 -78755 -25858
rect -78699 -25866 -78655 -25858
rect -78599 -25866 -78555 -25858
rect -78499 -25866 -78455 -25858
rect -78399 -25866 -78355 -25858
rect -78299 -25866 -78255 -25858
rect -78199 -25866 -78155 -25858
rect -78099 -25866 -78055 -25858
rect -77999 -25866 -77955 -25858
rect -77899 -25866 -77855 -25858
rect -77799 -25866 -77755 -25858
rect -77699 -25866 -77655 -25858
rect -77599 -25866 -77555 -25858
rect -77499 -25866 -77455 -25858
rect -77399 -25866 -77355 -25858
rect -77299 -25866 -77255 -25858
rect -76799 -25866 -76755 -25858
rect -76699 -25866 -76655 -25858
rect -76599 -25866 -76555 -25858
rect -76499 -25866 -76455 -25858
rect -76399 -25866 -76355 -25858
rect -76299 -25866 -76255 -25858
rect -76199 -25866 -76155 -25858
rect -76099 -25866 -76055 -25858
rect -75999 -25866 -75955 -25858
rect -75899 -25866 -75855 -25858
rect -75799 -25866 -75755 -25858
rect -75699 -25866 -75655 -25858
rect -75599 -25866 -75555 -25858
rect -75499 -25866 -75455 -25858
rect -75399 -25866 -75355 -25858
rect -75299 -25866 -75255 -25858
rect -82755 -25910 -82747 -25866
rect -82655 -25910 -82647 -25866
rect -82555 -25910 -82547 -25866
rect -82455 -25910 -82447 -25866
rect -82355 -25910 -82347 -25866
rect -82255 -25910 -82247 -25866
rect -82155 -25910 -82147 -25866
rect -82055 -25910 -82047 -25866
rect -81955 -25910 -81947 -25866
rect -81855 -25910 -81847 -25866
rect -81755 -25910 -81747 -25866
rect -81655 -25910 -81647 -25866
rect -81555 -25910 -81547 -25866
rect -81455 -25910 -81447 -25866
rect -81355 -25910 -81347 -25866
rect -81255 -25910 -81247 -25866
rect -80755 -25910 -80747 -25866
rect -80655 -25910 -80647 -25866
rect -80555 -25910 -80547 -25866
rect -80455 -25910 -80447 -25866
rect -80355 -25910 -80347 -25866
rect -80255 -25910 -80247 -25866
rect -80155 -25910 -80147 -25866
rect -80055 -25910 -80047 -25866
rect -79955 -25910 -79947 -25866
rect -79855 -25910 -79847 -25866
rect -79755 -25910 -79747 -25866
rect -79655 -25910 -79647 -25866
rect -79555 -25910 -79547 -25866
rect -79455 -25910 -79447 -25866
rect -79355 -25910 -79347 -25866
rect -79255 -25910 -79247 -25866
rect -78755 -25910 -78747 -25866
rect -78655 -25910 -78647 -25866
rect -78555 -25910 -78547 -25866
rect -78455 -25910 -78447 -25866
rect -78355 -25910 -78347 -25866
rect -78255 -25910 -78247 -25866
rect -78155 -25910 -78147 -25866
rect -78055 -25910 -78047 -25866
rect -77955 -25910 -77947 -25866
rect -77855 -25910 -77847 -25866
rect -77755 -25910 -77747 -25866
rect -77655 -25910 -77647 -25866
rect -77555 -25910 -77547 -25866
rect -77455 -25910 -77447 -25866
rect -77355 -25910 -77347 -25866
rect -77255 -25910 -77247 -25866
rect -76755 -25910 -76747 -25866
rect -76655 -25910 -76647 -25866
rect -76555 -25910 -76547 -25866
rect -76455 -25910 -76447 -25866
rect -76355 -25910 -76347 -25866
rect -76255 -25910 -76247 -25866
rect -76155 -25910 -76147 -25866
rect -76055 -25910 -76047 -25866
rect -75955 -25910 -75947 -25866
rect -75855 -25910 -75847 -25866
rect -75755 -25910 -75747 -25866
rect -75655 -25910 -75647 -25866
rect -75555 -25910 -75547 -25866
rect -75455 -25910 -75447 -25866
rect -75355 -25910 -75347 -25866
rect -75255 -25910 -75247 -25866
rect 145268 -165615 145312 -165607
rect 145368 -165615 145412 -165607
rect 145468 -165615 145512 -165607
rect 145568 -165615 145612 -165607
rect 145668 -165615 145712 -165607
rect 145768 -165615 145812 -165607
rect 145868 -165615 145912 -165607
rect 145968 -165615 146012 -165607
rect 146068 -165615 146112 -165607
rect 146168 -165615 146212 -165607
rect 146268 -165615 146312 -165607
rect 146368 -165615 146412 -165607
rect 146468 -165615 146512 -165607
rect 146568 -165615 146612 -165607
rect 146668 -165615 146712 -165607
rect 146768 -165615 146812 -165607
rect 147268 -165615 147312 -165607
rect 147368 -165615 147412 -165607
rect 147468 -165615 147512 -165607
rect 147568 -165615 147612 -165607
rect 147668 -165615 147712 -165607
rect 147768 -165615 147812 -165607
rect 147868 -165615 147912 -165607
rect 147968 -165615 148012 -165607
rect 148068 -165615 148112 -165607
rect 148168 -165615 148212 -165607
rect 148268 -165615 148312 -165607
rect 148368 -165615 148412 -165607
rect 148468 -165615 148512 -165607
rect 148568 -165615 148612 -165607
rect 148668 -165615 148712 -165607
rect 148768 -165615 148812 -165607
rect 149268 -165615 149312 -165607
rect 149368 -165615 149412 -165607
rect 149468 -165615 149512 -165607
rect 149568 -165615 149612 -165607
rect 149668 -165615 149712 -165607
rect 149768 -165615 149812 -165607
rect 149868 -165615 149912 -165607
rect 149968 -165615 150012 -165607
rect 150068 -165615 150112 -165607
rect 150168 -165615 150212 -165607
rect 150268 -165615 150312 -165607
rect 150368 -165615 150412 -165607
rect 150468 -165615 150512 -165607
rect 150568 -165615 150612 -165607
rect 150668 -165615 150712 -165607
rect 150768 -165615 150812 -165607
rect 151268 -165615 151312 -165607
rect 151368 -165615 151412 -165607
rect 151468 -165615 151512 -165607
rect 151568 -165615 151612 -165607
rect 151668 -165615 151712 -165607
rect 151768 -165615 151812 -165607
rect 151868 -165615 151912 -165607
rect 151968 -165615 152012 -165607
rect 152068 -165615 152112 -165607
rect 152168 -165615 152212 -165607
rect 152268 -165615 152312 -165607
rect 152368 -165615 152412 -165607
rect 152468 -165615 152512 -165607
rect 152568 -165615 152612 -165607
rect 152668 -165615 152712 -165607
rect 152768 -165615 152812 -165607
rect 145312 -165659 145320 -165615
rect 145412 -165659 145420 -165615
rect 145512 -165659 145520 -165615
rect 145612 -165659 145620 -165615
rect 145712 -165659 145720 -165615
rect 145812 -165659 145820 -165615
rect 145912 -165659 145920 -165615
rect 146012 -165659 146020 -165615
rect 146112 -165659 146120 -165615
rect 146212 -165659 146220 -165615
rect 146312 -165659 146320 -165615
rect 146412 -165659 146420 -165615
rect 146512 -165659 146520 -165615
rect 146612 -165659 146620 -165615
rect 146712 -165659 146720 -165615
rect 146812 -165659 146820 -165615
rect 147312 -165659 147320 -165615
rect 147412 -165659 147420 -165615
rect 147512 -165659 147520 -165615
rect 147612 -165659 147620 -165615
rect 147712 -165659 147720 -165615
rect 147812 -165659 147820 -165615
rect 147912 -165659 147920 -165615
rect 148012 -165659 148020 -165615
rect 148112 -165659 148120 -165615
rect 148212 -165659 148220 -165615
rect 148312 -165659 148320 -165615
rect 148412 -165659 148420 -165615
rect 148512 -165659 148520 -165615
rect 148612 -165659 148620 -165615
rect 148712 -165659 148720 -165615
rect 148812 -165659 148820 -165615
rect 149312 -165659 149320 -165615
rect 149412 -165659 149420 -165615
rect 149512 -165659 149520 -165615
rect 149612 -165659 149620 -165615
rect 149712 -165659 149720 -165615
rect 149812 -165659 149820 -165615
rect 149912 -165659 149920 -165615
rect 150012 -165659 150020 -165615
rect 150112 -165659 150120 -165615
rect 150212 -165659 150220 -165615
rect 150312 -165659 150320 -165615
rect 150412 -165659 150420 -165615
rect 150512 -165659 150520 -165615
rect 150612 -165659 150620 -165615
rect 150712 -165659 150720 -165615
rect 150812 -165659 150820 -165615
rect 151312 -165659 151320 -165615
rect 151412 -165659 151420 -165615
rect 151512 -165659 151520 -165615
rect 151612 -165659 151620 -165615
rect 151712 -165659 151720 -165615
rect 151812 -165659 151820 -165615
rect 151912 -165659 151920 -165615
rect 152012 -165659 152020 -165615
rect 152112 -165659 152120 -165615
rect 152212 -165659 152220 -165615
rect 152312 -165659 152320 -165615
rect 152412 -165659 152420 -165615
rect 152512 -165659 152520 -165615
rect 152612 -165659 152620 -165615
rect 152712 -165659 152720 -165615
rect 152812 -165659 152820 -165615
rect 145268 -165715 145312 -165707
rect 145368 -165715 145412 -165707
rect 145468 -165715 145512 -165707
rect 145568 -165715 145612 -165707
rect 145668 -165715 145712 -165707
rect 145768 -165715 145812 -165707
rect 145868 -165715 145912 -165707
rect 145968 -165715 146012 -165707
rect 146068 -165715 146112 -165707
rect 146168 -165715 146212 -165707
rect 146268 -165715 146312 -165707
rect 146368 -165715 146412 -165707
rect 146468 -165715 146512 -165707
rect 146568 -165715 146612 -165707
rect 146668 -165715 146712 -165707
rect 146768 -165715 146812 -165707
rect 147268 -165715 147312 -165707
rect 147368 -165715 147412 -165707
rect 147468 -165715 147512 -165707
rect 147568 -165715 147612 -165707
rect 147668 -165715 147712 -165707
rect 147768 -165715 147812 -165707
rect 147868 -165715 147912 -165707
rect 147968 -165715 148012 -165707
rect 148068 -165715 148112 -165707
rect 148168 -165715 148212 -165707
rect 148268 -165715 148312 -165707
rect 148368 -165715 148412 -165707
rect 148468 -165715 148512 -165707
rect 148568 -165715 148612 -165707
rect 148668 -165715 148712 -165707
rect 148768 -165715 148812 -165707
rect 149268 -165715 149312 -165707
rect 149368 -165715 149412 -165707
rect 149468 -165715 149512 -165707
rect 149568 -165715 149612 -165707
rect 149668 -165715 149712 -165707
rect 149768 -165715 149812 -165707
rect 149868 -165715 149912 -165707
rect 149968 -165715 150012 -165707
rect 150068 -165715 150112 -165707
rect 150168 -165715 150212 -165707
rect 150268 -165715 150312 -165707
rect 150368 -165715 150412 -165707
rect 150468 -165715 150512 -165707
rect 150568 -165715 150612 -165707
rect 150668 -165715 150712 -165707
rect 150768 -165715 150812 -165707
rect 151268 -165715 151312 -165707
rect 151368 -165715 151412 -165707
rect 151468 -165715 151512 -165707
rect 151568 -165715 151612 -165707
rect 151668 -165715 151712 -165707
rect 151768 -165715 151812 -165707
rect 151868 -165715 151912 -165707
rect 151968 -165715 152012 -165707
rect 152068 -165715 152112 -165707
rect 152168 -165715 152212 -165707
rect 152268 -165715 152312 -165707
rect 152368 -165715 152412 -165707
rect 152468 -165715 152512 -165707
rect 152568 -165715 152612 -165707
rect 152668 -165715 152712 -165707
rect 152768 -165715 152812 -165707
rect 145312 -165759 145320 -165715
rect 145412 -165759 145420 -165715
rect 145512 -165759 145520 -165715
rect 145612 -165759 145620 -165715
rect 145712 -165759 145720 -165715
rect 145812 -165759 145820 -165715
rect 145912 -165759 145920 -165715
rect 146012 -165759 146020 -165715
rect 146112 -165759 146120 -165715
rect 146212 -165759 146220 -165715
rect 146312 -165759 146320 -165715
rect 146412 -165759 146420 -165715
rect 146512 -165759 146520 -165715
rect 146612 -165759 146620 -165715
rect 146712 -165759 146720 -165715
rect 146812 -165759 146820 -165715
rect 147312 -165759 147320 -165715
rect 147412 -165759 147420 -165715
rect 147512 -165759 147520 -165715
rect 147612 -165759 147620 -165715
rect 147712 -165759 147720 -165715
rect 147812 -165759 147820 -165715
rect 147912 -165759 147920 -165715
rect 148012 -165759 148020 -165715
rect 148112 -165759 148120 -165715
rect 148212 -165759 148220 -165715
rect 148312 -165759 148320 -165715
rect 148412 -165759 148420 -165715
rect 148512 -165759 148520 -165715
rect 148612 -165759 148620 -165715
rect 148712 -165759 148720 -165715
rect 148812 -165759 148820 -165715
rect 149312 -165759 149320 -165715
rect 149412 -165759 149420 -165715
rect 149512 -165759 149520 -165715
rect 149612 -165759 149620 -165715
rect 149712 -165759 149720 -165715
rect 149812 -165759 149820 -165715
rect 149912 -165759 149920 -165715
rect 150012 -165759 150020 -165715
rect 150112 -165759 150120 -165715
rect 150212 -165759 150220 -165715
rect 150312 -165759 150320 -165715
rect 150412 -165759 150420 -165715
rect 150512 -165759 150520 -165715
rect 150612 -165759 150620 -165715
rect 150712 -165759 150720 -165715
rect 150812 -165759 150820 -165715
rect 151312 -165759 151320 -165715
rect 151412 -165759 151420 -165715
rect 151512 -165759 151520 -165715
rect 151612 -165759 151620 -165715
rect 151712 -165759 151720 -165715
rect 151812 -165759 151820 -165715
rect 151912 -165759 151920 -165715
rect 152012 -165759 152020 -165715
rect 152112 -165759 152120 -165715
rect 152212 -165759 152220 -165715
rect 152312 -165759 152320 -165715
rect 152412 -165759 152420 -165715
rect 152512 -165759 152520 -165715
rect 152612 -165759 152620 -165715
rect 152712 -165759 152720 -165715
rect 152812 -165759 152820 -165715
rect 145268 -165815 145312 -165807
rect 145368 -165815 145412 -165807
rect 145468 -165815 145512 -165807
rect 145568 -165815 145612 -165807
rect 145668 -165815 145712 -165807
rect 145768 -165815 145812 -165807
rect 145868 -165815 145912 -165807
rect 145968 -165815 146012 -165807
rect 146068 -165815 146112 -165807
rect 146168 -165815 146212 -165807
rect 146268 -165815 146312 -165807
rect 146368 -165815 146412 -165807
rect 146468 -165815 146512 -165807
rect 146568 -165815 146612 -165807
rect 146668 -165815 146712 -165807
rect 146768 -165815 146812 -165807
rect 147268 -165815 147312 -165807
rect 147368 -165815 147412 -165807
rect 147468 -165815 147512 -165807
rect 147568 -165815 147612 -165807
rect 147668 -165815 147712 -165807
rect 147768 -165815 147812 -165807
rect 147868 -165815 147912 -165807
rect 147968 -165815 148012 -165807
rect 148068 -165815 148112 -165807
rect 148168 -165815 148212 -165807
rect 148268 -165815 148312 -165807
rect 148368 -165815 148412 -165807
rect 148468 -165815 148512 -165807
rect 148568 -165815 148612 -165807
rect 148668 -165815 148712 -165807
rect 148768 -165815 148812 -165807
rect 149268 -165815 149312 -165807
rect 149368 -165815 149412 -165807
rect 149468 -165815 149512 -165807
rect 149568 -165815 149612 -165807
rect 149668 -165815 149712 -165807
rect 149768 -165815 149812 -165807
rect 149868 -165815 149912 -165807
rect 149968 -165815 150012 -165807
rect 150068 -165815 150112 -165807
rect 150168 -165815 150212 -165807
rect 150268 -165815 150312 -165807
rect 150368 -165815 150412 -165807
rect 150468 -165815 150512 -165807
rect 150568 -165815 150612 -165807
rect 150668 -165815 150712 -165807
rect 150768 -165815 150812 -165807
rect 151268 -165815 151312 -165807
rect 151368 -165815 151412 -165807
rect 151468 -165815 151512 -165807
rect 151568 -165815 151612 -165807
rect 151668 -165815 151712 -165807
rect 151768 -165815 151812 -165807
rect 151868 -165815 151912 -165807
rect 151968 -165815 152012 -165807
rect 152068 -165815 152112 -165807
rect 152168 -165815 152212 -165807
rect 152268 -165815 152312 -165807
rect 152368 -165815 152412 -165807
rect 152468 -165815 152512 -165807
rect 152568 -165815 152612 -165807
rect 152668 -165815 152712 -165807
rect 152768 -165815 152812 -165807
rect 145312 -165859 145320 -165815
rect 145412 -165859 145420 -165815
rect 145512 -165859 145520 -165815
rect 145612 -165859 145620 -165815
rect 145712 -165859 145720 -165815
rect 145812 -165859 145820 -165815
rect 145912 -165859 145920 -165815
rect 146012 -165859 146020 -165815
rect 146112 -165859 146120 -165815
rect 146212 -165859 146220 -165815
rect 146312 -165859 146320 -165815
rect 146412 -165859 146420 -165815
rect 146512 -165859 146520 -165815
rect 146612 -165859 146620 -165815
rect 146712 -165859 146720 -165815
rect 146812 -165859 146820 -165815
rect 147312 -165859 147320 -165815
rect 147412 -165859 147420 -165815
rect 147512 -165859 147520 -165815
rect 147612 -165859 147620 -165815
rect 147712 -165859 147720 -165815
rect 147812 -165859 147820 -165815
rect 147912 -165859 147920 -165815
rect 148012 -165859 148020 -165815
rect 148112 -165859 148120 -165815
rect 148212 -165859 148220 -165815
rect 148312 -165859 148320 -165815
rect 148412 -165859 148420 -165815
rect 148512 -165859 148520 -165815
rect 148612 -165859 148620 -165815
rect 148712 -165859 148720 -165815
rect 148812 -165859 148820 -165815
rect 149312 -165859 149320 -165815
rect 149412 -165859 149420 -165815
rect 149512 -165859 149520 -165815
rect 149612 -165859 149620 -165815
rect 149712 -165859 149720 -165815
rect 149812 -165859 149820 -165815
rect 149912 -165859 149920 -165815
rect 150012 -165859 150020 -165815
rect 150112 -165859 150120 -165815
rect 150212 -165859 150220 -165815
rect 150312 -165859 150320 -165815
rect 150412 -165859 150420 -165815
rect 150512 -165859 150520 -165815
rect 150612 -165859 150620 -165815
rect 150712 -165859 150720 -165815
rect 150812 -165859 150820 -165815
rect 151312 -165859 151320 -165815
rect 151412 -165859 151420 -165815
rect 151512 -165859 151520 -165815
rect 151612 -165859 151620 -165815
rect 151712 -165859 151720 -165815
rect 151812 -165859 151820 -165815
rect 151912 -165859 151920 -165815
rect 152012 -165859 152020 -165815
rect 152112 -165859 152120 -165815
rect 152212 -165859 152220 -165815
rect 152312 -165859 152320 -165815
rect 152412 -165859 152420 -165815
rect 152512 -165859 152520 -165815
rect 152612 -165859 152620 -165815
rect 152712 -165859 152720 -165815
rect 152812 -165859 152820 -165815
rect 145268 -165915 145312 -165907
rect 145368 -165915 145412 -165907
rect 145468 -165915 145512 -165907
rect 145568 -165915 145612 -165907
rect 145668 -165915 145712 -165907
rect 145768 -165915 145812 -165907
rect 145868 -165915 145912 -165907
rect 145968 -165915 146012 -165907
rect 146068 -165915 146112 -165907
rect 146168 -165915 146212 -165907
rect 146268 -165915 146312 -165907
rect 146368 -165915 146412 -165907
rect 146468 -165915 146512 -165907
rect 146568 -165915 146612 -165907
rect 146668 -165915 146712 -165907
rect 146768 -165915 146812 -165907
rect 147268 -165915 147312 -165907
rect 147368 -165915 147412 -165907
rect 147468 -165915 147512 -165907
rect 147568 -165915 147612 -165907
rect 147668 -165915 147712 -165907
rect 147768 -165915 147812 -165907
rect 147868 -165915 147912 -165907
rect 147968 -165915 148012 -165907
rect 148068 -165915 148112 -165907
rect 148168 -165915 148212 -165907
rect 148268 -165915 148312 -165907
rect 148368 -165915 148412 -165907
rect 148468 -165915 148512 -165907
rect 148568 -165915 148612 -165907
rect 148668 -165915 148712 -165907
rect 148768 -165915 148812 -165907
rect 149268 -165915 149312 -165907
rect 149368 -165915 149412 -165907
rect 149468 -165915 149512 -165907
rect 149568 -165915 149612 -165907
rect 149668 -165915 149712 -165907
rect 149768 -165915 149812 -165907
rect 149868 -165915 149912 -165907
rect 149968 -165915 150012 -165907
rect 150068 -165915 150112 -165907
rect 150168 -165915 150212 -165907
rect 150268 -165915 150312 -165907
rect 150368 -165915 150412 -165907
rect 150468 -165915 150512 -165907
rect 150568 -165915 150612 -165907
rect 150668 -165915 150712 -165907
rect 150768 -165915 150812 -165907
rect 151268 -165915 151312 -165907
rect 151368 -165915 151412 -165907
rect 151468 -165915 151512 -165907
rect 151568 -165915 151612 -165907
rect 151668 -165915 151712 -165907
rect 151768 -165915 151812 -165907
rect 151868 -165915 151912 -165907
rect 151968 -165915 152012 -165907
rect 152068 -165915 152112 -165907
rect 152168 -165915 152212 -165907
rect 152268 -165915 152312 -165907
rect 152368 -165915 152412 -165907
rect 152468 -165915 152512 -165907
rect 152568 -165915 152612 -165907
rect 152668 -165915 152712 -165907
rect 152768 -165915 152812 -165907
rect 145312 -165959 145320 -165915
rect 145412 -165959 145420 -165915
rect 145512 -165959 145520 -165915
rect 145612 -165959 145620 -165915
rect 145712 -165959 145720 -165915
rect 145812 -165959 145820 -165915
rect 145912 -165959 145920 -165915
rect 146012 -165959 146020 -165915
rect 146112 -165959 146120 -165915
rect 146212 -165959 146220 -165915
rect 146312 -165959 146320 -165915
rect 146412 -165959 146420 -165915
rect 146512 -165959 146520 -165915
rect 146612 -165959 146620 -165915
rect 146712 -165959 146720 -165915
rect 146812 -165959 146820 -165915
rect 147312 -165959 147320 -165915
rect 147412 -165959 147420 -165915
rect 147512 -165959 147520 -165915
rect 147612 -165959 147620 -165915
rect 147712 -165959 147720 -165915
rect 147812 -165959 147820 -165915
rect 147912 -165959 147920 -165915
rect 148012 -165959 148020 -165915
rect 148112 -165959 148120 -165915
rect 148212 -165959 148220 -165915
rect 148312 -165959 148320 -165915
rect 148412 -165959 148420 -165915
rect 148512 -165959 148520 -165915
rect 148612 -165959 148620 -165915
rect 148712 -165959 148720 -165915
rect 148812 -165959 148820 -165915
rect 149312 -165959 149320 -165915
rect 149412 -165959 149420 -165915
rect 149512 -165959 149520 -165915
rect 149612 -165959 149620 -165915
rect 149712 -165959 149720 -165915
rect 149812 -165959 149820 -165915
rect 149912 -165959 149920 -165915
rect 150012 -165959 150020 -165915
rect 150112 -165959 150120 -165915
rect 150212 -165959 150220 -165915
rect 150312 -165959 150320 -165915
rect 150412 -165959 150420 -165915
rect 150512 -165959 150520 -165915
rect 150612 -165959 150620 -165915
rect 150712 -165959 150720 -165915
rect 150812 -165959 150820 -165915
rect 151312 -165959 151320 -165915
rect 151412 -165959 151420 -165915
rect 151512 -165959 151520 -165915
rect 151612 -165959 151620 -165915
rect 151712 -165959 151720 -165915
rect 151812 -165959 151820 -165915
rect 151912 -165959 151920 -165915
rect 152012 -165959 152020 -165915
rect 152112 -165959 152120 -165915
rect 152212 -165959 152220 -165915
rect 152312 -165959 152320 -165915
rect 152412 -165959 152420 -165915
rect 152512 -165959 152520 -165915
rect 152612 -165959 152620 -165915
rect 152712 -165959 152720 -165915
rect 152812 -165959 152820 -165915
rect 145268 -166015 145312 -166007
rect 145368 -166015 145412 -166007
rect 145468 -166015 145512 -166007
rect 145568 -166015 145612 -166007
rect 145668 -166015 145712 -166007
rect 145768 -166015 145812 -166007
rect 145868 -166015 145912 -166007
rect 145968 -166015 146012 -166007
rect 146068 -166015 146112 -166007
rect 146168 -166015 146212 -166007
rect 146268 -166015 146312 -166007
rect 146368 -166015 146412 -166007
rect 146468 -166015 146512 -166007
rect 146568 -166015 146612 -166007
rect 146668 -166015 146712 -166007
rect 146768 -166015 146812 -166007
rect 147268 -166015 147312 -166007
rect 147368 -166015 147412 -166007
rect 147468 -166015 147512 -166007
rect 147568 -166015 147612 -166007
rect 147668 -166015 147712 -166007
rect 147768 -166015 147812 -166007
rect 147868 -166015 147912 -166007
rect 147968 -166015 148012 -166007
rect 148068 -166015 148112 -166007
rect 148168 -166015 148212 -166007
rect 148268 -166015 148312 -166007
rect 148368 -166015 148412 -166007
rect 148468 -166015 148512 -166007
rect 148568 -166015 148612 -166007
rect 148668 -166015 148712 -166007
rect 148768 -166015 148812 -166007
rect 149268 -166015 149312 -166007
rect 149368 -166015 149412 -166007
rect 149468 -166015 149512 -166007
rect 149568 -166015 149612 -166007
rect 149668 -166015 149712 -166007
rect 149768 -166015 149812 -166007
rect 149868 -166015 149912 -166007
rect 149968 -166015 150012 -166007
rect 150068 -166015 150112 -166007
rect 150168 -166015 150212 -166007
rect 150268 -166015 150312 -166007
rect 150368 -166015 150412 -166007
rect 150468 -166015 150512 -166007
rect 150568 -166015 150612 -166007
rect 150668 -166015 150712 -166007
rect 150768 -166015 150812 -166007
rect 151268 -166015 151312 -166007
rect 151368 -166015 151412 -166007
rect 151468 -166015 151512 -166007
rect 151568 -166015 151612 -166007
rect 151668 -166015 151712 -166007
rect 151768 -166015 151812 -166007
rect 151868 -166015 151912 -166007
rect 151968 -166015 152012 -166007
rect 152068 -166015 152112 -166007
rect 152168 -166015 152212 -166007
rect 152268 -166015 152312 -166007
rect 152368 -166015 152412 -166007
rect 152468 -166015 152512 -166007
rect 152568 -166015 152612 -166007
rect 152668 -166015 152712 -166007
rect 152768 -166015 152812 -166007
rect 145312 -166059 145320 -166015
rect 145412 -166059 145420 -166015
rect 145512 -166059 145520 -166015
rect 145612 -166059 145620 -166015
rect 145712 -166059 145720 -166015
rect 145812 -166059 145820 -166015
rect 145912 -166059 145920 -166015
rect 146012 -166059 146020 -166015
rect 146112 -166059 146120 -166015
rect 146212 -166059 146220 -166015
rect 146312 -166059 146320 -166015
rect 146412 -166059 146420 -166015
rect 146512 -166059 146520 -166015
rect 146612 -166059 146620 -166015
rect 146712 -166059 146720 -166015
rect 146812 -166059 146820 -166015
rect 147312 -166059 147320 -166015
rect 147412 -166059 147420 -166015
rect 147512 -166059 147520 -166015
rect 147612 -166059 147620 -166015
rect 147712 -166059 147720 -166015
rect 147812 -166059 147820 -166015
rect 147912 -166059 147920 -166015
rect 148012 -166059 148020 -166015
rect 148112 -166059 148120 -166015
rect 148212 -166059 148220 -166015
rect 148312 -166059 148320 -166015
rect 148412 -166059 148420 -166015
rect 148512 -166059 148520 -166015
rect 148612 -166059 148620 -166015
rect 148712 -166059 148720 -166015
rect 148812 -166059 148820 -166015
rect 149312 -166059 149320 -166015
rect 149412 -166059 149420 -166015
rect 149512 -166059 149520 -166015
rect 149612 -166059 149620 -166015
rect 149712 -166059 149720 -166015
rect 149812 -166059 149820 -166015
rect 149912 -166059 149920 -166015
rect 150012 -166059 150020 -166015
rect 150112 -166059 150120 -166015
rect 150212 -166059 150220 -166015
rect 150312 -166059 150320 -166015
rect 150412 -166059 150420 -166015
rect 150512 -166059 150520 -166015
rect 150612 -166059 150620 -166015
rect 150712 -166059 150720 -166015
rect 150812 -166059 150820 -166015
rect 151312 -166059 151320 -166015
rect 151412 -166059 151420 -166015
rect 151512 -166059 151520 -166015
rect 151612 -166059 151620 -166015
rect 151712 -166059 151720 -166015
rect 151812 -166059 151820 -166015
rect 151912 -166059 151920 -166015
rect 152012 -166059 152020 -166015
rect 152112 -166059 152120 -166015
rect 152212 -166059 152220 -166015
rect 152312 -166059 152320 -166015
rect 152412 -166059 152420 -166015
rect 152512 -166059 152520 -166015
rect 152612 -166059 152620 -166015
rect 152712 -166059 152720 -166015
rect 152812 -166059 152820 -166015
rect 145268 -166115 145312 -166107
rect 145368 -166115 145412 -166107
rect 145468 -166115 145512 -166107
rect 145568 -166115 145612 -166107
rect 145668 -166115 145712 -166107
rect 145768 -166115 145812 -166107
rect 145868 -166115 145912 -166107
rect 145968 -166115 146012 -166107
rect 146068 -166115 146112 -166107
rect 146168 -166115 146212 -166107
rect 146268 -166115 146312 -166107
rect 146368 -166115 146412 -166107
rect 146468 -166115 146512 -166107
rect 146568 -166115 146612 -166107
rect 146668 -166115 146712 -166107
rect 146768 -166115 146812 -166107
rect 147268 -166115 147312 -166107
rect 147368 -166115 147412 -166107
rect 147468 -166115 147512 -166107
rect 147568 -166115 147612 -166107
rect 147668 -166115 147712 -166107
rect 147768 -166115 147812 -166107
rect 147868 -166115 147912 -166107
rect 147968 -166115 148012 -166107
rect 148068 -166115 148112 -166107
rect 148168 -166115 148212 -166107
rect 148268 -166115 148312 -166107
rect 148368 -166115 148412 -166107
rect 148468 -166115 148512 -166107
rect 148568 -166115 148612 -166107
rect 148668 -166115 148712 -166107
rect 148768 -166115 148812 -166107
rect 149268 -166115 149312 -166107
rect 149368 -166115 149412 -166107
rect 149468 -166115 149512 -166107
rect 149568 -166115 149612 -166107
rect 149668 -166115 149712 -166107
rect 149768 -166115 149812 -166107
rect 149868 -166115 149912 -166107
rect 149968 -166115 150012 -166107
rect 150068 -166115 150112 -166107
rect 150168 -166115 150212 -166107
rect 150268 -166115 150312 -166107
rect 150368 -166115 150412 -166107
rect 150468 -166115 150512 -166107
rect 150568 -166115 150612 -166107
rect 150668 -166115 150712 -166107
rect 150768 -166115 150812 -166107
rect 151268 -166115 151312 -166107
rect 151368 -166115 151412 -166107
rect 151468 -166115 151512 -166107
rect 151568 -166115 151612 -166107
rect 151668 -166115 151712 -166107
rect 151768 -166115 151812 -166107
rect 151868 -166115 151912 -166107
rect 151968 -166115 152012 -166107
rect 152068 -166115 152112 -166107
rect 152168 -166115 152212 -166107
rect 152268 -166115 152312 -166107
rect 152368 -166115 152412 -166107
rect 152468 -166115 152512 -166107
rect 152568 -166115 152612 -166107
rect 152668 -166115 152712 -166107
rect 152768 -166115 152812 -166107
rect 145312 -166159 145320 -166115
rect 145412 -166159 145420 -166115
rect 145512 -166159 145520 -166115
rect 145612 -166159 145620 -166115
rect 145712 -166159 145720 -166115
rect 145812 -166159 145820 -166115
rect 145912 -166159 145920 -166115
rect 146012 -166159 146020 -166115
rect 146112 -166159 146120 -166115
rect 146212 -166159 146220 -166115
rect 146312 -166159 146320 -166115
rect 146412 -166159 146420 -166115
rect 146512 -166159 146520 -166115
rect 146612 -166159 146620 -166115
rect 146712 -166159 146720 -166115
rect 146812 -166159 146820 -166115
rect 147312 -166159 147320 -166115
rect 147412 -166159 147420 -166115
rect 147512 -166159 147520 -166115
rect 147612 -166159 147620 -166115
rect 147712 -166159 147720 -166115
rect 147812 -166159 147820 -166115
rect 147912 -166159 147920 -166115
rect 148012 -166159 148020 -166115
rect 148112 -166159 148120 -166115
rect 148212 -166159 148220 -166115
rect 148312 -166159 148320 -166115
rect 148412 -166159 148420 -166115
rect 148512 -166159 148520 -166115
rect 148612 -166159 148620 -166115
rect 148712 -166159 148720 -166115
rect 148812 -166159 148820 -166115
rect 149312 -166159 149320 -166115
rect 149412 -166159 149420 -166115
rect 149512 -166159 149520 -166115
rect 149612 -166159 149620 -166115
rect 149712 -166159 149720 -166115
rect 149812 -166159 149820 -166115
rect 149912 -166159 149920 -166115
rect 150012 -166159 150020 -166115
rect 150112 -166159 150120 -166115
rect 150212 -166159 150220 -166115
rect 150312 -166159 150320 -166115
rect 150412 -166159 150420 -166115
rect 150512 -166159 150520 -166115
rect 150612 -166159 150620 -166115
rect 150712 -166159 150720 -166115
rect 150812 -166159 150820 -166115
rect 151312 -166159 151320 -166115
rect 151412 -166159 151420 -166115
rect 151512 -166159 151520 -166115
rect 151612 -166159 151620 -166115
rect 151712 -166159 151720 -166115
rect 151812 -166159 151820 -166115
rect 151912 -166159 151920 -166115
rect 152012 -166159 152020 -166115
rect 152112 -166159 152120 -166115
rect 152212 -166159 152220 -166115
rect 152312 -166159 152320 -166115
rect 152412 -166159 152420 -166115
rect 152512 -166159 152520 -166115
rect 152612 -166159 152620 -166115
rect 152712 -166159 152720 -166115
rect 152812 -166159 152820 -166115
rect 145268 -166215 145312 -166207
rect 145368 -166215 145412 -166207
rect 145468 -166215 145512 -166207
rect 145568 -166215 145612 -166207
rect 145668 -166215 145712 -166207
rect 145768 -166215 145812 -166207
rect 145868 -166215 145912 -166207
rect 145968 -166215 146012 -166207
rect 146068 -166215 146112 -166207
rect 146168 -166215 146212 -166207
rect 146268 -166215 146312 -166207
rect 146368 -166215 146412 -166207
rect 146468 -166215 146512 -166207
rect 146568 -166215 146612 -166207
rect 146668 -166215 146712 -166207
rect 146768 -166215 146812 -166207
rect 147268 -166215 147312 -166207
rect 147368 -166215 147412 -166207
rect 147468 -166215 147512 -166207
rect 147568 -166215 147612 -166207
rect 147668 -166215 147712 -166207
rect 147768 -166215 147812 -166207
rect 147868 -166215 147912 -166207
rect 147968 -166215 148012 -166207
rect 148068 -166215 148112 -166207
rect 148168 -166215 148212 -166207
rect 148268 -166215 148312 -166207
rect 148368 -166215 148412 -166207
rect 148468 -166215 148512 -166207
rect 148568 -166215 148612 -166207
rect 148668 -166215 148712 -166207
rect 148768 -166215 148812 -166207
rect 149268 -166215 149312 -166207
rect 149368 -166215 149412 -166207
rect 149468 -166215 149512 -166207
rect 149568 -166215 149612 -166207
rect 149668 -166215 149712 -166207
rect 149768 -166215 149812 -166207
rect 149868 -166215 149912 -166207
rect 149968 -166215 150012 -166207
rect 150068 -166215 150112 -166207
rect 150168 -166215 150212 -166207
rect 150268 -166215 150312 -166207
rect 150368 -166215 150412 -166207
rect 150468 -166215 150512 -166207
rect 150568 -166215 150612 -166207
rect 150668 -166215 150712 -166207
rect 150768 -166215 150812 -166207
rect 151268 -166215 151312 -166207
rect 151368 -166215 151412 -166207
rect 151468 -166215 151512 -166207
rect 151568 -166215 151612 -166207
rect 151668 -166215 151712 -166207
rect 151768 -166215 151812 -166207
rect 151868 -166215 151912 -166207
rect 151968 -166215 152012 -166207
rect 152068 -166215 152112 -166207
rect 152168 -166215 152212 -166207
rect 152268 -166215 152312 -166207
rect 152368 -166215 152412 -166207
rect 152468 -166215 152512 -166207
rect 152568 -166215 152612 -166207
rect 152668 -166215 152712 -166207
rect 152768 -166215 152812 -166207
rect 145312 -166259 145320 -166215
rect 145412 -166259 145420 -166215
rect 145512 -166259 145520 -166215
rect 145612 -166259 145620 -166215
rect 145712 -166259 145720 -166215
rect 145812 -166259 145820 -166215
rect 145912 -166259 145920 -166215
rect 146012 -166259 146020 -166215
rect 146112 -166259 146120 -166215
rect 146212 -166259 146220 -166215
rect 146312 -166259 146320 -166215
rect 146412 -166259 146420 -166215
rect 146512 -166259 146520 -166215
rect 146612 -166259 146620 -166215
rect 146712 -166259 146720 -166215
rect 146812 -166259 146820 -166215
rect 147312 -166259 147320 -166215
rect 147412 -166259 147420 -166215
rect 147512 -166259 147520 -166215
rect 147612 -166259 147620 -166215
rect 147712 -166259 147720 -166215
rect 147812 -166259 147820 -166215
rect 147912 -166259 147920 -166215
rect 148012 -166259 148020 -166215
rect 148112 -166259 148120 -166215
rect 148212 -166259 148220 -166215
rect 148312 -166259 148320 -166215
rect 148412 -166259 148420 -166215
rect 148512 -166259 148520 -166215
rect 148612 -166259 148620 -166215
rect 148712 -166259 148720 -166215
rect 148812 -166259 148820 -166215
rect 149312 -166259 149320 -166215
rect 149412 -166259 149420 -166215
rect 149512 -166259 149520 -166215
rect 149612 -166259 149620 -166215
rect 149712 -166259 149720 -166215
rect 149812 -166259 149820 -166215
rect 149912 -166259 149920 -166215
rect 150012 -166259 150020 -166215
rect 150112 -166259 150120 -166215
rect 150212 -166259 150220 -166215
rect 150312 -166259 150320 -166215
rect 150412 -166259 150420 -166215
rect 150512 -166259 150520 -166215
rect 150612 -166259 150620 -166215
rect 150712 -166259 150720 -166215
rect 150812 -166259 150820 -166215
rect 151312 -166259 151320 -166215
rect 151412 -166259 151420 -166215
rect 151512 -166259 151520 -166215
rect 151612 -166259 151620 -166215
rect 151712 -166259 151720 -166215
rect 151812 -166259 151820 -166215
rect 151912 -166259 151920 -166215
rect 152012 -166259 152020 -166215
rect 152112 -166259 152120 -166215
rect 152212 -166259 152220 -166215
rect 152312 -166259 152320 -166215
rect 152412 -166259 152420 -166215
rect 152512 -166259 152520 -166215
rect 152612 -166259 152620 -166215
rect 152712 -166259 152720 -166215
rect 152812 -166259 152820 -166215
rect 145268 -166315 145312 -166307
rect 145368 -166315 145412 -166307
rect 145468 -166315 145512 -166307
rect 145568 -166315 145612 -166307
rect 145668 -166315 145712 -166307
rect 145768 -166315 145812 -166307
rect 145868 -166315 145912 -166307
rect 145968 -166315 146012 -166307
rect 146068 -166315 146112 -166307
rect 146168 -166315 146212 -166307
rect 146268 -166315 146312 -166307
rect 146368 -166315 146412 -166307
rect 146468 -166315 146512 -166307
rect 146568 -166315 146612 -166307
rect 146668 -166315 146712 -166307
rect 146768 -166315 146812 -166307
rect 147268 -166315 147312 -166307
rect 147368 -166315 147412 -166307
rect 147468 -166315 147512 -166307
rect 147568 -166315 147612 -166307
rect 147668 -166315 147712 -166307
rect 147768 -166315 147812 -166307
rect 147868 -166315 147912 -166307
rect 147968 -166315 148012 -166307
rect 148068 -166315 148112 -166307
rect 148168 -166315 148212 -166307
rect 148268 -166315 148312 -166307
rect 148368 -166315 148412 -166307
rect 148468 -166315 148512 -166307
rect 148568 -166315 148612 -166307
rect 148668 -166315 148712 -166307
rect 148768 -166315 148812 -166307
rect 149268 -166315 149312 -166307
rect 149368 -166315 149412 -166307
rect 149468 -166315 149512 -166307
rect 149568 -166315 149612 -166307
rect 149668 -166315 149712 -166307
rect 149768 -166315 149812 -166307
rect 149868 -166315 149912 -166307
rect 149968 -166315 150012 -166307
rect 150068 -166315 150112 -166307
rect 150168 -166315 150212 -166307
rect 150268 -166315 150312 -166307
rect 150368 -166315 150412 -166307
rect 150468 -166315 150512 -166307
rect 150568 -166315 150612 -166307
rect 150668 -166315 150712 -166307
rect 150768 -166315 150812 -166307
rect 151268 -166315 151312 -166307
rect 151368 -166315 151412 -166307
rect 151468 -166315 151512 -166307
rect 151568 -166315 151612 -166307
rect 151668 -166315 151712 -166307
rect 151768 -166315 151812 -166307
rect 151868 -166315 151912 -166307
rect 151968 -166315 152012 -166307
rect 152068 -166315 152112 -166307
rect 152168 -166315 152212 -166307
rect 152268 -166315 152312 -166307
rect 152368 -166315 152412 -166307
rect 152468 -166315 152512 -166307
rect 152568 -166315 152612 -166307
rect 152668 -166315 152712 -166307
rect 152768 -166315 152812 -166307
rect 145312 -166359 145320 -166315
rect 145412 -166359 145420 -166315
rect 145512 -166359 145520 -166315
rect 145612 -166359 145620 -166315
rect 145712 -166359 145720 -166315
rect 145812 -166359 145820 -166315
rect 145912 -166359 145920 -166315
rect 146012 -166359 146020 -166315
rect 146112 -166359 146120 -166315
rect 146212 -166359 146220 -166315
rect 146312 -166359 146320 -166315
rect 146412 -166359 146420 -166315
rect 146512 -166359 146520 -166315
rect 146612 -166359 146620 -166315
rect 146712 -166359 146720 -166315
rect 146812 -166359 146820 -166315
rect 147312 -166359 147320 -166315
rect 147412 -166359 147420 -166315
rect 147512 -166359 147520 -166315
rect 147612 -166359 147620 -166315
rect 147712 -166359 147720 -166315
rect 147812 -166359 147820 -166315
rect 147912 -166359 147920 -166315
rect 148012 -166359 148020 -166315
rect 148112 -166359 148120 -166315
rect 148212 -166359 148220 -166315
rect 148312 -166359 148320 -166315
rect 148412 -166359 148420 -166315
rect 148512 -166359 148520 -166315
rect 148612 -166359 148620 -166315
rect 148712 -166359 148720 -166315
rect 148812 -166359 148820 -166315
rect 149312 -166359 149320 -166315
rect 149412 -166359 149420 -166315
rect 149512 -166359 149520 -166315
rect 149612 -166359 149620 -166315
rect 149712 -166359 149720 -166315
rect 149812 -166359 149820 -166315
rect 149912 -166359 149920 -166315
rect 150012 -166359 150020 -166315
rect 150112 -166359 150120 -166315
rect 150212 -166359 150220 -166315
rect 150312 -166359 150320 -166315
rect 150412 -166359 150420 -166315
rect 150512 -166359 150520 -166315
rect 150612 -166359 150620 -166315
rect 150712 -166359 150720 -166315
rect 150812 -166359 150820 -166315
rect 151312 -166359 151320 -166315
rect 151412 -166359 151420 -166315
rect 151512 -166359 151520 -166315
rect 151612 -166359 151620 -166315
rect 151712 -166359 151720 -166315
rect 151812 -166359 151820 -166315
rect 151912 -166359 151920 -166315
rect 152012 -166359 152020 -166315
rect 152112 -166359 152120 -166315
rect 152212 -166359 152220 -166315
rect 152312 -166359 152320 -166315
rect 152412 -166359 152420 -166315
rect 152512 -166359 152520 -166315
rect 152612 -166359 152620 -166315
rect 152712 -166359 152720 -166315
rect 152812 -166359 152820 -166315
rect 145268 -166415 145312 -166407
rect 145368 -166415 145412 -166407
rect 145468 -166415 145512 -166407
rect 145568 -166415 145612 -166407
rect 145668 -166415 145712 -166407
rect 145768 -166415 145812 -166407
rect 145868 -166415 145912 -166407
rect 145968 -166415 146012 -166407
rect 146068 -166415 146112 -166407
rect 146168 -166415 146212 -166407
rect 146268 -166415 146312 -166407
rect 146368 -166415 146412 -166407
rect 146468 -166415 146512 -166407
rect 146568 -166415 146612 -166407
rect 146668 -166415 146712 -166407
rect 146768 -166415 146812 -166407
rect 147268 -166415 147312 -166407
rect 147368 -166415 147412 -166407
rect 147468 -166415 147512 -166407
rect 147568 -166415 147612 -166407
rect 147668 -166415 147712 -166407
rect 147768 -166415 147812 -166407
rect 147868 -166415 147912 -166407
rect 147968 -166415 148012 -166407
rect 148068 -166415 148112 -166407
rect 148168 -166415 148212 -166407
rect 148268 -166415 148312 -166407
rect 148368 -166415 148412 -166407
rect 148468 -166415 148512 -166407
rect 148568 -166415 148612 -166407
rect 148668 -166415 148712 -166407
rect 148768 -166415 148812 -166407
rect 149268 -166415 149312 -166407
rect 149368 -166415 149412 -166407
rect 149468 -166415 149512 -166407
rect 149568 -166415 149612 -166407
rect 149668 -166415 149712 -166407
rect 149768 -166415 149812 -166407
rect 149868 -166415 149912 -166407
rect 149968 -166415 150012 -166407
rect 150068 -166415 150112 -166407
rect 150168 -166415 150212 -166407
rect 150268 -166415 150312 -166407
rect 150368 -166415 150412 -166407
rect 150468 -166415 150512 -166407
rect 150568 -166415 150612 -166407
rect 150668 -166415 150712 -166407
rect 150768 -166415 150812 -166407
rect 151268 -166415 151312 -166407
rect 151368 -166415 151412 -166407
rect 151468 -166415 151512 -166407
rect 151568 -166415 151612 -166407
rect 151668 -166415 151712 -166407
rect 151768 -166415 151812 -166407
rect 151868 -166415 151912 -166407
rect 151968 -166415 152012 -166407
rect 152068 -166415 152112 -166407
rect 152168 -166415 152212 -166407
rect 152268 -166415 152312 -166407
rect 152368 -166415 152412 -166407
rect 152468 -166415 152512 -166407
rect 152568 -166415 152612 -166407
rect 152668 -166415 152712 -166407
rect 152768 -166415 152812 -166407
rect 145312 -166459 145320 -166415
rect 145412 -166459 145420 -166415
rect 145512 -166459 145520 -166415
rect 145612 -166459 145620 -166415
rect 145712 -166459 145720 -166415
rect 145812 -166459 145820 -166415
rect 145912 -166459 145920 -166415
rect 146012 -166459 146020 -166415
rect 146112 -166459 146120 -166415
rect 146212 -166459 146220 -166415
rect 146312 -166459 146320 -166415
rect 146412 -166459 146420 -166415
rect 146512 -166459 146520 -166415
rect 146612 -166459 146620 -166415
rect 146712 -166459 146720 -166415
rect 146812 -166459 146820 -166415
rect 147312 -166459 147320 -166415
rect 147412 -166459 147420 -166415
rect 147512 -166459 147520 -166415
rect 147612 -166459 147620 -166415
rect 147712 -166459 147720 -166415
rect 147812 -166459 147820 -166415
rect 147912 -166459 147920 -166415
rect 148012 -166459 148020 -166415
rect 148112 -166459 148120 -166415
rect 148212 -166459 148220 -166415
rect 148312 -166459 148320 -166415
rect 148412 -166459 148420 -166415
rect 148512 -166459 148520 -166415
rect 148612 -166459 148620 -166415
rect 148712 -166459 148720 -166415
rect 148812 -166459 148820 -166415
rect 149312 -166459 149320 -166415
rect 149412 -166459 149420 -166415
rect 149512 -166459 149520 -166415
rect 149612 -166459 149620 -166415
rect 149712 -166459 149720 -166415
rect 149812 -166459 149820 -166415
rect 149912 -166459 149920 -166415
rect 150012 -166459 150020 -166415
rect 150112 -166459 150120 -166415
rect 150212 -166459 150220 -166415
rect 150312 -166459 150320 -166415
rect 150412 -166459 150420 -166415
rect 150512 -166459 150520 -166415
rect 150612 -166459 150620 -166415
rect 150712 -166459 150720 -166415
rect 150812 -166459 150820 -166415
rect 151312 -166459 151320 -166415
rect 151412 -166459 151420 -166415
rect 151512 -166459 151520 -166415
rect 151612 -166459 151620 -166415
rect 151712 -166459 151720 -166415
rect 151812 -166459 151820 -166415
rect 151912 -166459 151920 -166415
rect 152012 -166459 152020 -166415
rect 152112 -166459 152120 -166415
rect 152212 -166459 152220 -166415
rect 152312 -166459 152320 -166415
rect 152412 -166459 152420 -166415
rect 152512 -166459 152520 -166415
rect 152612 -166459 152620 -166415
rect 152712 -166459 152720 -166415
rect 152812 -166459 152820 -166415
rect 145268 -166515 145312 -166507
rect 145368 -166515 145412 -166507
rect 145468 -166515 145512 -166507
rect 145568 -166515 145612 -166507
rect 145668 -166515 145712 -166507
rect 145768 -166515 145812 -166507
rect 145868 -166515 145912 -166507
rect 145968 -166515 146012 -166507
rect 146068 -166515 146112 -166507
rect 146168 -166515 146212 -166507
rect 146268 -166515 146312 -166507
rect 146368 -166515 146412 -166507
rect 146468 -166515 146512 -166507
rect 146568 -166515 146612 -166507
rect 146668 -166515 146712 -166507
rect 146768 -166515 146812 -166507
rect 147268 -166515 147312 -166507
rect 147368 -166515 147412 -166507
rect 147468 -166515 147512 -166507
rect 147568 -166515 147612 -166507
rect 147668 -166515 147712 -166507
rect 147768 -166515 147812 -166507
rect 147868 -166515 147912 -166507
rect 147968 -166515 148012 -166507
rect 148068 -166515 148112 -166507
rect 148168 -166515 148212 -166507
rect 148268 -166515 148312 -166507
rect 148368 -166515 148412 -166507
rect 148468 -166515 148512 -166507
rect 148568 -166515 148612 -166507
rect 148668 -166515 148712 -166507
rect 148768 -166515 148812 -166507
rect 149268 -166515 149312 -166507
rect 149368 -166515 149412 -166507
rect 149468 -166515 149512 -166507
rect 149568 -166515 149612 -166507
rect 149668 -166515 149712 -166507
rect 149768 -166515 149812 -166507
rect 149868 -166515 149912 -166507
rect 149968 -166515 150012 -166507
rect 150068 -166515 150112 -166507
rect 150168 -166515 150212 -166507
rect 150268 -166515 150312 -166507
rect 150368 -166515 150412 -166507
rect 150468 -166515 150512 -166507
rect 150568 -166515 150612 -166507
rect 150668 -166515 150712 -166507
rect 150768 -166515 150812 -166507
rect 151268 -166515 151312 -166507
rect 151368 -166515 151412 -166507
rect 151468 -166515 151512 -166507
rect 151568 -166515 151612 -166507
rect 151668 -166515 151712 -166507
rect 151768 -166515 151812 -166507
rect 151868 -166515 151912 -166507
rect 151968 -166515 152012 -166507
rect 152068 -166515 152112 -166507
rect 152168 -166515 152212 -166507
rect 152268 -166515 152312 -166507
rect 152368 -166515 152412 -166507
rect 152468 -166515 152512 -166507
rect 152568 -166515 152612 -166507
rect 152668 -166515 152712 -166507
rect 152768 -166515 152812 -166507
rect 145312 -166559 145320 -166515
rect 145412 -166559 145420 -166515
rect 145512 -166559 145520 -166515
rect 145612 -166559 145620 -166515
rect 145712 -166559 145720 -166515
rect 145812 -166559 145820 -166515
rect 145912 -166559 145920 -166515
rect 146012 -166559 146020 -166515
rect 146112 -166559 146120 -166515
rect 146212 -166559 146220 -166515
rect 146312 -166559 146320 -166515
rect 146412 -166559 146420 -166515
rect 146512 -166559 146520 -166515
rect 146612 -166559 146620 -166515
rect 146712 -166559 146720 -166515
rect 146812 -166559 146820 -166515
rect 147312 -166559 147320 -166515
rect 147412 -166559 147420 -166515
rect 147512 -166559 147520 -166515
rect 147612 -166559 147620 -166515
rect 147712 -166559 147720 -166515
rect 147812 -166559 147820 -166515
rect 147912 -166559 147920 -166515
rect 148012 -166559 148020 -166515
rect 148112 -166559 148120 -166515
rect 148212 -166559 148220 -166515
rect 148312 -166559 148320 -166515
rect 148412 -166559 148420 -166515
rect 148512 -166559 148520 -166515
rect 148612 -166559 148620 -166515
rect 148712 -166559 148720 -166515
rect 148812 -166559 148820 -166515
rect 149312 -166559 149320 -166515
rect 149412 -166559 149420 -166515
rect 149512 -166559 149520 -166515
rect 149612 -166559 149620 -166515
rect 149712 -166559 149720 -166515
rect 149812 -166559 149820 -166515
rect 149912 -166559 149920 -166515
rect 150012 -166559 150020 -166515
rect 150112 -166559 150120 -166515
rect 150212 -166559 150220 -166515
rect 150312 -166559 150320 -166515
rect 150412 -166559 150420 -166515
rect 150512 -166559 150520 -166515
rect 150612 -166559 150620 -166515
rect 150712 -166559 150720 -166515
rect 150812 -166559 150820 -166515
rect 151312 -166559 151320 -166515
rect 151412 -166559 151420 -166515
rect 151512 -166559 151520 -166515
rect 151612 -166559 151620 -166515
rect 151712 -166559 151720 -166515
rect 151812 -166559 151820 -166515
rect 151912 -166559 151920 -166515
rect 152012 -166559 152020 -166515
rect 152112 -166559 152120 -166515
rect 152212 -166559 152220 -166515
rect 152312 -166559 152320 -166515
rect 152412 -166559 152420 -166515
rect 152512 -166559 152520 -166515
rect 152612 -166559 152620 -166515
rect 152712 -166559 152720 -166515
rect 152812 -166559 152820 -166515
rect 145268 -166615 145312 -166607
rect 145368 -166615 145412 -166607
rect 145468 -166615 145512 -166607
rect 145568 -166615 145612 -166607
rect 145668 -166615 145712 -166607
rect 145768 -166615 145812 -166607
rect 145868 -166615 145912 -166607
rect 145968 -166615 146012 -166607
rect 146068 -166615 146112 -166607
rect 146168 -166615 146212 -166607
rect 146268 -166615 146312 -166607
rect 146368 -166615 146412 -166607
rect 146468 -166615 146512 -166607
rect 146568 -166615 146612 -166607
rect 146668 -166615 146712 -166607
rect 146768 -166615 146812 -166607
rect 147268 -166615 147312 -166607
rect 147368 -166615 147412 -166607
rect 147468 -166615 147512 -166607
rect 147568 -166615 147612 -166607
rect 147668 -166615 147712 -166607
rect 147768 -166615 147812 -166607
rect 147868 -166615 147912 -166607
rect 147968 -166615 148012 -166607
rect 148068 -166615 148112 -166607
rect 148168 -166615 148212 -166607
rect 148268 -166615 148312 -166607
rect 148368 -166615 148412 -166607
rect 148468 -166615 148512 -166607
rect 148568 -166615 148612 -166607
rect 148668 -166615 148712 -166607
rect 148768 -166615 148812 -166607
rect 149268 -166615 149312 -166607
rect 149368 -166615 149412 -166607
rect 149468 -166615 149512 -166607
rect 149568 -166615 149612 -166607
rect 149668 -166615 149712 -166607
rect 149768 -166615 149812 -166607
rect 149868 -166615 149912 -166607
rect 149968 -166615 150012 -166607
rect 150068 -166615 150112 -166607
rect 150168 -166615 150212 -166607
rect 150268 -166615 150312 -166607
rect 150368 -166615 150412 -166607
rect 150468 -166615 150512 -166607
rect 150568 -166615 150612 -166607
rect 150668 -166615 150712 -166607
rect 150768 -166615 150812 -166607
rect 151268 -166615 151312 -166607
rect 151368 -166615 151412 -166607
rect 151468 -166615 151512 -166607
rect 151568 -166615 151612 -166607
rect 151668 -166615 151712 -166607
rect 151768 -166615 151812 -166607
rect 151868 -166615 151912 -166607
rect 151968 -166615 152012 -166607
rect 152068 -166615 152112 -166607
rect 152168 -166615 152212 -166607
rect 152268 -166615 152312 -166607
rect 152368 -166615 152412 -166607
rect 152468 -166615 152512 -166607
rect 152568 -166615 152612 -166607
rect 152668 -166615 152712 -166607
rect 152768 -166615 152812 -166607
rect 145312 -166659 145320 -166615
rect 145412 -166659 145420 -166615
rect 145512 -166659 145520 -166615
rect 145612 -166659 145620 -166615
rect 145712 -166659 145720 -166615
rect 145812 -166659 145820 -166615
rect 145912 -166659 145920 -166615
rect 146012 -166659 146020 -166615
rect 146112 -166659 146120 -166615
rect 146212 -166659 146220 -166615
rect 146312 -166659 146320 -166615
rect 146412 -166659 146420 -166615
rect 146512 -166659 146520 -166615
rect 146612 -166659 146620 -166615
rect 146712 -166659 146720 -166615
rect 146812 -166659 146820 -166615
rect 147312 -166659 147320 -166615
rect 147412 -166659 147420 -166615
rect 147512 -166659 147520 -166615
rect 147612 -166659 147620 -166615
rect 147712 -166659 147720 -166615
rect 147812 -166659 147820 -166615
rect 147912 -166659 147920 -166615
rect 148012 -166659 148020 -166615
rect 148112 -166659 148120 -166615
rect 148212 -166659 148220 -166615
rect 148312 -166659 148320 -166615
rect 148412 -166659 148420 -166615
rect 148512 -166659 148520 -166615
rect 148612 -166659 148620 -166615
rect 148712 -166659 148720 -166615
rect 148812 -166659 148820 -166615
rect 149312 -166659 149320 -166615
rect 149412 -166659 149420 -166615
rect 149512 -166659 149520 -166615
rect 149612 -166659 149620 -166615
rect 149712 -166659 149720 -166615
rect 149812 -166659 149820 -166615
rect 149912 -166659 149920 -166615
rect 150012 -166659 150020 -166615
rect 150112 -166659 150120 -166615
rect 150212 -166659 150220 -166615
rect 150312 -166659 150320 -166615
rect 150412 -166659 150420 -166615
rect 150512 -166659 150520 -166615
rect 150612 -166659 150620 -166615
rect 150712 -166659 150720 -166615
rect 150812 -166659 150820 -166615
rect 151312 -166659 151320 -166615
rect 151412 -166659 151420 -166615
rect 151512 -166659 151520 -166615
rect 151612 -166659 151620 -166615
rect 151712 -166659 151720 -166615
rect 151812 -166659 151820 -166615
rect 151912 -166659 151920 -166615
rect 152012 -166659 152020 -166615
rect 152112 -166659 152120 -166615
rect 152212 -166659 152220 -166615
rect 152312 -166659 152320 -166615
rect 152412 -166659 152420 -166615
rect 152512 -166659 152520 -166615
rect 152612 -166659 152620 -166615
rect 152712 -166659 152720 -166615
rect 152812 -166659 152820 -166615
rect 145268 -166715 145312 -166707
rect 145368 -166715 145412 -166707
rect 145468 -166715 145512 -166707
rect 145568 -166715 145612 -166707
rect 145668 -166715 145712 -166707
rect 145768 -166715 145812 -166707
rect 145868 -166715 145912 -166707
rect 145968 -166715 146012 -166707
rect 146068 -166715 146112 -166707
rect 146168 -166715 146212 -166707
rect 146268 -166715 146312 -166707
rect 146368 -166715 146412 -166707
rect 146468 -166715 146512 -166707
rect 146568 -166715 146612 -166707
rect 146668 -166715 146712 -166707
rect 146768 -166715 146812 -166707
rect 147268 -166715 147312 -166707
rect 147368 -166715 147412 -166707
rect 147468 -166715 147512 -166707
rect 147568 -166715 147612 -166707
rect 147668 -166715 147712 -166707
rect 147768 -166715 147812 -166707
rect 147868 -166715 147912 -166707
rect 147968 -166715 148012 -166707
rect 148068 -166715 148112 -166707
rect 148168 -166715 148212 -166707
rect 148268 -166715 148312 -166707
rect 148368 -166715 148412 -166707
rect 148468 -166715 148512 -166707
rect 148568 -166715 148612 -166707
rect 148668 -166715 148712 -166707
rect 148768 -166715 148812 -166707
rect 149268 -166715 149312 -166707
rect 149368 -166715 149412 -166707
rect 149468 -166715 149512 -166707
rect 149568 -166715 149612 -166707
rect 149668 -166715 149712 -166707
rect 149768 -166715 149812 -166707
rect 149868 -166715 149912 -166707
rect 149968 -166715 150012 -166707
rect 150068 -166715 150112 -166707
rect 150168 -166715 150212 -166707
rect 150268 -166715 150312 -166707
rect 150368 -166715 150412 -166707
rect 150468 -166715 150512 -166707
rect 150568 -166715 150612 -166707
rect 150668 -166715 150712 -166707
rect 150768 -166715 150812 -166707
rect 151268 -166715 151312 -166707
rect 151368 -166715 151412 -166707
rect 151468 -166715 151512 -166707
rect 151568 -166715 151612 -166707
rect 151668 -166715 151712 -166707
rect 151768 -166715 151812 -166707
rect 151868 -166715 151912 -166707
rect 151968 -166715 152012 -166707
rect 152068 -166715 152112 -166707
rect 152168 -166715 152212 -166707
rect 152268 -166715 152312 -166707
rect 152368 -166715 152412 -166707
rect 152468 -166715 152512 -166707
rect 152568 -166715 152612 -166707
rect 152668 -166715 152712 -166707
rect 152768 -166715 152812 -166707
rect 145312 -166759 145320 -166715
rect 145412 -166759 145420 -166715
rect 145512 -166759 145520 -166715
rect 145612 -166759 145620 -166715
rect 145712 -166759 145720 -166715
rect 145812 -166759 145820 -166715
rect 145912 -166759 145920 -166715
rect 146012 -166759 146020 -166715
rect 146112 -166759 146120 -166715
rect 146212 -166759 146220 -166715
rect 146312 -166759 146320 -166715
rect 146412 -166759 146420 -166715
rect 146512 -166759 146520 -166715
rect 146612 -166759 146620 -166715
rect 146712 -166759 146720 -166715
rect 146812 -166759 146820 -166715
rect 147312 -166759 147320 -166715
rect 147412 -166759 147420 -166715
rect 147512 -166759 147520 -166715
rect 147612 -166759 147620 -166715
rect 147712 -166759 147720 -166715
rect 147812 -166759 147820 -166715
rect 147912 -166759 147920 -166715
rect 148012 -166759 148020 -166715
rect 148112 -166759 148120 -166715
rect 148212 -166759 148220 -166715
rect 148312 -166759 148320 -166715
rect 148412 -166759 148420 -166715
rect 148512 -166759 148520 -166715
rect 148612 -166759 148620 -166715
rect 148712 -166759 148720 -166715
rect 148812 -166759 148820 -166715
rect 149312 -166759 149320 -166715
rect 149412 -166759 149420 -166715
rect 149512 -166759 149520 -166715
rect 149612 -166759 149620 -166715
rect 149712 -166759 149720 -166715
rect 149812 -166759 149820 -166715
rect 149912 -166759 149920 -166715
rect 150012 -166759 150020 -166715
rect 150112 -166759 150120 -166715
rect 150212 -166759 150220 -166715
rect 150312 -166759 150320 -166715
rect 150412 -166759 150420 -166715
rect 150512 -166759 150520 -166715
rect 150612 -166759 150620 -166715
rect 150712 -166759 150720 -166715
rect 150812 -166759 150820 -166715
rect 151312 -166759 151320 -166715
rect 151412 -166759 151420 -166715
rect 151512 -166759 151520 -166715
rect 151612 -166759 151620 -166715
rect 151712 -166759 151720 -166715
rect 151812 -166759 151820 -166715
rect 151912 -166759 151920 -166715
rect 152012 -166759 152020 -166715
rect 152112 -166759 152120 -166715
rect 152212 -166759 152220 -166715
rect 152312 -166759 152320 -166715
rect 152412 -166759 152420 -166715
rect 152512 -166759 152520 -166715
rect 152612 -166759 152620 -166715
rect 152712 -166759 152720 -166715
rect 152812 -166759 152820 -166715
rect 145268 -166815 145312 -166807
rect 145368 -166815 145412 -166807
rect 145468 -166815 145512 -166807
rect 145568 -166815 145612 -166807
rect 145668 -166815 145712 -166807
rect 145768 -166815 145812 -166807
rect 145868 -166815 145912 -166807
rect 145968 -166815 146012 -166807
rect 146068 -166815 146112 -166807
rect 146168 -166815 146212 -166807
rect 146268 -166815 146312 -166807
rect 146368 -166815 146412 -166807
rect 146468 -166815 146512 -166807
rect 146568 -166815 146612 -166807
rect 146668 -166815 146712 -166807
rect 146768 -166815 146812 -166807
rect 147268 -166815 147312 -166807
rect 147368 -166815 147412 -166807
rect 147468 -166815 147512 -166807
rect 147568 -166815 147612 -166807
rect 147668 -166815 147712 -166807
rect 147768 -166815 147812 -166807
rect 147868 -166815 147912 -166807
rect 147968 -166815 148012 -166807
rect 148068 -166815 148112 -166807
rect 148168 -166815 148212 -166807
rect 148268 -166815 148312 -166807
rect 148368 -166815 148412 -166807
rect 148468 -166815 148512 -166807
rect 148568 -166815 148612 -166807
rect 148668 -166815 148712 -166807
rect 148768 -166815 148812 -166807
rect 149268 -166815 149312 -166807
rect 149368 -166815 149412 -166807
rect 149468 -166815 149512 -166807
rect 149568 -166815 149612 -166807
rect 149668 -166815 149712 -166807
rect 149768 -166815 149812 -166807
rect 149868 -166815 149912 -166807
rect 149968 -166815 150012 -166807
rect 150068 -166815 150112 -166807
rect 150168 -166815 150212 -166807
rect 150268 -166815 150312 -166807
rect 150368 -166815 150412 -166807
rect 150468 -166815 150512 -166807
rect 150568 -166815 150612 -166807
rect 150668 -166815 150712 -166807
rect 150768 -166815 150812 -166807
rect 151268 -166815 151312 -166807
rect 151368 -166815 151412 -166807
rect 151468 -166815 151512 -166807
rect 151568 -166815 151612 -166807
rect 151668 -166815 151712 -166807
rect 151768 -166815 151812 -166807
rect 151868 -166815 151912 -166807
rect 151968 -166815 152012 -166807
rect 152068 -166815 152112 -166807
rect 152168 -166815 152212 -166807
rect 152268 -166815 152312 -166807
rect 152368 -166815 152412 -166807
rect 152468 -166815 152512 -166807
rect 152568 -166815 152612 -166807
rect 152668 -166815 152712 -166807
rect 152768 -166815 152812 -166807
rect 145312 -166859 145320 -166815
rect 145412 -166859 145420 -166815
rect 145512 -166859 145520 -166815
rect 145612 -166859 145620 -166815
rect 145712 -166859 145720 -166815
rect 145812 -166859 145820 -166815
rect 145912 -166859 145920 -166815
rect 146012 -166859 146020 -166815
rect 146112 -166859 146120 -166815
rect 146212 -166859 146220 -166815
rect 146312 -166859 146320 -166815
rect 146412 -166859 146420 -166815
rect 146512 -166859 146520 -166815
rect 146612 -166859 146620 -166815
rect 146712 -166859 146720 -166815
rect 146812 -166859 146820 -166815
rect 147312 -166859 147320 -166815
rect 147412 -166859 147420 -166815
rect 147512 -166859 147520 -166815
rect 147612 -166859 147620 -166815
rect 147712 -166859 147720 -166815
rect 147812 -166859 147820 -166815
rect 147912 -166859 147920 -166815
rect 148012 -166859 148020 -166815
rect 148112 -166859 148120 -166815
rect 148212 -166859 148220 -166815
rect 148312 -166859 148320 -166815
rect 148412 -166859 148420 -166815
rect 148512 -166859 148520 -166815
rect 148612 -166859 148620 -166815
rect 148712 -166859 148720 -166815
rect 148812 -166859 148820 -166815
rect 149312 -166859 149320 -166815
rect 149412 -166859 149420 -166815
rect 149512 -166859 149520 -166815
rect 149612 -166859 149620 -166815
rect 149712 -166859 149720 -166815
rect 149812 -166859 149820 -166815
rect 149912 -166859 149920 -166815
rect 150012 -166859 150020 -166815
rect 150112 -166859 150120 -166815
rect 150212 -166859 150220 -166815
rect 150312 -166859 150320 -166815
rect 150412 -166859 150420 -166815
rect 150512 -166859 150520 -166815
rect 150612 -166859 150620 -166815
rect 150712 -166859 150720 -166815
rect 150812 -166859 150820 -166815
rect 151312 -166859 151320 -166815
rect 151412 -166859 151420 -166815
rect 151512 -166859 151520 -166815
rect 151612 -166859 151620 -166815
rect 151712 -166859 151720 -166815
rect 151812 -166859 151820 -166815
rect 151912 -166859 151920 -166815
rect 152012 -166859 152020 -166815
rect 152112 -166859 152120 -166815
rect 152212 -166859 152220 -166815
rect 152312 -166859 152320 -166815
rect 152412 -166859 152420 -166815
rect 152512 -166859 152520 -166815
rect 152612 -166859 152620 -166815
rect 152712 -166859 152720 -166815
rect 152812 -166859 152820 -166815
rect 145268 -166915 145312 -166907
rect 145368 -166915 145412 -166907
rect 145468 -166915 145512 -166907
rect 145568 -166915 145612 -166907
rect 145668 -166915 145712 -166907
rect 145768 -166915 145812 -166907
rect 145868 -166915 145912 -166907
rect 145968 -166915 146012 -166907
rect 146068 -166915 146112 -166907
rect 146168 -166915 146212 -166907
rect 146268 -166915 146312 -166907
rect 146368 -166915 146412 -166907
rect 146468 -166915 146512 -166907
rect 146568 -166915 146612 -166907
rect 146668 -166915 146712 -166907
rect 146768 -166915 146812 -166907
rect 147268 -166915 147312 -166907
rect 147368 -166915 147412 -166907
rect 147468 -166915 147512 -166907
rect 147568 -166915 147612 -166907
rect 147668 -166915 147712 -166907
rect 147768 -166915 147812 -166907
rect 147868 -166915 147912 -166907
rect 147968 -166915 148012 -166907
rect 148068 -166915 148112 -166907
rect 148168 -166915 148212 -166907
rect 148268 -166915 148312 -166907
rect 148368 -166915 148412 -166907
rect 148468 -166915 148512 -166907
rect 148568 -166915 148612 -166907
rect 148668 -166915 148712 -166907
rect 148768 -166915 148812 -166907
rect 149268 -166915 149312 -166907
rect 149368 -166915 149412 -166907
rect 149468 -166915 149512 -166907
rect 149568 -166915 149612 -166907
rect 149668 -166915 149712 -166907
rect 149768 -166915 149812 -166907
rect 149868 -166915 149912 -166907
rect 149968 -166915 150012 -166907
rect 150068 -166915 150112 -166907
rect 150168 -166915 150212 -166907
rect 150268 -166915 150312 -166907
rect 150368 -166915 150412 -166907
rect 150468 -166915 150512 -166907
rect 150568 -166915 150612 -166907
rect 150668 -166915 150712 -166907
rect 150768 -166915 150812 -166907
rect 151268 -166915 151312 -166907
rect 151368 -166915 151412 -166907
rect 151468 -166915 151512 -166907
rect 151568 -166915 151612 -166907
rect 151668 -166915 151712 -166907
rect 151768 -166915 151812 -166907
rect 151868 -166915 151912 -166907
rect 151968 -166915 152012 -166907
rect 152068 -166915 152112 -166907
rect 152168 -166915 152212 -166907
rect 152268 -166915 152312 -166907
rect 152368 -166915 152412 -166907
rect 152468 -166915 152512 -166907
rect 152568 -166915 152612 -166907
rect 152668 -166915 152712 -166907
rect 152768 -166915 152812 -166907
rect 145312 -166959 145320 -166915
rect 145412 -166959 145420 -166915
rect 145512 -166959 145520 -166915
rect 145612 -166959 145620 -166915
rect 145712 -166959 145720 -166915
rect 145812 -166959 145820 -166915
rect 145912 -166959 145920 -166915
rect 146012 -166959 146020 -166915
rect 146112 -166959 146120 -166915
rect 146212 -166959 146220 -166915
rect 146312 -166959 146320 -166915
rect 146412 -166959 146420 -166915
rect 146512 -166959 146520 -166915
rect 146612 -166959 146620 -166915
rect 146712 -166959 146720 -166915
rect 146812 -166959 146820 -166915
rect 147312 -166959 147320 -166915
rect 147412 -166959 147420 -166915
rect 147512 -166959 147520 -166915
rect 147612 -166959 147620 -166915
rect 147712 -166959 147720 -166915
rect 147812 -166959 147820 -166915
rect 147912 -166959 147920 -166915
rect 148012 -166959 148020 -166915
rect 148112 -166959 148120 -166915
rect 148212 -166959 148220 -166915
rect 148312 -166959 148320 -166915
rect 148412 -166959 148420 -166915
rect 148512 -166959 148520 -166915
rect 148612 -166959 148620 -166915
rect 148712 -166959 148720 -166915
rect 148812 -166959 148820 -166915
rect 149312 -166959 149320 -166915
rect 149412 -166959 149420 -166915
rect 149512 -166959 149520 -166915
rect 149612 -166959 149620 -166915
rect 149712 -166959 149720 -166915
rect 149812 -166959 149820 -166915
rect 149912 -166959 149920 -166915
rect 150012 -166959 150020 -166915
rect 150112 -166959 150120 -166915
rect 150212 -166959 150220 -166915
rect 150312 -166959 150320 -166915
rect 150412 -166959 150420 -166915
rect 150512 -166959 150520 -166915
rect 150612 -166959 150620 -166915
rect 150712 -166959 150720 -166915
rect 150812 -166959 150820 -166915
rect 151312 -166959 151320 -166915
rect 151412 -166959 151420 -166915
rect 151512 -166959 151520 -166915
rect 151612 -166959 151620 -166915
rect 151712 -166959 151720 -166915
rect 151812 -166959 151820 -166915
rect 151912 -166959 151920 -166915
rect 152012 -166959 152020 -166915
rect 152112 -166959 152120 -166915
rect 152212 -166959 152220 -166915
rect 152312 -166959 152320 -166915
rect 152412 -166959 152420 -166915
rect 152512 -166959 152520 -166915
rect 152612 -166959 152620 -166915
rect 152712 -166959 152720 -166915
rect 152812 -166959 152820 -166915
rect 145268 -167015 145312 -167007
rect 145368 -167015 145412 -167007
rect 145468 -167015 145512 -167007
rect 145568 -167015 145612 -167007
rect 145668 -167015 145712 -167007
rect 145768 -167015 145812 -167007
rect 145868 -167015 145912 -167007
rect 145968 -167015 146012 -167007
rect 146068 -167015 146112 -167007
rect 146168 -167015 146212 -167007
rect 146268 -167015 146312 -167007
rect 146368 -167015 146412 -167007
rect 146468 -167015 146512 -167007
rect 146568 -167015 146612 -167007
rect 146668 -167015 146712 -167007
rect 146768 -167015 146812 -167007
rect 147268 -167015 147312 -167007
rect 147368 -167015 147412 -167007
rect 147468 -167015 147512 -167007
rect 147568 -167015 147612 -167007
rect 147668 -167015 147712 -167007
rect 147768 -167015 147812 -167007
rect 147868 -167015 147912 -167007
rect 147968 -167015 148012 -167007
rect 148068 -167015 148112 -167007
rect 148168 -167015 148212 -167007
rect 148268 -167015 148312 -167007
rect 148368 -167015 148412 -167007
rect 148468 -167015 148512 -167007
rect 148568 -167015 148612 -167007
rect 148668 -167015 148712 -167007
rect 148768 -167015 148812 -167007
rect 149268 -167015 149312 -167007
rect 149368 -167015 149412 -167007
rect 149468 -167015 149512 -167007
rect 149568 -167015 149612 -167007
rect 149668 -167015 149712 -167007
rect 149768 -167015 149812 -167007
rect 149868 -167015 149912 -167007
rect 149968 -167015 150012 -167007
rect 150068 -167015 150112 -167007
rect 150168 -167015 150212 -167007
rect 150268 -167015 150312 -167007
rect 150368 -167015 150412 -167007
rect 150468 -167015 150512 -167007
rect 150568 -167015 150612 -167007
rect 150668 -167015 150712 -167007
rect 150768 -167015 150812 -167007
rect 151268 -167015 151312 -167007
rect 151368 -167015 151412 -167007
rect 151468 -167015 151512 -167007
rect 151568 -167015 151612 -167007
rect 151668 -167015 151712 -167007
rect 151768 -167015 151812 -167007
rect 151868 -167015 151912 -167007
rect 151968 -167015 152012 -167007
rect 152068 -167015 152112 -167007
rect 152168 -167015 152212 -167007
rect 152268 -167015 152312 -167007
rect 152368 -167015 152412 -167007
rect 152468 -167015 152512 -167007
rect 152568 -167015 152612 -167007
rect 152668 -167015 152712 -167007
rect 152768 -167015 152812 -167007
rect 145312 -167059 145320 -167015
rect 145412 -167059 145420 -167015
rect 145512 -167059 145520 -167015
rect 145612 -167059 145620 -167015
rect 145712 -167059 145720 -167015
rect 145812 -167059 145820 -167015
rect 145912 -167059 145920 -167015
rect 146012 -167059 146020 -167015
rect 146112 -167059 146120 -167015
rect 146212 -167059 146220 -167015
rect 146312 -167059 146320 -167015
rect 146412 -167059 146420 -167015
rect 146512 -167059 146520 -167015
rect 146612 -167059 146620 -167015
rect 146712 -167059 146720 -167015
rect 146812 -167059 146820 -167015
rect 147312 -167059 147320 -167015
rect 147412 -167059 147420 -167015
rect 147512 -167059 147520 -167015
rect 147612 -167059 147620 -167015
rect 147712 -167059 147720 -167015
rect 147812 -167059 147820 -167015
rect 147912 -167059 147920 -167015
rect 148012 -167059 148020 -167015
rect 148112 -167059 148120 -167015
rect 148212 -167059 148220 -167015
rect 148312 -167059 148320 -167015
rect 148412 -167059 148420 -167015
rect 148512 -167059 148520 -167015
rect 148612 -167059 148620 -167015
rect 148712 -167059 148720 -167015
rect 148812 -167059 148820 -167015
rect 149312 -167059 149320 -167015
rect 149412 -167059 149420 -167015
rect 149512 -167059 149520 -167015
rect 149612 -167059 149620 -167015
rect 149712 -167059 149720 -167015
rect 149812 -167059 149820 -167015
rect 149912 -167059 149920 -167015
rect 150012 -167059 150020 -167015
rect 150112 -167059 150120 -167015
rect 150212 -167059 150220 -167015
rect 150312 -167059 150320 -167015
rect 150412 -167059 150420 -167015
rect 150512 -167059 150520 -167015
rect 150612 -167059 150620 -167015
rect 150712 -167059 150720 -167015
rect 150812 -167059 150820 -167015
rect 151312 -167059 151320 -167015
rect 151412 -167059 151420 -167015
rect 151512 -167059 151520 -167015
rect 151612 -167059 151620 -167015
rect 151712 -167059 151720 -167015
rect 151812 -167059 151820 -167015
rect 151912 -167059 151920 -167015
rect 152012 -167059 152020 -167015
rect 152112 -167059 152120 -167015
rect 152212 -167059 152220 -167015
rect 152312 -167059 152320 -167015
rect 152412 -167059 152420 -167015
rect 152512 -167059 152520 -167015
rect 152612 -167059 152620 -167015
rect 152712 -167059 152720 -167015
rect 152812 -167059 152820 -167015
rect 145268 -167115 145312 -167107
rect 145368 -167115 145412 -167107
rect 145468 -167115 145512 -167107
rect 145568 -167115 145612 -167107
rect 145668 -167115 145712 -167107
rect 145768 -167115 145812 -167107
rect 145868 -167115 145912 -167107
rect 145968 -167115 146012 -167107
rect 146068 -167115 146112 -167107
rect 146168 -167115 146212 -167107
rect 146268 -167115 146312 -167107
rect 146368 -167115 146412 -167107
rect 146468 -167115 146512 -167107
rect 146568 -167115 146612 -167107
rect 146668 -167115 146712 -167107
rect 146768 -167115 146812 -167107
rect 147268 -167115 147312 -167107
rect 147368 -167115 147412 -167107
rect 147468 -167115 147512 -167107
rect 147568 -167115 147612 -167107
rect 147668 -167115 147712 -167107
rect 147768 -167115 147812 -167107
rect 147868 -167115 147912 -167107
rect 147968 -167115 148012 -167107
rect 148068 -167115 148112 -167107
rect 148168 -167115 148212 -167107
rect 148268 -167115 148312 -167107
rect 148368 -167115 148412 -167107
rect 148468 -167115 148512 -167107
rect 148568 -167115 148612 -167107
rect 148668 -167115 148712 -167107
rect 148768 -167115 148812 -167107
rect 149268 -167115 149312 -167107
rect 149368 -167115 149412 -167107
rect 149468 -167115 149512 -167107
rect 149568 -167115 149612 -167107
rect 149668 -167115 149712 -167107
rect 149768 -167115 149812 -167107
rect 149868 -167115 149912 -167107
rect 149968 -167115 150012 -167107
rect 150068 -167115 150112 -167107
rect 150168 -167115 150212 -167107
rect 150268 -167115 150312 -167107
rect 150368 -167115 150412 -167107
rect 150468 -167115 150512 -167107
rect 150568 -167115 150612 -167107
rect 150668 -167115 150712 -167107
rect 150768 -167115 150812 -167107
rect 151268 -167115 151312 -167107
rect 151368 -167115 151412 -167107
rect 151468 -167115 151512 -167107
rect 151568 -167115 151612 -167107
rect 151668 -167115 151712 -167107
rect 151768 -167115 151812 -167107
rect 151868 -167115 151912 -167107
rect 151968 -167115 152012 -167107
rect 152068 -167115 152112 -167107
rect 152168 -167115 152212 -167107
rect 152268 -167115 152312 -167107
rect 152368 -167115 152412 -167107
rect 152468 -167115 152512 -167107
rect 152568 -167115 152612 -167107
rect 152668 -167115 152712 -167107
rect 152768 -167115 152812 -167107
rect 145312 -167159 145320 -167115
rect 145412 -167159 145420 -167115
rect 145512 -167159 145520 -167115
rect 145612 -167159 145620 -167115
rect 145712 -167159 145720 -167115
rect 145812 -167159 145820 -167115
rect 145912 -167159 145920 -167115
rect 146012 -167159 146020 -167115
rect 146112 -167159 146120 -167115
rect 146212 -167159 146220 -167115
rect 146312 -167159 146320 -167115
rect 146412 -167159 146420 -167115
rect 146512 -167159 146520 -167115
rect 146612 -167159 146620 -167115
rect 146712 -167159 146720 -167115
rect 146812 -167159 146820 -167115
rect 147312 -167159 147320 -167115
rect 147412 -167159 147420 -167115
rect 147512 -167159 147520 -167115
rect 147612 -167159 147620 -167115
rect 147712 -167159 147720 -167115
rect 147812 -167159 147820 -167115
rect 147912 -167159 147920 -167115
rect 148012 -167159 148020 -167115
rect 148112 -167159 148120 -167115
rect 148212 -167159 148220 -167115
rect 148312 -167159 148320 -167115
rect 148412 -167159 148420 -167115
rect 148512 -167159 148520 -167115
rect 148612 -167159 148620 -167115
rect 148712 -167159 148720 -167115
rect 148812 -167159 148820 -167115
rect 149312 -167159 149320 -167115
rect 149412 -167159 149420 -167115
rect 149512 -167159 149520 -167115
rect 149612 -167159 149620 -167115
rect 149712 -167159 149720 -167115
rect 149812 -167159 149820 -167115
rect 149912 -167159 149920 -167115
rect 150012 -167159 150020 -167115
rect 150112 -167159 150120 -167115
rect 150212 -167159 150220 -167115
rect 150312 -167159 150320 -167115
rect 150412 -167159 150420 -167115
rect 150512 -167159 150520 -167115
rect 150612 -167159 150620 -167115
rect 150712 -167159 150720 -167115
rect 150812 -167159 150820 -167115
rect 151312 -167159 151320 -167115
rect 151412 -167159 151420 -167115
rect 151512 -167159 151520 -167115
rect 151612 -167159 151620 -167115
rect 151712 -167159 151720 -167115
rect 151812 -167159 151820 -167115
rect 151912 -167159 151920 -167115
rect 152012 -167159 152020 -167115
rect 152112 -167159 152120 -167115
rect 152212 -167159 152220 -167115
rect 152312 -167159 152320 -167115
rect 152412 -167159 152420 -167115
rect 152512 -167159 152520 -167115
rect 152612 -167159 152620 -167115
rect 152712 -167159 152720 -167115
rect 152812 -167159 152820 -167115
rect 165525 -172989 165569 -172981
rect 165625 -172989 165669 -172981
rect 165725 -172989 165769 -172981
rect 165825 -172989 165869 -172981
rect 165925 -172989 165969 -172981
rect 166025 -172989 166069 -172981
rect 166125 -172989 166169 -172981
rect 166225 -172989 166269 -172981
rect 166325 -172989 166369 -172981
rect 166425 -172989 166469 -172981
rect 166525 -172989 166569 -172981
rect 166625 -172989 166669 -172981
rect 166725 -172989 166769 -172981
rect 166825 -172989 166869 -172981
rect 166925 -172989 166969 -172981
rect 167025 -172989 167069 -172981
rect 167525 -172989 167569 -172981
rect 167625 -172989 167669 -172981
rect 167725 -172989 167769 -172981
rect 167825 -172989 167869 -172981
rect 167925 -172989 167969 -172981
rect 168025 -172989 168069 -172981
rect 168125 -172989 168169 -172981
rect 168225 -172989 168269 -172981
rect 168325 -172989 168369 -172981
rect 168425 -172989 168469 -172981
rect 168525 -172989 168569 -172981
rect 168625 -172989 168669 -172981
rect 168725 -172989 168769 -172981
rect 168825 -172989 168869 -172981
rect 168925 -172989 168969 -172981
rect 169025 -172989 169069 -172981
rect 169525 -172989 169569 -172981
rect 169625 -172989 169669 -172981
rect 169725 -172989 169769 -172981
rect 169825 -172989 169869 -172981
rect 169925 -172989 169969 -172981
rect 170025 -172989 170069 -172981
rect 170125 -172989 170169 -172981
rect 170225 -172989 170269 -172981
rect 170325 -172989 170369 -172981
rect 170425 -172989 170469 -172981
rect 170525 -172989 170569 -172981
rect 170625 -172989 170669 -172981
rect 170725 -172989 170769 -172981
rect 170825 -172989 170869 -172981
rect 170925 -172989 170969 -172981
rect 171025 -172989 171069 -172981
rect 171525 -172989 171569 -172981
rect 171625 -172989 171669 -172981
rect 171725 -172989 171769 -172981
rect 171825 -172989 171869 -172981
rect 171925 -172989 171969 -172981
rect 172025 -172989 172069 -172981
rect 172125 -172989 172169 -172981
rect 172225 -172989 172269 -172981
rect 172325 -172989 172369 -172981
rect 172425 -172989 172469 -172981
rect 172525 -172989 172569 -172981
rect 172625 -172989 172669 -172981
rect 172725 -172989 172769 -172981
rect 172825 -172989 172869 -172981
rect 172925 -172989 172969 -172981
rect 173025 -172989 173069 -172981
rect 165569 -173033 165577 -172989
rect 165669 -173033 165677 -172989
rect 165769 -173033 165777 -172989
rect 165869 -173033 165877 -172989
rect 165969 -173033 165977 -172989
rect 166069 -173033 166077 -172989
rect 166169 -173033 166177 -172989
rect 166269 -173033 166277 -172989
rect 166369 -173033 166377 -172989
rect 166469 -173033 166477 -172989
rect 166569 -173033 166577 -172989
rect 166669 -173033 166677 -172989
rect 166769 -173033 166777 -172989
rect 166869 -173033 166877 -172989
rect 166969 -173033 166977 -172989
rect 167069 -173033 167077 -172989
rect 167569 -173033 167577 -172989
rect 167669 -173033 167677 -172989
rect 167769 -173033 167777 -172989
rect 167869 -173033 167877 -172989
rect 167969 -173033 167977 -172989
rect 168069 -173033 168077 -172989
rect 168169 -173033 168177 -172989
rect 168269 -173033 168277 -172989
rect 168369 -173033 168377 -172989
rect 168469 -173033 168477 -172989
rect 168569 -173033 168577 -172989
rect 168669 -173033 168677 -172989
rect 168769 -173033 168777 -172989
rect 168869 -173033 168877 -172989
rect 168969 -173033 168977 -172989
rect 169069 -173033 169077 -172989
rect 169569 -173033 169577 -172989
rect 169669 -173033 169677 -172989
rect 169769 -173033 169777 -172989
rect 169869 -173033 169877 -172989
rect 169969 -173033 169977 -172989
rect 170069 -173033 170077 -172989
rect 170169 -173033 170177 -172989
rect 170269 -173033 170277 -172989
rect 170369 -173033 170377 -172989
rect 170469 -173033 170477 -172989
rect 170569 -173033 170577 -172989
rect 170669 -173033 170677 -172989
rect 170769 -173033 170777 -172989
rect 170869 -173033 170877 -172989
rect 170969 -173033 170977 -172989
rect 171069 -173033 171077 -172989
rect 171569 -173033 171577 -172989
rect 171669 -173033 171677 -172989
rect 171769 -173033 171777 -172989
rect 171869 -173033 171877 -172989
rect 171969 -173033 171977 -172989
rect 172069 -173033 172077 -172989
rect 172169 -173033 172177 -172989
rect 172269 -173033 172277 -172989
rect 172369 -173033 172377 -172989
rect 172469 -173033 172477 -172989
rect 172569 -173033 172577 -172989
rect 172669 -173033 172677 -172989
rect 172769 -173033 172777 -172989
rect 172869 -173033 172877 -172989
rect 172969 -173033 172977 -172989
rect 173069 -173033 173077 -172989
rect 81627 -173049 81671 -173041
rect 81727 -173049 81771 -173041
rect 81827 -173049 81871 -173041
rect 81927 -173049 81971 -173041
rect 82027 -173049 82071 -173041
rect 82127 -173049 82171 -173041
rect 82227 -173049 82271 -173041
rect 82327 -173049 82371 -173041
rect 82427 -173049 82471 -173041
rect 82527 -173049 82571 -173041
rect 82627 -173049 82671 -173041
rect 82727 -173049 82771 -173041
rect 82827 -173049 82871 -173041
rect 82927 -173049 82971 -173041
rect 83027 -173049 83071 -173041
rect 83127 -173049 83171 -173041
rect 83627 -173049 83671 -173041
rect 83727 -173049 83771 -173041
rect 83827 -173049 83871 -173041
rect 83927 -173049 83971 -173041
rect 84027 -173049 84071 -173041
rect 84127 -173049 84171 -173041
rect 84227 -173049 84271 -173041
rect 84327 -173049 84371 -173041
rect 84427 -173049 84471 -173041
rect 84527 -173049 84571 -173041
rect 84627 -173049 84671 -173041
rect 84727 -173049 84771 -173041
rect 84827 -173049 84871 -173041
rect 84927 -173049 84971 -173041
rect 85027 -173049 85071 -173041
rect 85127 -173049 85171 -173041
rect 85627 -173049 85671 -173041
rect 85727 -173049 85771 -173041
rect 85827 -173049 85871 -173041
rect 85927 -173049 85971 -173041
rect 86027 -173049 86071 -173041
rect 86127 -173049 86171 -173041
rect 86227 -173049 86271 -173041
rect 86327 -173049 86371 -173041
rect 86427 -173049 86471 -173041
rect 86527 -173049 86571 -173041
rect 86627 -173049 86671 -173041
rect 86727 -173049 86771 -173041
rect 86827 -173049 86871 -173041
rect 86927 -173049 86971 -173041
rect 87027 -173049 87071 -173041
rect 87127 -173049 87171 -173041
rect 87627 -173049 87671 -173041
rect 87727 -173049 87771 -173041
rect 87827 -173049 87871 -173041
rect 87927 -173049 87971 -173041
rect 88027 -173049 88071 -173041
rect 88127 -173049 88171 -173041
rect 88227 -173049 88271 -173041
rect 88327 -173049 88371 -173041
rect 88427 -173049 88471 -173041
rect 88527 -173049 88571 -173041
rect 88627 -173049 88671 -173041
rect 88727 -173049 88771 -173041
rect 88827 -173049 88871 -173041
rect 88927 -173049 88971 -173041
rect 89027 -173049 89071 -173041
rect 89127 -173049 89171 -173041
rect 81671 -173093 81679 -173049
rect 81771 -173093 81779 -173049
rect 81871 -173093 81879 -173049
rect 81971 -173093 81979 -173049
rect 82071 -173093 82079 -173049
rect 82171 -173093 82179 -173049
rect 82271 -173093 82279 -173049
rect 82371 -173093 82379 -173049
rect 82471 -173093 82479 -173049
rect 82571 -173093 82579 -173049
rect 82671 -173093 82679 -173049
rect 82771 -173093 82779 -173049
rect 82871 -173093 82879 -173049
rect 82971 -173093 82979 -173049
rect 83071 -173093 83079 -173049
rect 83171 -173093 83179 -173049
rect 83671 -173093 83679 -173049
rect 83771 -173093 83779 -173049
rect 83871 -173093 83879 -173049
rect 83971 -173093 83979 -173049
rect 84071 -173093 84079 -173049
rect 84171 -173093 84179 -173049
rect 84271 -173093 84279 -173049
rect 84371 -173093 84379 -173049
rect 84471 -173093 84479 -173049
rect 84571 -173093 84579 -173049
rect 84671 -173093 84679 -173049
rect 84771 -173093 84779 -173049
rect 84871 -173093 84879 -173049
rect 84971 -173093 84979 -173049
rect 85071 -173093 85079 -173049
rect 85171 -173093 85179 -173049
rect 85671 -173093 85679 -173049
rect 85771 -173093 85779 -173049
rect 85871 -173093 85879 -173049
rect 85971 -173093 85979 -173049
rect 86071 -173093 86079 -173049
rect 86171 -173093 86179 -173049
rect 86271 -173093 86279 -173049
rect 86371 -173093 86379 -173049
rect 86471 -173093 86479 -173049
rect 86571 -173093 86579 -173049
rect 86671 -173093 86679 -173049
rect 86771 -173093 86779 -173049
rect 86871 -173093 86879 -173049
rect 86971 -173093 86979 -173049
rect 87071 -173093 87079 -173049
rect 87171 -173093 87179 -173049
rect 87671 -173093 87679 -173049
rect 87771 -173093 87779 -173049
rect 87871 -173093 87879 -173049
rect 87971 -173093 87979 -173049
rect 88071 -173093 88079 -173049
rect 88171 -173093 88179 -173049
rect 88271 -173093 88279 -173049
rect 88371 -173093 88379 -173049
rect 88471 -173093 88479 -173049
rect 88571 -173093 88579 -173049
rect 88671 -173093 88679 -173049
rect 88771 -173093 88779 -173049
rect 88871 -173093 88879 -173049
rect 88971 -173093 88979 -173049
rect 89071 -173093 89079 -173049
rect 89171 -173093 89179 -173049
rect 165525 -173089 165569 -173081
rect 165625 -173089 165669 -173081
rect 165725 -173089 165769 -173081
rect 165825 -173089 165869 -173081
rect 165925 -173089 165969 -173081
rect 166025 -173089 166069 -173081
rect 166125 -173089 166169 -173081
rect 166225 -173089 166269 -173081
rect 166325 -173089 166369 -173081
rect 166425 -173089 166469 -173081
rect 166525 -173089 166569 -173081
rect 166625 -173089 166669 -173081
rect 166725 -173089 166769 -173081
rect 166825 -173089 166869 -173081
rect 166925 -173089 166969 -173081
rect 167025 -173089 167069 -173081
rect 167525 -173089 167569 -173081
rect 167625 -173089 167669 -173081
rect 167725 -173089 167769 -173081
rect 167825 -173089 167869 -173081
rect 167925 -173089 167969 -173081
rect 168025 -173089 168069 -173081
rect 168125 -173089 168169 -173081
rect 168225 -173089 168269 -173081
rect 168325 -173089 168369 -173081
rect 168425 -173089 168469 -173081
rect 168525 -173089 168569 -173081
rect 168625 -173089 168669 -173081
rect 168725 -173089 168769 -173081
rect 168825 -173089 168869 -173081
rect 168925 -173089 168969 -173081
rect 169025 -173089 169069 -173081
rect 169525 -173089 169569 -173081
rect 169625 -173089 169669 -173081
rect 169725 -173089 169769 -173081
rect 169825 -173089 169869 -173081
rect 169925 -173089 169969 -173081
rect 170025 -173089 170069 -173081
rect 170125 -173089 170169 -173081
rect 170225 -173089 170269 -173081
rect 170325 -173089 170369 -173081
rect 170425 -173089 170469 -173081
rect 170525 -173089 170569 -173081
rect 170625 -173089 170669 -173081
rect 170725 -173089 170769 -173081
rect 170825 -173089 170869 -173081
rect 170925 -173089 170969 -173081
rect 171025 -173089 171069 -173081
rect 171525 -173089 171569 -173081
rect 171625 -173089 171669 -173081
rect 171725 -173089 171769 -173081
rect 171825 -173089 171869 -173081
rect 171925 -173089 171969 -173081
rect 172025 -173089 172069 -173081
rect 172125 -173089 172169 -173081
rect 172225 -173089 172269 -173081
rect 172325 -173089 172369 -173081
rect 172425 -173089 172469 -173081
rect 172525 -173089 172569 -173081
rect 172625 -173089 172669 -173081
rect 172725 -173089 172769 -173081
rect 172825 -173089 172869 -173081
rect 172925 -173089 172969 -173081
rect 173025 -173089 173069 -173081
rect 165569 -173133 165577 -173089
rect 165669 -173133 165677 -173089
rect 165769 -173133 165777 -173089
rect 165869 -173133 165877 -173089
rect 165969 -173133 165977 -173089
rect 166069 -173133 166077 -173089
rect 166169 -173133 166177 -173089
rect 166269 -173133 166277 -173089
rect 166369 -173133 166377 -173089
rect 166469 -173133 166477 -173089
rect 166569 -173133 166577 -173089
rect 166669 -173133 166677 -173089
rect 166769 -173133 166777 -173089
rect 166869 -173133 166877 -173089
rect 166969 -173133 166977 -173089
rect 167069 -173133 167077 -173089
rect 167569 -173133 167577 -173089
rect 167669 -173133 167677 -173089
rect 167769 -173133 167777 -173089
rect 167869 -173133 167877 -173089
rect 167969 -173133 167977 -173089
rect 168069 -173133 168077 -173089
rect 168169 -173133 168177 -173089
rect 168269 -173133 168277 -173089
rect 168369 -173133 168377 -173089
rect 168469 -173133 168477 -173089
rect 168569 -173133 168577 -173089
rect 168669 -173133 168677 -173089
rect 168769 -173133 168777 -173089
rect 168869 -173133 168877 -173089
rect 168969 -173133 168977 -173089
rect 169069 -173133 169077 -173089
rect 169569 -173133 169577 -173089
rect 169669 -173133 169677 -173089
rect 169769 -173133 169777 -173089
rect 169869 -173133 169877 -173089
rect 169969 -173133 169977 -173089
rect 170069 -173133 170077 -173089
rect 170169 -173133 170177 -173089
rect 170269 -173133 170277 -173089
rect 170369 -173133 170377 -173089
rect 170469 -173133 170477 -173089
rect 170569 -173133 170577 -173089
rect 170669 -173133 170677 -173089
rect 170769 -173133 170777 -173089
rect 170869 -173133 170877 -173089
rect 170969 -173133 170977 -173089
rect 171069 -173133 171077 -173089
rect 171569 -173133 171577 -173089
rect 171669 -173133 171677 -173089
rect 171769 -173133 171777 -173089
rect 171869 -173133 171877 -173089
rect 171969 -173133 171977 -173089
rect 172069 -173133 172077 -173089
rect 172169 -173133 172177 -173089
rect 172269 -173133 172277 -173089
rect 172369 -173133 172377 -173089
rect 172469 -173133 172477 -173089
rect 172569 -173133 172577 -173089
rect 172669 -173133 172677 -173089
rect 172769 -173133 172777 -173089
rect 172869 -173133 172877 -173089
rect 172969 -173133 172977 -173089
rect 173069 -173133 173077 -173089
rect 81627 -173149 81671 -173141
rect 81727 -173149 81771 -173141
rect 81827 -173149 81871 -173141
rect 81927 -173149 81971 -173141
rect 82027 -173149 82071 -173141
rect 82127 -173149 82171 -173141
rect 82227 -173149 82271 -173141
rect 82327 -173149 82371 -173141
rect 82427 -173149 82471 -173141
rect 82527 -173149 82571 -173141
rect 82627 -173149 82671 -173141
rect 82727 -173149 82771 -173141
rect 82827 -173149 82871 -173141
rect 82927 -173149 82971 -173141
rect 83027 -173149 83071 -173141
rect 83127 -173149 83171 -173141
rect 83627 -173149 83671 -173141
rect 83727 -173149 83771 -173141
rect 83827 -173149 83871 -173141
rect 83927 -173149 83971 -173141
rect 84027 -173149 84071 -173141
rect 84127 -173149 84171 -173141
rect 84227 -173149 84271 -173141
rect 84327 -173149 84371 -173141
rect 84427 -173149 84471 -173141
rect 84527 -173149 84571 -173141
rect 84627 -173149 84671 -173141
rect 84727 -173149 84771 -173141
rect 84827 -173149 84871 -173141
rect 84927 -173149 84971 -173141
rect 85027 -173149 85071 -173141
rect 85127 -173149 85171 -173141
rect 85627 -173149 85671 -173141
rect 85727 -173149 85771 -173141
rect 85827 -173149 85871 -173141
rect 85927 -173149 85971 -173141
rect 86027 -173149 86071 -173141
rect 86127 -173149 86171 -173141
rect 86227 -173149 86271 -173141
rect 86327 -173149 86371 -173141
rect 86427 -173149 86471 -173141
rect 86527 -173149 86571 -173141
rect 86627 -173149 86671 -173141
rect 86727 -173149 86771 -173141
rect 86827 -173149 86871 -173141
rect 86927 -173149 86971 -173141
rect 87027 -173149 87071 -173141
rect 87127 -173149 87171 -173141
rect 87627 -173149 87671 -173141
rect 87727 -173149 87771 -173141
rect 87827 -173149 87871 -173141
rect 87927 -173149 87971 -173141
rect 88027 -173149 88071 -173141
rect 88127 -173149 88171 -173141
rect 88227 -173149 88271 -173141
rect 88327 -173149 88371 -173141
rect 88427 -173149 88471 -173141
rect 88527 -173149 88571 -173141
rect 88627 -173149 88671 -173141
rect 88727 -173149 88771 -173141
rect 88827 -173149 88871 -173141
rect 88927 -173149 88971 -173141
rect 89027 -173149 89071 -173141
rect 89127 -173149 89171 -173141
rect 81671 -173193 81679 -173149
rect 81771 -173193 81779 -173149
rect 81871 -173193 81879 -173149
rect 81971 -173193 81979 -173149
rect 82071 -173193 82079 -173149
rect 82171 -173193 82179 -173149
rect 82271 -173193 82279 -173149
rect 82371 -173193 82379 -173149
rect 82471 -173193 82479 -173149
rect 82571 -173193 82579 -173149
rect 82671 -173193 82679 -173149
rect 82771 -173193 82779 -173149
rect 82871 -173193 82879 -173149
rect 82971 -173193 82979 -173149
rect 83071 -173193 83079 -173149
rect 83171 -173193 83179 -173149
rect 83671 -173193 83679 -173149
rect 83771 -173193 83779 -173149
rect 83871 -173193 83879 -173149
rect 83971 -173193 83979 -173149
rect 84071 -173193 84079 -173149
rect 84171 -173193 84179 -173149
rect 84271 -173193 84279 -173149
rect 84371 -173193 84379 -173149
rect 84471 -173193 84479 -173149
rect 84571 -173193 84579 -173149
rect 84671 -173193 84679 -173149
rect 84771 -173193 84779 -173149
rect 84871 -173193 84879 -173149
rect 84971 -173193 84979 -173149
rect 85071 -173193 85079 -173149
rect 85171 -173193 85179 -173149
rect 85671 -173193 85679 -173149
rect 85771 -173193 85779 -173149
rect 85871 -173193 85879 -173149
rect 85971 -173193 85979 -173149
rect 86071 -173193 86079 -173149
rect 86171 -173193 86179 -173149
rect 86271 -173193 86279 -173149
rect 86371 -173193 86379 -173149
rect 86471 -173193 86479 -173149
rect 86571 -173193 86579 -173149
rect 86671 -173193 86679 -173149
rect 86771 -173193 86779 -173149
rect 86871 -173193 86879 -173149
rect 86971 -173193 86979 -173149
rect 87071 -173193 87079 -173149
rect 87171 -173193 87179 -173149
rect 87671 -173193 87679 -173149
rect 87771 -173193 87779 -173149
rect 87871 -173193 87879 -173149
rect 87971 -173193 87979 -173149
rect 88071 -173193 88079 -173149
rect 88171 -173193 88179 -173149
rect 88271 -173193 88279 -173149
rect 88371 -173193 88379 -173149
rect 88471 -173193 88479 -173149
rect 88571 -173193 88579 -173149
rect 88671 -173193 88679 -173149
rect 88771 -173193 88779 -173149
rect 88871 -173193 88879 -173149
rect 88971 -173193 88979 -173149
rect 89071 -173193 89079 -173149
rect 89171 -173193 89179 -173149
rect 165525 -173189 165569 -173181
rect 165625 -173189 165669 -173181
rect 165725 -173189 165769 -173181
rect 165825 -173189 165869 -173181
rect 165925 -173189 165969 -173181
rect 166025 -173189 166069 -173181
rect 166125 -173189 166169 -173181
rect 166225 -173189 166269 -173181
rect 166325 -173189 166369 -173181
rect 166425 -173189 166469 -173181
rect 166525 -173189 166569 -173181
rect 166625 -173189 166669 -173181
rect 166725 -173189 166769 -173181
rect 166825 -173189 166869 -173181
rect 166925 -173189 166969 -173181
rect 167025 -173189 167069 -173181
rect 167525 -173189 167569 -173181
rect 167625 -173189 167669 -173181
rect 167725 -173189 167769 -173181
rect 167825 -173189 167869 -173181
rect 167925 -173189 167969 -173181
rect 168025 -173189 168069 -173181
rect 168125 -173189 168169 -173181
rect 168225 -173189 168269 -173181
rect 168325 -173189 168369 -173181
rect 168425 -173189 168469 -173181
rect 168525 -173189 168569 -173181
rect 168625 -173189 168669 -173181
rect 168725 -173189 168769 -173181
rect 168825 -173189 168869 -173181
rect 168925 -173189 168969 -173181
rect 169025 -173189 169069 -173181
rect 169525 -173189 169569 -173181
rect 169625 -173189 169669 -173181
rect 169725 -173189 169769 -173181
rect 169825 -173189 169869 -173181
rect 169925 -173189 169969 -173181
rect 170025 -173189 170069 -173181
rect 170125 -173189 170169 -173181
rect 170225 -173189 170269 -173181
rect 170325 -173189 170369 -173181
rect 170425 -173189 170469 -173181
rect 170525 -173189 170569 -173181
rect 170625 -173189 170669 -173181
rect 170725 -173189 170769 -173181
rect 170825 -173189 170869 -173181
rect 170925 -173189 170969 -173181
rect 171025 -173189 171069 -173181
rect 171525 -173189 171569 -173181
rect 171625 -173189 171669 -173181
rect 171725 -173189 171769 -173181
rect 171825 -173189 171869 -173181
rect 171925 -173189 171969 -173181
rect 172025 -173189 172069 -173181
rect 172125 -173189 172169 -173181
rect 172225 -173189 172269 -173181
rect 172325 -173189 172369 -173181
rect 172425 -173189 172469 -173181
rect 172525 -173189 172569 -173181
rect 172625 -173189 172669 -173181
rect 172725 -173189 172769 -173181
rect 172825 -173189 172869 -173181
rect 172925 -173189 172969 -173181
rect 173025 -173189 173069 -173181
rect 165569 -173233 165577 -173189
rect 165669 -173233 165677 -173189
rect 165769 -173233 165777 -173189
rect 165869 -173233 165877 -173189
rect 165969 -173233 165977 -173189
rect 166069 -173233 166077 -173189
rect 166169 -173233 166177 -173189
rect 166269 -173233 166277 -173189
rect 166369 -173233 166377 -173189
rect 166469 -173233 166477 -173189
rect 166569 -173233 166577 -173189
rect 166669 -173233 166677 -173189
rect 166769 -173233 166777 -173189
rect 166869 -173233 166877 -173189
rect 166969 -173233 166977 -173189
rect 167069 -173233 167077 -173189
rect 167569 -173233 167577 -173189
rect 167669 -173233 167677 -173189
rect 167769 -173233 167777 -173189
rect 167869 -173233 167877 -173189
rect 167969 -173233 167977 -173189
rect 168069 -173233 168077 -173189
rect 168169 -173233 168177 -173189
rect 168269 -173233 168277 -173189
rect 168369 -173233 168377 -173189
rect 168469 -173233 168477 -173189
rect 168569 -173233 168577 -173189
rect 168669 -173233 168677 -173189
rect 168769 -173233 168777 -173189
rect 168869 -173233 168877 -173189
rect 168969 -173233 168977 -173189
rect 169069 -173233 169077 -173189
rect 169569 -173233 169577 -173189
rect 169669 -173233 169677 -173189
rect 169769 -173233 169777 -173189
rect 169869 -173233 169877 -173189
rect 169969 -173233 169977 -173189
rect 170069 -173233 170077 -173189
rect 170169 -173233 170177 -173189
rect 170269 -173233 170277 -173189
rect 170369 -173233 170377 -173189
rect 170469 -173233 170477 -173189
rect 170569 -173233 170577 -173189
rect 170669 -173233 170677 -173189
rect 170769 -173233 170777 -173189
rect 170869 -173233 170877 -173189
rect 170969 -173233 170977 -173189
rect 171069 -173233 171077 -173189
rect 171569 -173233 171577 -173189
rect 171669 -173233 171677 -173189
rect 171769 -173233 171777 -173189
rect 171869 -173233 171877 -173189
rect 171969 -173233 171977 -173189
rect 172069 -173233 172077 -173189
rect 172169 -173233 172177 -173189
rect 172269 -173233 172277 -173189
rect 172369 -173233 172377 -173189
rect 172469 -173233 172477 -173189
rect 172569 -173233 172577 -173189
rect 172669 -173233 172677 -173189
rect 172769 -173233 172777 -173189
rect 172869 -173233 172877 -173189
rect 172969 -173233 172977 -173189
rect 173069 -173233 173077 -173189
rect 81627 -173249 81671 -173241
rect 81727 -173249 81771 -173241
rect 81827 -173249 81871 -173241
rect 81927 -173249 81971 -173241
rect 82027 -173249 82071 -173241
rect 82127 -173249 82171 -173241
rect 82227 -173249 82271 -173241
rect 82327 -173249 82371 -173241
rect 82427 -173249 82471 -173241
rect 82527 -173249 82571 -173241
rect 82627 -173249 82671 -173241
rect 82727 -173249 82771 -173241
rect 82827 -173249 82871 -173241
rect 82927 -173249 82971 -173241
rect 83027 -173249 83071 -173241
rect 83127 -173249 83171 -173241
rect 83627 -173249 83671 -173241
rect 83727 -173249 83771 -173241
rect 83827 -173249 83871 -173241
rect 83927 -173249 83971 -173241
rect 84027 -173249 84071 -173241
rect 84127 -173249 84171 -173241
rect 84227 -173249 84271 -173241
rect 84327 -173249 84371 -173241
rect 84427 -173249 84471 -173241
rect 84527 -173249 84571 -173241
rect 84627 -173249 84671 -173241
rect 84727 -173249 84771 -173241
rect 84827 -173249 84871 -173241
rect 84927 -173249 84971 -173241
rect 85027 -173249 85071 -173241
rect 85127 -173249 85171 -173241
rect 85627 -173249 85671 -173241
rect 85727 -173249 85771 -173241
rect 85827 -173249 85871 -173241
rect 85927 -173249 85971 -173241
rect 86027 -173249 86071 -173241
rect 86127 -173249 86171 -173241
rect 86227 -173249 86271 -173241
rect 86327 -173249 86371 -173241
rect 86427 -173249 86471 -173241
rect 86527 -173249 86571 -173241
rect 86627 -173249 86671 -173241
rect 86727 -173249 86771 -173241
rect 86827 -173249 86871 -173241
rect 86927 -173249 86971 -173241
rect 87027 -173249 87071 -173241
rect 87127 -173249 87171 -173241
rect 87627 -173249 87671 -173241
rect 87727 -173249 87771 -173241
rect 87827 -173249 87871 -173241
rect 87927 -173249 87971 -173241
rect 88027 -173249 88071 -173241
rect 88127 -173249 88171 -173241
rect 88227 -173249 88271 -173241
rect 88327 -173249 88371 -173241
rect 88427 -173249 88471 -173241
rect 88527 -173249 88571 -173241
rect 88627 -173249 88671 -173241
rect 88727 -173249 88771 -173241
rect 88827 -173249 88871 -173241
rect 88927 -173249 88971 -173241
rect 89027 -173249 89071 -173241
rect 89127 -173249 89171 -173241
rect 81671 -173293 81679 -173249
rect 81771 -173293 81779 -173249
rect 81871 -173293 81879 -173249
rect 81971 -173293 81979 -173249
rect 82071 -173293 82079 -173249
rect 82171 -173293 82179 -173249
rect 82271 -173293 82279 -173249
rect 82371 -173293 82379 -173249
rect 82471 -173293 82479 -173249
rect 82571 -173293 82579 -173249
rect 82671 -173293 82679 -173249
rect 82771 -173293 82779 -173249
rect 82871 -173293 82879 -173249
rect 82971 -173293 82979 -173249
rect 83071 -173293 83079 -173249
rect 83171 -173293 83179 -173249
rect 83671 -173293 83679 -173249
rect 83771 -173293 83779 -173249
rect 83871 -173293 83879 -173249
rect 83971 -173293 83979 -173249
rect 84071 -173293 84079 -173249
rect 84171 -173293 84179 -173249
rect 84271 -173293 84279 -173249
rect 84371 -173293 84379 -173249
rect 84471 -173293 84479 -173249
rect 84571 -173293 84579 -173249
rect 84671 -173293 84679 -173249
rect 84771 -173293 84779 -173249
rect 84871 -173293 84879 -173249
rect 84971 -173293 84979 -173249
rect 85071 -173293 85079 -173249
rect 85171 -173293 85179 -173249
rect 85671 -173293 85679 -173249
rect 85771 -173293 85779 -173249
rect 85871 -173293 85879 -173249
rect 85971 -173293 85979 -173249
rect 86071 -173293 86079 -173249
rect 86171 -173293 86179 -173249
rect 86271 -173293 86279 -173249
rect 86371 -173293 86379 -173249
rect 86471 -173293 86479 -173249
rect 86571 -173293 86579 -173249
rect 86671 -173293 86679 -173249
rect 86771 -173293 86779 -173249
rect 86871 -173293 86879 -173249
rect 86971 -173293 86979 -173249
rect 87071 -173293 87079 -173249
rect 87171 -173293 87179 -173249
rect 87671 -173293 87679 -173249
rect 87771 -173293 87779 -173249
rect 87871 -173293 87879 -173249
rect 87971 -173293 87979 -173249
rect 88071 -173293 88079 -173249
rect 88171 -173293 88179 -173249
rect 88271 -173293 88279 -173249
rect 88371 -173293 88379 -173249
rect 88471 -173293 88479 -173249
rect 88571 -173293 88579 -173249
rect 88671 -173293 88679 -173249
rect 88771 -173293 88779 -173249
rect 88871 -173293 88879 -173249
rect 88971 -173293 88979 -173249
rect 89071 -173293 89079 -173249
rect 89171 -173293 89179 -173249
rect 165525 -173289 165569 -173281
rect 165625 -173289 165669 -173281
rect 165725 -173289 165769 -173281
rect 165825 -173289 165869 -173281
rect 165925 -173289 165969 -173281
rect 166025 -173289 166069 -173281
rect 166125 -173289 166169 -173281
rect 166225 -173289 166269 -173281
rect 166325 -173289 166369 -173281
rect 166425 -173289 166469 -173281
rect 166525 -173289 166569 -173281
rect 166625 -173289 166669 -173281
rect 166725 -173289 166769 -173281
rect 166825 -173289 166869 -173281
rect 166925 -173289 166969 -173281
rect 167025 -173289 167069 -173281
rect 167525 -173289 167569 -173281
rect 167625 -173289 167669 -173281
rect 167725 -173289 167769 -173281
rect 167825 -173289 167869 -173281
rect 167925 -173289 167969 -173281
rect 168025 -173289 168069 -173281
rect 168125 -173289 168169 -173281
rect 168225 -173289 168269 -173281
rect 168325 -173289 168369 -173281
rect 168425 -173289 168469 -173281
rect 168525 -173289 168569 -173281
rect 168625 -173289 168669 -173281
rect 168725 -173289 168769 -173281
rect 168825 -173289 168869 -173281
rect 168925 -173289 168969 -173281
rect 169025 -173289 169069 -173281
rect 169525 -173289 169569 -173281
rect 169625 -173289 169669 -173281
rect 169725 -173289 169769 -173281
rect 169825 -173289 169869 -173281
rect 169925 -173289 169969 -173281
rect 170025 -173289 170069 -173281
rect 170125 -173289 170169 -173281
rect 170225 -173289 170269 -173281
rect 170325 -173289 170369 -173281
rect 170425 -173289 170469 -173281
rect 170525 -173289 170569 -173281
rect 170625 -173289 170669 -173281
rect 170725 -173289 170769 -173281
rect 170825 -173289 170869 -173281
rect 170925 -173289 170969 -173281
rect 171025 -173289 171069 -173281
rect 171525 -173289 171569 -173281
rect 171625 -173289 171669 -173281
rect 171725 -173289 171769 -173281
rect 171825 -173289 171869 -173281
rect 171925 -173289 171969 -173281
rect 172025 -173289 172069 -173281
rect 172125 -173289 172169 -173281
rect 172225 -173289 172269 -173281
rect 172325 -173289 172369 -173281
rect 172425 -173289 172469 -173281
rect 172525 -173289 172569 -173281
rect 172625 -173289 172669 -173281
rect 172725 -173289 172769 -173281
rect 172825 -173289 172869 -173281
rect 172925 -173289 172969 -173281
rect 173025 -173289 173069 -173281
rect 165569 -173333 165577 -173289
rect 165669 -173333 165677 -173289
rect 165769 -173333 165777 -173289
rect 165869 -173333 165877 -173289
rect 165969 -173333 165977 -173289
rect 166069 -173333 166077 -173289
rect 166169 -173333 166177 -173289
rect 166269 -173333 166277 -173289
rect 166369 -173333 166377 -173289
rect 166469 -173333 166477 -173289
rect 166569 -173333 166577 -173289
rect 166669 -173333 166677 -173289
rect 166769 -173333 166777 -173289
rect 166869 -173333 166877 -173289
rect 166969 -173333 166977 -173289
rect 167069 -173333 167077 -173289
rect 167569 -173333 167577 -173289
rect 167669 -173333 167677 -173289
rect 167769 -173333 167777 -173289
rect 167869 -173333 167877 -173289
rect 167969 -173333 167977 -173289
rect 168069 -173333 168077 -173289
rect 168169 -173333 168177 -173289
rect 168269 -173333 168277 -173289
rect 168369 -173333 168377 -173289
rect 168469 -173333 168477 -173289
rect 168569 -173333 168577 -173289
rect 168669 -173333 168677 -173289
rect 168769 -173333 168777 -173289
rect 168869 -173333 168877 -173289
rect 168969 -173333 168977 -173289
rect 169069 -173333 169077 -173289
rect 169569 -173333 169577 -173289
rect 169669 -173333 169677 -173289
rect 169769 -173333 169777 -173289
rect 169869 -173333 169877 -173289
rect 169969 -173333 169977 -173289
rect 170069 -173333 170077 -173289
rect 170169 -173333 170177 -173289
rect 170269 -173333 170277 -173289
rect 170369 -173333 170377 -173289
rect 170469 -173333 170477 -173289
rect 170569 -173333 170577 -173289
rect 170669 -173333 170677 -173289
rect 170769 -173333 170777 -173289
rect 170869 -173333 170877 -173289
rect 170969 -173333 170977 -173289
rect 171069 -173333 171077 -173289
rect 171569 -173333 171577 -173289
rect 171669 -173333 171677 -173289
rect 171769 -173333 171777 -173289
rect 171869 -173333 171877 -173289
rect 171969 -173333 171977 -173289
rect 172069 -173333 172077 -173289
rect 172169 -173333 172177 -173289
rect 172269 -173333 172277 -173289
rect 172369 -173333 172377 -173289
rect 172469 -173333 172477 -173289
rect 172569 -173333 172577 -173289
rect 172669 -173333 172677 -173289
rect 172769 -173333 172777 -173289
rect 172869 -173333 172877 -173289
rect 172969 -173333 172977 -173289
rect 173069 -173333 173077 -173289
rect 81627 -173349 81671 -173341
rect 81727 -173349 81771 -173341
rect 81827 -173349 81871 -173341
rect 81927 -173349 81971 -173341
rect 82027 -173349 82071 -173341
rect 82127 -173349 82171 -173341
rect 82227 -173349 82271 -173341
rect 82327 -173349 82371 -173341
rect 82427 -173349 82471 -173341
rect 82527 -173349 82571 -173341
rect 82627 -173349 82671 -173341
rect 82727 -173349 82771 -173341
rect 82827 -173349 82871 -173341
rect 82927 -173349 82971 -173341
rect 83027 -173349 83071 -173341
rect 83127 -173349 83171 -173341
rect 83627 -173349 83671 -173341
rect 83727 -173349 83771 -173341
rect 83827 -173349 83871 -173341
rect 83927 -173349 83971 -173341
rect 84027 -173349 84071 -173341
rect 84127 -173349 84171 -173341
rect 84227 -173349 84271 -173341
rect 84327 -173349 84371 -173341
rect 84427 -173349 84471 -173341
rect 84527 -173349 84571 -173341
rect 84627 -173349 84671 -173341
rect 84727 -173349 84771 -173341
rect 84827 -173349 84871 -173341
rect 84927 -173349 84971 -173341
rect 85027 -173349 85071 -173341
rect 85127 -173349 85171 -173341
rect 85627 -173349 85671 -173341
rect 85727 -173349 85771 -173341
rect 85827 -173349 85871 -173341
rect 85927 -173349 85971 -173341
rect 86027 -173349 86071 -173341
rect 86127 -173349 86171 -173341
rect 86227 -173349 86271 -173341
rect 86327 -173349 86371 -173341
rect 86427 -173349 86471 -173341
rect 86527 -173349 86571 -173341
rect 86627 -173349 86671 -173341
rect 86727 -173349 86771 -173341
rect 86827 -173349 86871 -173341
rect 86927 -173349 86971 -173341
rect 87027 -173349 87071 -173341
rect 87127 -173349 87171 -173341
rect 87627 -173349 87671 -173341
rect 87727 -173349 87771 -173341
rect 87827 -173349 87871 -173341
rect 87927 -173349 87971 -173341
rect 88027 -173349 88071 -173341
rect 88127 -173349 88171 -173341
rect 88227 -173349 88271 -173341
rect 88327 -173349 88371 -173341
rect 88427 -173349 88471 -173341
rect 88527 -173349 88571 -173341
rect 88627 -173349 88671 -173341
rect 88727 -173349 88771 -173341
rect 88827 -173349 88871 -173341
rect 88927 -173349 88971 -173341
rect 89027 -173349 89071 -173341
rect 89127 -173349 89171 -173341
rect 81671 -173393 81679 -173349
rect 81771 -173393 81779 -173349
rect 81871 -173393 81879 -173349
rect 81971 -173393 81979 -173349
rect 82071 -173393 82079 -173349
rect 82171 -173393 82179 -173349
rect 82271 -173393 82279 -173349
rect 82371 -173393 82379 -173349
rect 82471 -173393 82479 -173349
rect 82571 -173393 82579 -173349
rect 82671 -173393 82679 -173349
rect 82771 -173393 82779 -173349
rect 82871 -173393 82879 -173349
rect 82971 -173393 82979 -173349
rect 83071 -173393 83079 -173349
rect 83171 -173393 83179 -173349
rect 83671 -173393 83679 -173349
rect 83771 -173393 83779 -173349
rect 83871 -173393 83879 -173349
rect 83971 -173393 83979 -173349
rect 84071 -173393 84079 -173349
rect 84171 -173393 84179 -173349
rect 84271 -173393 84279 -173349
rect 84371 -173393 84379 -173349
rect 84471 -173393 84479 -173349
rect 84571 -173393 84579 -173349
rect 84671 -173393 84679 -173349
rect 84771 -173393 84779 -173349
rect 84871 -173393 84879 -173349
rect 84971 -173393 84979 -173349
rect 85071 -173393 85079 -173349
rect 85171 -173393 85179 -173349
rect 85671 -173393 85679 -173349
rect 85771 -173393 85779 -173349
rect 85871 -173393 85879 -173349
rect 85971 -173393 85979 -173349
rect 86071 -173393 86079 -173349
rect 86171 -173393 86179 -173349
rect 86271 -173393 86279 -173349
rect 86371 -173393 86379 -173349
rect 86471 -173393 86479 -173349
rect 86571 -173393 86579 -173349
rect 86671 -173393 86679 -173349
rect 86771 -173393 86779 -173349
rect 86871 -173393 86879 -173349
rect 86971 -173393 86979 -173349
rect 87071 -173393 87079 -173349
rect 87171 -173393 87179 -173349
rect 87671 -173393 87679 -173349
rect 87771 -173393 87779 -173349
rect 87871 -173393 87879 -173349
rect 87971 -173393 87979 -173349
rect 88071 -173393 88079 -173349
rect 88171 -173393 88179 -173349
rect 88271 -173393 88279 -173349
rect 88371 -173393 88379 -173349
rect 88471 -173393 88479 -173349
rect 88571 -173393 88579 -173349
rect 88671 -173393 88679 -173349
rect 88771 -173393 88779 -173349
rect 88871 -173393 88879 -173349
rect 88971 -173393 88979 -173349
rect 89071 -173393 89079 -173349
rect 89171 -173393 89179 -173349
rect 165525 -173389 165569 -173381
rect 165625 -173389 165669 -173381
rect 165725 -173389 165769 -173381
rect 165825 -173389 165869 -173381
rect 165925 -173389 165969 -173381
rect 166025 -173389 166069 -173381
rect 166125 -173389 166169 -173381
rect 166225 -173389 166269 -173381
rect 166325 -173389 166369 -173381
rect 166425 -173389 166469 -173381
rect 166525 -173389 166569 -173381
rect 166625 -173389 166669 -173381
rect 166725 -173389 166769 -173381
rect 166825 -173389 166869 -173381
rect 166925 -173389 166969 -173381
rect 167025 -173389 167069 -173381
rect 167525 -173389 167569 -173381
rect 167625 -173389 167669 -173381
rect 167725 -173389 167769 -173381
rect 167825 -173389 167869 -173381
rect 167925 -173389 167969 -173381
rect 168025 -173389 168069 -173381
rect 168125 -173389 168169 -173381
rect 168225 -173389 168269 -173381
rect 168325 -173389 168369 -173381
rect 168425 -173389 168469 -173381
rect 168525 -173389 168569 -173381
rect 168625 -173389 168669 -173381
rect 168725 -173389 168769 -173381
rect 168825 -173389 168869 -173381
rect 168925 -173389 168969 -173381
rect 169025 -173389 169069 -173381
rect 169525 -173389 169569 -173381
rect 169625 -173389 169669 -173381
rect 169725 -173389 169769 -173381
rect 169825 -173389 169869 -173381
rect 169925 -173389 169969 -173381
rect 170025 -173389 170069 -173381
rect 170125 -173389 170169 -173381
rect 170225 -173389 170269 -173381
rect 170325 -173389 170369 -173381
rect 170425 -173389 170469 -173381
rect 170525 -173389 170569 -173381
rect 170625 -173389 170669 -173381
rect 170725 -173389 170769 -173381
rect 170825 -173389 170869 -173381
rect 170925 -173389 170969 -173381
rect 171025 -173389 171069 -173381
rect 171525 -173389 171569 -173381
rect 171625 -173389 171669 -173381
rect 171725 -173389 171769 -173381
rect 171825 -173389 171869 -173381
rect 171925 -173389 171969 -173381
rect 172025 -173389 172069 -173381
rect 172125 -173389 172169 -173381
rect 172225 -173389 172269 -173381
rect 172325 -173389 172369 -173381
rect 172425 -173389 172469 -173381
rect 172525 -173389 172569 -173381
rect 172625 -173389 172669 -173381
rect 172725 -173389 172769 -173381
rect 172825 -173389 172869 -173381
rect 172925 -173389 172969 -173381
rect 173025 -173389 173069 -173381
rect 165569 -173433 165577 -173389
rect 165669 -173433 165677 -173389
rect 165769 -173433 165777 -173389
rect 165869 -173433 165877 -173389
rect 165969 -173433 165977 -173389
rect 166069 -173433 166077 -173389
rect 166169 -173433 166177 -173389
rect 166269 -173433 166277 -173389
rect 166369 -173433 166377 -173389
rect 166469 -173433 166477 -173389
rect 166569 -173433 166577 -173389
rect 166669 -173433 166677 -173389
rect 166769 -173433 166777 -173389
rect 166869 -173433 166877 -173389
rect 166969 -173433 166977 -173389
rect 167069 -173433 167077 -173389
rect 167569 -173433 167577 -173389
rect 167669 -173433 167677 -173389
rect 167769 -173433 167777 -173389
rect 167869 -173433 167877 -173389
rect 167969 -173433 167977 -173389
rect 168069 -173433 168077 -173389
rect 168169 -173433 168177 -173389
rect 168269 -173433 168277 -173389
rect 168369 -173433 168377 -173389
rect 168469 -173433 168477 -173389
rect 168569 -173433 168577 -173389
rect 168669 -173433 168677 -173389
rect 168769 -173433 168777 -173389
rect 168869 -173433 168877 -173389
rect 168969 -173433 168977 -173389
rect 169069 -173433 169077 -173389
rect 169569 -173433 169577 -173389
rect 169669 -173433 169677 -173389
rect 169769 -173433 169777 -173389
rect 169869 -173433 169877 -173389
rect 169969 -173433 169977 -173389
rect 170069 -173433 170077 -173389
rect 170169 -173433 170177 -173389
rect 170269 -173433 170277 -173389
rect 170369 -173433 170377 -173389
rect 170469 -173433 170477 -173389
rect 170569 -173433 170577 -173389
rect 170669 -173433 170677 -173389
rect 170769 -173433 170777 -173389
rect 170869 -173433 170877 -173389
rect 170969 -173433 170977 -173389
rect 171069 -173433 171077 -173389
rect 171569 -173433 171577 -173389
rect 171669 -173433 171677 -173389
rect 171769 -173433 171777 -173389
rect 171869 -173433 171877 -173389
rect 171969 -173433 171977 -173389
rect 172069 -173433 172077 -173389
rect 172169 -173433 172177 -173389
rect 172269 -173433 172277 -173389
rect 172369 -173433 172377 -173389
rect 172469 -173433 172477 -173389
rect 172569 -173433 172577 -173389
rect 172669 -173433 172677 -173389
rect 172769 -173433 172777 -173389
rect 172869 -173433 172877 -173389
rect 172969 -173433 172977 -173389
rect 173069 -173433 173077 -173389
rect 81627 -173449 81671 -173441
rect 81727 -173449 81771 -173441
rect 81827 -173449 81871 -173441
rect 81927 -173449 81971 -173441
rect 82027 -173449 82071 -173441
rect 82127 -173449 82171 -173441
rect 82227 -173449 82271 -173441
rect 82327 -173449 82371 -173441
rect 82427 -173449 82471 -173441
rect 82527 -173449 82571 -173441
rect 82627 -173449 82671 -173441
rect 82727 -173449 82771 -173441
rect 82827 -173449 82871 -173441
rect 82927 -173449 82971 -173441
rect 83027 -173449 83071 -173441
rect 83127 -173449 83171 -173441
rect 83627 -173449 83671 -173441
rect 83727 -173449 83771 -173441
rect 83827 -173449 83871 -173441
rect 83927 -173449 83971 -173441
rect 84027 -173449 84071 -173441
rect 84127 -173449 84171 -173441
rect 84227 -173449 84271 -173441
rect 84327 -173449 84371 -173441
rect 84427 -173449 84471 -173441
rect 84527 -173449 84571 -173441
rect 84627 -173449 84671 -173441
rect 84727 -173449 84771 -173441
rect 84827 -173449 84871 -173441
rect 84927 -173449 84971 -173441
rect 85027 -173449 85071 -173441
rect 85127 -173449 85171 -173441
rect 85627 -173449 85671 -173441
rect 85727 -173449 85771 -173441
rect 85827 -173449 85871 -173441
rect 85927 -173449 85971 -173441
rect 86027 -173449 86071 -173441
rect 86127 -173449 86171 -173441
rect 86227 -173449 86271 -173441
rect 86327 -173449 86371 -173441
rect 86427 -173449 86471 -173441
rect 86527 -173449 86571 -173441
rect 86627 -173449 86671 -173441
rect 86727 -173449 86771 -173441
rect 86827 -173449 86871 -173441
rect 86927 -173449 86971 -173441
rect 87027 -173449 87071 -173441
rect 87127 -173449 87171 -173441
rect 87627 -173449 87671 -173441
rect 87727 -173449 87771 -173441
rect 87827 -173449 87871 -173441
rect 87927 -173449 87971 -173441
rect 88027 -173449 88071 -173441
rect 88127 -173449 88171 -173441
rect 88227 -173449 88271 -173441
rect 88327 -173449 88371 -173441
rect 88427 -173449 88471 -173441
rect 88527 -173449 88571 -173441
rect 88627 -173449 88671 -173441
rect 88727 -173449 88771 -173441
rect 88827 -173449 88871 -173441
rect 88927 -173449 88971 -173441
rect 89027 -173449 89071 -173441
rect 89127 -173449 89171 -173441
rect 81671 -173493 81679 -173449
rect 81771 -173493 81779 -173449
rect 81871 -173493 81879 -173449
rect 81971 -173493 81979 -173449
rect 82071 -173493 82079 -173449
rect 82171 -173493 82179 -173449
rect 82271 -173493 82279 -173449
rect 82371 -173493 82379 -173449
rect 82471 -173493 82479 -173449
rect 82571 -173493 82579 -173449
rect 82671 -173493 82679 -173449
rect 82771 -173493 82779 -173449
rect 82871 -173493 82879 -173449
rect 82971 -173493 82979 -173449
rect 83071 -173493 83079 -173449
rect 83171 -173493 83179 -173449
rect 83671 -173493 83679 -173449
rect 83771 -173493 83779 -173449
rect 83871 -173493 83879 -173449
rect 83971 -173493 83979 -173449
rect 84071 -173493 84079 -173449
rect 84171 -173493 84179 -173449
rect 84271 -173493 84279 -173449
rect 84371 -173493 84379 -173449
rect 84471 -173493 84479 -173449
rect 84571 -173493 84579 -173449
rect 84671 -173493 84679 -173449
rect 84771 -173493 84779 -173449
rect 84871 -173493 84879 -173449
rect 84971 -173493 84979 -173449
rect 85071 -173493 85079 -173449
rect 85171 -173493 85179 -173449
rect 85671 -173493 85679 -173449
rect 85771 -173493 85779 -173449
rect 85871 -173493 85879 -173449
rect 85971 -173493 85979 -173449
rect 86071 -173493 86079 -173449
rect 86171 -173493 86179 -173449
rect 86271 -173493 86279 -173449
rect 86371 -173493 86379 -173449
rect 86471 -173493 86479 -173449
rect 86571 -173493 86579 -173449
rect 86671 -173493 86679 -173449
rect 86771 -173493 86779 -173449
rect 86871 -173493 86879 -173449
rect 86971 -173493 86979 -173449
rect 87071 -173493 87079 -173449
rect 87171 -173493 87179 -173449
rect 87671 -173493 87679 -173449
rect 87771 -173493 87779 -173449
rect 87871 -173493 87879 -173449
rect 87971 -173493 87979 -173449
rect 88071 -173493 88079 -173449
rect 88171 -173493 88179 -173449
rect 88271 -173493 88279 -173449
rect 88371 -173493 88379 -173449
rect 88471 -173493 88479 -173449
rect 88571 -173493 88579 -173449
rect 88671 -173493 88679 -173449
rect 88771 -173493 88779 -173449
rect 88871 -173493 88879 -173449
rect 88971 -173493 88979 -173449
rect 89071 -173493 89079 -173449
rect 89171 -173493 89179 -173449
rect 165525 -173489 165569 -173481
rect 165625 -173489 165669 -173481
rect 165725 -173489 165769 -173481
rect 165825 -173489 165869 -173481
rect 165925 -173489 165969 -173481
rect 166025 -173489 166069 -173481
rect 166125 -173489 166169 -173481
rect 166225 -173489 166269 -173481
rect 166325 -173489 166369 -173481
rect 166425 -173489 166469 -173481
rect 166525 -173489 166569 -173481
rect 166625 -173489 166669 -173481
rect 166725 -173489 166769 -173481
rect 166825 -173489 166869 -173481
rect 166925 -173489 166969 -173481
rect 167025 -173489 167069 -173481
rect 167525 -173489 167569 -173481
rect 167625 -173489 167669 -173481
rect 167725 -173489 167769 -173481
rect 167825 -173489 167869 -173481
rect 167925 -173489 167969 -173481
rect 168025 -173489 168069 -173481
rect 168125 -173489 168169 -173481
rect 168225 -173489 168269 -173481
rect 168325 -173489 168369 -173481
rect 168425 -173489 168469 -173481
rect 168525 -173489 168569 -173481
rect 168625 -173489 168669 -173481
rect 168725 -173489 168769 -173481
rect 168825 -173489 168869 -173481
rect 168925 -173489 168969 -173481
rect 169025 -173489 169069 -173481
rect 169525 -173489 169569 -173481
rect 169625 -173489 169669 -173481
rect 169725 -173489 169769 -173481
rect 169825 -173489 169869 -173481
rect 169925 -173489 169969 -173481
rect 170025 -173489 170069 -173481
rect 170125 -173489 170169 -173481
rect 170225 -173489 170269 -173481
rect 170325 -173489 170369 -173481
rect 170425 -173489 170469 -173481
rect 170525 -173489 170569 -173481
rect 170625 -173489 170669 -173481
rect 170725 -173489 170769 -173481
rect 170825 -173489 170869 -173481
rect 170925 -173489 170969 -173481
rect 171025 -173489 171069 -173481
rect 171525 -173489 171569 -173481
rect 171625 -173489 171669 -173481
rect 171725 -173489 171769 -173481
rect 171825 -173489 171869 -173481
rect 171925 -173489 171969 -173481
rect 172025 -173489 172069 -173481
rect 172125 -173489 172169 -173481
rect 172225 -173489 172269 -173481
rect 172325 -173489 172369 -173481
rect 172425 -173489 172469 -173481
rect 172525 -173489 172569 -173481
rect 172625 -173489 172669 -173481
rect 172725 -173489 172769 -173481
rect 172825 -173489 172869 -173481
rect 172925 -173489 172969 -173481
rect 173025 -173489 173069 -173481
rect 165569 -173533 165577 -173489
rect 165669 -173533 165677 -173489
rect 165769 -173533 165777 -173489
rect 165869 -173533 165877 -173489
rect 165969 -173533 165977 -173489
rect 166069 -173533 166077 -173489
rect 166169 -173533 166177 -173489
rect 166269 -173533 166277 -173489
rect 166369 -173533 166377 -173489
rect 166469 -173533 166477 -173489
rect 166569 -173533 166577 -173489
rect 166669 -173533 166677 -173489
rect 166769 -173533 166777 -173489
rect 166869 -173533 166877 -173489
rect 166969 -173533 166977 -173489
rect 167069 -173533 167077 -173489
rect 167569 -173533 167577 -173489
rect 167669 -173533 167677 -173489
rect 167769 -173533 167777 -173489
rect 167869 -173533 167877 -173489
rect 167969 -173533 167977 -173489
rect 168069 -173533 168077 -173489
rect 168169 -173533 168177 -173489
rect 168269 -173533 168277 -173489
rect 168369 -173533 168377 -173489
rect 168469 -173533 168477 -173489
rect 168569 -173533 168577 -173489
rect 168669 -173533 168677 -173489
rect 168769 -173533 168777 -173489
rect 168869 -173533 168877 -173489
rect 168969 -173533 168977 -173489
rect 169069 -173533 169077 -173489
rect 169569 -173533 169577 -173489
rect 169669 -173533 169677 -173489
rect 169769 -173533 169777 -173489
rect 169869 -173533 169877 -173489
rect 169969 -173533 169977 -173489
rect 170069 -173533 170077 -173489
rect 170169 -173533 170177 -173489
rect 170269 -173533 170277 -173489
rect 170369 -173533 170377 -173489
rect 170469 -173533 170477 -173489
rect 170569 -173533 170577 -173489
rect 170669 -173533 170677 -173489
rect 170769 -173533 170777 -173489
rect 170869 -173533 170877 -173489
rect 170969 -173533 170977 -173489
rect 171069 -173533 171077 -173489
rect 171569 -173533 171577 -173489
rect 171669 -173533 171677 -173489
rect 171769 -173533 171777 -173489
rect 171869 -173533 171877 -173489
rect 171969 -173533 171977 -173489
rect 172069 -173533 172077 -173489
rect 172169 -173533 172177 -173489
rect 172269 -173533 172277 -173489
rect 172369 -173533 172377 -173489
rect 172469 -173533 172477 -173489
rect 172569 -173533 172577 -173489
rect 172669 -173533 172677 -173489
rect 172769 -173533 172777 -173489
rect 172869 -173533 172877 -173489
rect 172969 -173533 172977 -173489
rect 173069 -173533 173077 -173489
rect 81627 -173549 81671 -173541
rect 81727 -173549 81771 -173541
rect 81827 -173549 81871 -173541
rect 81927 -173549 81971 -173541
rect 82027 -173549 82071 -173541
rect 82127 -173549 82171 -173541
rect 82227 -173549 82271 -173541
rect 82327 -173549 82371 -173541
rect 82427 -173549 82471 -173541
rect 82527 -173549 82571 -173541
rect 82627 -173549 82671 -173541
rect 82727 -173549 82771 -173541
rect 82827 -173549 82871 -173541
rect 82927 -173549 82971 -173541
rect 83027 -173549 83071 -173541
rect 83127 -173549 83171 -173541
rect 83627 -173549 83671 -173541
rect 83727 -173549 83771 -173541
rect 83827 -173549 83871 -173541
rect 83927 -173549 83971 -173541
rect 84027 -173549 84071 -173541
rect 84127 -173549 84171 -173541
rect 84227 -173549 84271 -173541
rect 84327 -173549 84371 -173541
rect 84427 -173549 84471 -173541
rect 84527 -173549 84571 -173541
rect 84627 -173549 84671 -173541
rect 84727 -173549 84771 -173541
rect 84827 -173549 84871 -173541
rect 84927 -173549 84971 -173541
rect 85027 -173549 85071 -173541
rect 85127 -173549 85171 -173541
rect 85627 -173549 85671 -173541
rect 85727 -173549 85771 -173541
rect 85827 -173549 85871 -173541
rect 85927 -173549 85971 -173541
rect 86027 -173549 86071 -173541
rect 86127 -173549 86171 -173541
rect 86227 -173549 86271 -173541
rect 86327 -173549 86371 -173541
rect 86427 -173549 86471 -173541
rect 86527 -173549 86571 -173541
rect 86627 -173549 86671 -173541
rect 86727 -173549 86771 -173541
rect 86827 -173549 86871 -173541
rect 86927 -173549 86971 -173541
rect 87027 -173549 87071 -173541
rect 87127 -173549 87171 -173541
rect 87627 -173549 87671 -173541
rect 87727 -173549 87771 -173541
rect 87827 -173549 87871 -173541
rect 87927 -173549 87971 -173541
rect 88027 -173549 88071 -173541
rect 88127 -173549 88171 -173541
rect 88227 -173549 88271 -173541
rect 88327 -173549 88371 -173541
rect 88427 -173549 88471 -173541
rect 88527 -173549 88571 -173541
rect 88627 -173549 88671 -173541
rect 88727 -173549 88771 -173541
rect 88827 -173549 88871 -173541
rect 88927 -173549 88971 -173541
rect 89027 -173549 89071 -173541
rect 89127 -173549 89171 -173541
rect 81671 -173593 81679 -173549
rect 81771 -173593 81779 -173549
rect 81871 -173593 81879 -173549
rect 81971 -173593 81979 -173549
rect 82071 -173593 82079 -173549
rect 82171 -173593 82179 -173549
rect 82271 -173593 82279 -173549
rect 82371 -173593 82379 -173549
rect 82471 -173593 82479 -173549
rect 82571 -173593 82579 -173549
rect 82671 -173593 82679 -173549
rect 82771 -173593 82779 -173549
rect 82871 -173593 82879 -173549
rect 82971 -173593 82979 -173549
rect 83071 -173593 83079 -173549
rect 83171 -173593 83179 -173549
rect 83671 -173593 83679 -173549
rect 83771 -173593 83779 -173549
rect 83871 -173593 83879 -173549
rect 83971 -173593 83979 -173549
rect 84071 -173593 84079 -173549
rect 84171 -173593 84179 -173549
rect 84271 -173593 84279 -173549
rect 84371 -173593 84379 -173549
rect 84471 -173593 84479 -173549
rect 84571 -173593 84579 -173549
rect 84671 -173593 84679 -173549
rect 84771 -173593 84779 -173549
rect 84871 -173593 84879 -173549
rect 84971 -173593 84979 -173549
rect 85071 -173593 85079 -173549
rect 85171 -173593 85179 -173549
rect 85671 -173593 85679 -173549
rect 85771 -173593 85779 -173549
rect 85871 -173593 85879 -173549
rect 85971 -173593 85979 -173549
rect 86071 -173593 86079 -173549
rect 86171 -173593 86179 -173549
rect 86271 -173593 86279 -173549
rect 86371 -173593 86379 -173549
rect 86471 -173593 86479 -173549
rect 86571 -173593 86579 -173549
rect 86671 -173593 86679 -173549
rect 86771 -173593 86779 -173549
rect 86871 -173593 86879 -173549
rect 86971 -173593 86979 -173549
rect 87071 -173593 87079 -173549
rect 87171 -173593 87179 -173549
rect 87671 -173593 87679 -173549
rect 87771 -173593 87779 -173549
rect 87871 -173593 87879 -173549
rect 87971 -173593 87979 -173549
rect 88071 -173593 88079 -173549
rect 88171 -173593 88179 -173549
rect 88271 -173593 88279 -173549
rect 88371 -173593 88379 -173549
rect 88471 -173593 88479 -173549
rect 88571 -173593 88579 -173549
rect 88671 -173593 88679 -173549
rect 88771 -173593 88779 -173549
rect 88871 -173593 88879 -173549
rect 88971 -173593 88979 -173549
rect 89071 -173593 89079 -173549
rect 89171 -173593 89179 -173549
rect 165525 -173589 165569 -173581
rect 165625 -173589 165669 -173581
rect 165725 -173589 165769 -173581
rect 165825 -173589 165869 -173581
rect 165925 -173589 165969 -173581
rect 166025 -173589 166069 -173581
rect 166125 -173589 166169 -173581
rect 166225 -173589 166269 -173581
rect 166325 -173589 166369 -173581
rect 166425 -173589 166469 -173581
rect 166525 -173589 166569 -173581
rect 166625 -173589 166669 -173581
rect 166725 -173589 166769 -173581
rect 166825 -173589 166869 -173581
rect 166925 -173589 166969 -173581
rect 167025 -173589 167069 -173581
rect 167525 -173589 167569 -173581
rect 167625 -173589 167669 -173581
rect 167725 -173589 167769 -173581
rect 167825 -173589 167869 -173581
rect 167925 -173589 167969 -173581
rect 168025 -173589 168069 -173581
rect 168125 -173589 168169 -173581
rect 168225 -173589 168269 -173581
rect 168325 -173589 168369 -173581
rect 168425 -173589 168469 -173581
rect 168525 -173589 168569 -173581
rect 168625 -173589 168669 -173581
rect 168725 -173589 168769 -173581
rect 168825 -173589 168869 -173581
rect 168925 -173589 168969 -173581
rect 169025 -173589 169069 -173581
rect 169525 -173589 169569 -173581
rect 169625 -173589 169669 -173581
rect 169725 -173589 169769 -173581
rect 169825 -173589 169869 -173581
rect 169925 -173589 169969 -173581
rect 170025 -173589 170069 -173581
rect 170125 -173589 170169 -173581
rect 170225 -173589 170269 -173581
rect 170325 -173589 170369 -173581
rect 170425 -173589 170469 -173581
rect 170525 -173589 170569 -173581
rect 170625 -173589 170669 -173581
rect 170725 -173589 170769 -173581
rect 170825 -173589 170869 -173581
rect 170925 -173589 170969 -173581
rect 171025 -173589 171069 -173581
rect 171525 -173589 171569 -173581
rect 171625 -173589 171669 -173581
rect 171725 -173589 171769 -173581
rect 171825 -173589 171869 -173581
rect 171925 -173589 171969 -173581
rect 172025 -173589 172069 -173581
rect 172125 -173589 172169 -173581
rect 172225 -173589 172269 -173581
rect 172325 -173589 172369 -173581
rect 172425 -173589 172469 -173581
rect 172525 -173589 172569 -173581
rect 172625 -173589 172669 -173581
rect 172725 -173589 172769 -173581
rect 172825 -173589 172869 -173581
rect 172925 -173589 172969 -173581
rect 173025 -173589 173069 -173581
rect 165569 -173633 165577 -173589
rect 165669 -173633 165677 -173589
rect 165769 -173633 165777 -173589
rect 165869 -173633 165877 -173589
rect 165969 -173633 165977 -173589
rect 166069 -173633 166077 -173589
rect 166169 -173633 166177 -173589
rect 166269 -173633 166277 -173589
rect 166369 -173633 166377 -173589
rect 166469 -173633 166477 -173589
rect 166569 -173633 166577 -173589
rect 166669 -173633 166677 -173589
rect 166769 -173633 166777 -173589
rect 166869 -173633 166877 -173589
rect 166969 -173633 166977 -173589
rect 167069 -173633 167077 -173589
rect 167569 -173633 167577 -173589
rect 167669 -173633 167677 -173589
rect 167769 -173633 167777 -173589
rect 167869 -173633 167877 -173589
rect 167969 -173633 167977 -173589
rect 168069 -173633 168077 -173589
rect 168169 -173633 168177 -173589
rect 168269 -173633 168277 -173589
rect 168369 -173633 168377 -173589
rect 168469 -173633 168477 -173589
rect 168569 -173633 168577 -173589
rect 168669 -173633 168677 -173589
rect 168769 -173633 168777 -173589
rect 168869 -173633 168877 -173589
rect 168969 -173633 168977 -173589
rect 169069 -173633 169077 -173589
rect 169569 -173633 169577 -173589
rect 169669 -173633 169677 -173589
rect 169769 -173633 169777 -173589
rect 169869 -173633 169877 -173589
rect 169969 -173633 169977 -173589
rect 170069 -173633 170077 -173589
rect 170169 -173633 170177 -173589
rect 170269 -173633 170277 -173589
rect 170369 -173633 170377 -173589
rect 170469 -173633 170477 -173589
rect 170569 -173633 170577 -173589
rect 170669 -173633 170677 -173589
rect 170769 -173633 170777 -173589
rect 170869 -173633 170877 -173589
rect 170969 -173633 170977 -173589
rect 171069 -173633 171077 -173589
rect 171569 -173633 171577 -173589
rect 171669 -173633 171677 -173589
rect 171769 -173633 171777 -173589
rect 171869 -173633 171877 -173589
rect 171969 -173633 171977 -173589
rect 172069 -173633 172077 -173589
rect 172169 -173633 172177 -173589
rect 172269 -173633 172277 -173589
rect 172369 -173633 172377 -173589
rect 172469 -173633 172477 -173589
rect 172569 -173633 172577 -173589
rect 172669 -173633 172677 -173589
rect 172769 -173633 172777 -173589
rect 172869 -173633 172877 -173589
rect 172969 -173633 172977 -173589
rect 173069 -173633 173077 -173589
rect 81627 -173649 81671 -173641
rect 81727 -173649 81771 -173641
rect 81827 -173649 81871 -173641
rect 81927 -173649 81971 -173641
rect 82027 -173649 82071 -173641
rect 82127 -173649 82171 -173641
rect 82227 -173649 82271 -173641
rect 82327 -173649 82371 -173641
rect 82427 -173649 82471 -173641
rect 82527 -173649 82571 -173641
rect 82627 -173649 82671 -173641
rect 82727 -173649 82771 -173641
rect 82827 -173649 82871 -173641
rect 82927 -173649 82971 -173641
rect 83027 -173649 83071 -173641
rect 83127 -173649 83171 -173641
rect 83627 -173649 83671 -173641
rect 83727 -173649 83771 -173641
rect 83827 -173649 83871 -173641
rect 83927 -173649 83971 -173641
rect 84027 -173649 84071 -173641
rect 84127 -173649 84171 -173641
rect 84227 -173649 84271 -173641
rect 84327 -173649 84371 -173641
rect 84427 -173649 84471 -173641
rect 84527 -173649 84571 -173641
rect 84627 -173649 84671 -173641
rect 84727 -173649 84771 -173641
rect 84827 -173649 84871 -173641
rect 84927 -173649 84971 -173641
rect 85027 -173649 85071 -173641
rect 85127 -173649 85171 -173641
rect 85627 -173649 85671 -173641
rect 85727 -173649 85771 -173641
rect 85827 -173649 85871 -173641
rect 85927 -173649 85971 -173641
rect 86027 -173649 86071 -173641
rect 86127 -173649 86171 -173641
rect 86227 -173649 86271 -173641
rect 86327 -173649 86371 -173641
rect 86427 -173649 86471 -173641
rect 86527 -173649 86571 -173641
rect 86627 -173649 86671 -173641
rect 86727 -173649 86771 -173641
rect 86827 -173649 86871 -173641
rect 86927 -173649 86971 -173641
rect 87027 -173649 87071 -173641
rect 87127 -173649 87171 -173641
rect 87627 -173649 87671 -173641
rect 87727 -173649 87771 -173641
rect 87827 -173649 87871 -173641
rect 87927 -173649 87971 -173641
rect 88027 -173649 88071 -173641
rect 88127 -173649 88171 -173641
rect 88227 -173649 88271 -173641
rect 88327 -173649 88371 -173641
rect 88427 -173649 88471 -173641
rect 88527 -173649 88571 -173641
rect 88627 -173649 88671 -173641
rect 88727 -173649 88771 -173641
rect 88827 -173649 88871 -173641
rect 88927 -173649 88971 -173641
rect 89027 -173649 89071 -173641
rect 89127 -173649 89171 -173641
rect 81671 -173693 81679 -173649
rect 81771 -173693 81779 -173649
rect 81871 -173693 81879 -173649
rect 81971 -173693 81979 -173649
rect 82071 -173693 82079 -173649
rect 82171 -173693 82179 -173649
rect 82271 -173693 82279 -173649
rect 82371 -173693 82379 -173649
rect 82471 -173693 82479 -173649
rect 82571 -173693 82579 -173649
rect 82671 -173693 82679 -173649
rect 82771 -173693 82779 -173649
rect 82871 -173693 82879 -173649
rect 82971 -173693 82979 -173649
rect 83071 -173693 83079 -173649
rect 83171 -173693 83179 -173649
rect 83671 -173693 83679 -173649
rect 83771 -173693 83779 -173649
rect 83871 -173693 83879 -173649
rect 83971 -173693 83979 -173649
rect 84071 -173693 84079 -173649
rect 84171 -173693 84179 -173649
rect 84271 -173693 84279 -173649
rect 84371 -173693 84379 -173649
rect 84471 -173693 84479 -173649
rect 84571 -173693 84579 -173649
rect 84671 -173693 84679 -173649
rect 84771 -173693 84779 -173649
rect 84871 -173693 84879 -173649
rect 84971 -173693 84979 -173649
rect 85071 -173693 85079 -173649
rect 85171 -173693 85179 -173649
rect 85671 -173693 85679 -173649
rect 85771 -173693 85779 -173649
rect 85871 -173693 85879 -173649
rect 85971 -173693 85979 -173649
rect 86071 -173693 86079 -173649
rect 86171 -173693 86179 -173649
rect 86271 -173693 86279 -173649
rect 86371 -173693 86379 -173649
rect 86471 -173693 86479 -173649
rect 86571 -173693 86579 -173649
rect 86671 -173693 86679 -173649
rect 86771 -173693 86779 -173649
rect 86871 -173693 86879 -173649
rect 86971 -173693 86979 -173649
rect 87071 -173693 87079 -173649
rect 87171 -173693 87179 -173649
rect 87671 -173693 87679 -173649
rect 87771 -173693 87779 -173649
rect 87871 -173693 87879 -173649
rect 87971 -173693 87979 -173649
rect 88071 -173693 88079 -173649
rect 88171 -173693 88179 -173649
rect 88271 -173693 88279 -173649
rect 88371 -173693 88379 -173649
rect 88471 -173693 88479 -173649
rect 88571 -173693 88579 -173649
rect 88671 -173693 88679 -173649
rect 88771 -173693 88779 -173649
rect 88871 -173693 88879 -173649
rect 88971 -173693 88979 -173649
rect 89071 -173693 89079 -173649
rect 89171 -173693 89179 -173649
rect 165525 -173689 165569 -173681
rect 165625 -173689 165669 -173681
rect 165725 -173689 165769 -173681
rect 165825 -173689 165869 -173681
rect 165925 -173689 165969 -173681
rect 166025 -173689 166069 -173681
rect 166125 -173689 166169 -173681
rect 166225 -173689 166269 -173681
rect 166325 -173689 166369 -173681
rect 166425 -173689 166469 -173681
rect 166525 -173689 166569 -173681
rect 166625 -173689 166669 -173681
rect 166725 -173689 166769 -173681
rect 166825 -173689 166869 -173681
rect 166925 -173689 166969 -173681
rect 167025 -173689 167069 -173681
rect 167525 -173689 167569 -173681
rect 167625 -173689 167669 -173681
rect 167725 -173689 167769 -173681
rect 167825 -173689 167869 -173681
rect 167925 -173689 167969 -173681
rect 168025 -173689 168069 -173681
rect 168125 -173689 168169 -173681
rect 168225 -173689 168269 -173681
rect 168325 -173689 168369 -173681
rect 168425 -173689 168469 -173681
rect 168525 -173689 168569 -173681
rect 168625 -173689 168669 -173681
rect 168725 -173689 168769 -173681
rect 168825 -173689 168869 -173681
rect 168925 -173689 168969 -173681
rect 169025 -173689 169069 -173681
rect 169525 -173689 169569 -173681
rect 169625 -173689 169669 -173681
rect 169725 -173689 169769 -173681
rect 169825 -173689 169869 -173681
rect 169925 -173689 169969 -173681
rect 170025 -173689 170069 -173681
rect 170125 -173689 170169 -173681
rect 170225 -173689 170269 -173681
rect 170325 -173689 170369 -173681
rect 170425 -173689 170469 -173681
rect 170525 -173689 170569 -173681
rect 170625 -173689 170669 -173681
rect 170725 -173689 170769 -173681
rect 170825 -173689 170869 -173681
rect 170925 -173689 170969 -173681
rect 171025 -173689 171069 -173681
rect 171525 -173689 171569 -173681
rect 171625 -173689 171669 -173681
rect 171725 -173689 171769 -173681
rect 171825 -173689 171869 -173681
rect 171925 -173689 171969 -173681
rect 172025 -173689 172069 -173681
rect 172125 -173689 172169 -173681
rect 172225 -173689 172269 -173681
rect 172325 -173689 172369 -173681
rect 172425 -173689 172469 -173681
rect 172525 -173689 172569 -173681
rect 172625 -173689 172669 -173681
rect 172725 -173689 172769 -173681
rect 172825 -173689 172869 -173681
rect 172925 -173689 172969 -173681
rect 173025 -173689 173069 -173681
rect 165569 -173733 165577 -173689
rect 165669 -173733 165677 -173689
rect 165769 -173733 165777 -173689
rect 165869 -173733 165877 -173689
rect 165969 -173733 165977 -173689
rect 166069 -173733 166077 -173689
rect 166169 -173733 166177 -173689
rect 166269 -173733 166277 -173689
rect 166369 -173733 166377 -173689
rect 166469 -173733 166477 -173689
rect 166569 -173733 166577 -173689
rect 166669 -173733 166677 -173689
rect 166769 -173733 166777 -173689
rect 166869 -173733 166877 -173689
rect 166969 -173733 166977 -173689
rect 167069 -173733 167077 -173689
rect 167569 -173733 167577 -173689
rect 167669 -173733 167677 -173689
rect 167769 -173733 167777 -173689
rect 167869 -173733 167877 -173689
rect 167969 -173733 167977 -173689
rect 168069 -173733 168077 -173689
rect 168169 -173733 168177 -173689
rect 168269 -173733 168277 -173689
rect 168369 -173733 168377 -173689
rect 168469 -173733 168477 -173689
rect 168569 -173733 168577 -173689
rect 168669 -173733 168677 -173689
rect 168769 -173733 168777 -173689
rect 168869 -173733 168877 -173689
rect 168969 -173733 168977 -173689
rect 169069 -173733 169077 -173689
rect 169569 -173733 169577 -173689
rect 169669 -173733 169677 -173689
rect 169769 -173733 169777 -173689
rect 169869 -173733 169877 -173689
rect 169969 -173733 169977 -173689
rect 170069 -173733 170077 -173689
rect 170169 -173733 170177 -173689
rect 170269 -173733 170277 -173689
rect 170369 -173733 170377 -173689
rect 170469 -173733 170477 -173689
rect 170569 -173733 170577 -173689
rect 170669 -173733 170677 -173689
rect 170769 -173733 170777 -173689
rect 170869 -173733 170877 -173689
rect 170969 -173733 170977 -173689
rect 171069 -173733 171077 -173689
rect 171569 -173733 171577 -173689
rect 171669 -173733 171677 -173689
rect 171769 -173733 171777 -173689
rect 171869 -173733 171877 -173689
rect 171969 -173733 171977 -173689
rect 172069 -173733 172077 -173689
rect 172169 -173733 172177 -173689
rect 172269 -173733 172277 -173689
rect 172369 -173733 172377 -173689
rect 172469 -173733 172477 -173689
rect 172569 -173733 172577 -173689
rect 172669 -173733 172677 -173689
rect 172769 -173733 172777 -173689
rect 172869 -173733 172877 -173689
rect 172969 -173733 172977 -173689
rect 173069 -173733 173077 -173689
rect 81627 -173749 81671 -173741
rect 81727 -173749 81771 -173741
rect 81827 -173749 81871 -173741
rect 81927 -173749 81971 -173741
rect 82027 -173749 82071 -173741
rect 82127 -173749 82171 -173741
rect 82227 -173749 82271 -173741
rect 82327 -173749 82371 -173741
rect 82427 -173749 82471 -173741
rect 82527 -173749 82571 -173741
rect 82627 -173749 82671 -173741
rect 82727 -173749 82771 -173741
rect 82827 -173749 82871 -173741
rect 82927 -173749 82971 -173741
rect 83027 -173749 83071 -173741
rect 83127 -173749 83171 -173741
rect 83627 -173749 83671 -173741
rect 83727 -173749 83771 -173741
rect 83827 -173749 83871 -173741
rect 83927 -173749 83971 -173741
rect 84027 -173749 84071 -173741
rect 84127 -173749 84171 -173741
rect 84227 -173749 84271 -173741
rect 84327 -173749 84371 -173741
rect 84427 -173749 84471 -173741
rect 84527 -173749 84571 -173741
rect 84627 -173749 84671 -173741
rect 84727 -173749 84771 -173741
rect 84827 -173749 84871 -173741
rect 84927 -173749 84971 -173741
rect 85027 -173749 85071 -173741
rect 85127 -173749 85171 -173741
rect 85627 -173749 85671 -173741
rect 85727 -173749 85771 -173741
rect 85827 -173749 85871 -173741
rect 85927 -173749 85971 -173741
rect 86027 -173749 86071 -173741
rect 86127 -173749 86171 -173741
rect 86227 -173749 86271 -173741
rect 86327 -173749 86371 -173741
rect 86427 -173749 86471 -173741
rect 86527 -173749 86571 -173741
rect 86627 -173749 86671 -173741
rect 86727 -173749 86771 -173741
rect 86827 -173749 86871 -173741
rect 86927 -173749 86971 -173741
rect 87027 -173749 87071 -173741
rect 87127 -173749 87171 -173741
rect 87627 -173749 87671 -173741
rect 87727 -173749 87771 -173741
rect 87827 -173749 87871 -173741
rect 87927 -173749 87971 -173741
rect 88027 -173749 88071 -173741
rect 88127 -173749 88171 -173741
rect 88227 -173749 88271 -173741
rect 88327 -173749 88371 -173741
rect 88427 -173749 88471 -173741
rect 88527 -173749 88571 -173741
rect 88627 -173749 88671 -173741
rect 88727 -173749 88771 -173741
rect 88827 -173749 88871 -173741
rect 88927 -173749 88971 -173741
rect 89027 -173749 89071 -173741
rect 89127 -173749 89171 -173741
rect 81671 -173793 81679 -173749
rect 81771 -173793 81779 -173749
rect 81871 -173793 81879 -173749
rect 81971 -173793 81979 -173749
rect 82071 -173793 82079 -173749
rect 82171 -173793 82179 -173749
rect 82271 -173793 82279 -173749
rect 82371 -173793 82379 -173749
rect 82471 -173793 82479 -173749
rect 82571 -173793 82579 -173749
rect 82671 -173793 82679 -173749
rect 82771 -173793 82779 -173749
rect 82871 -173793 82879 -173749
rect 82971 -173793 82979 -173749
rect 83071 -173793 83079 -173749
rect 83171 -173793 83179 -173749
rect 83671 -173793 83679 -173749
rect 83771 -173793 83779 -173749
rect 83871 -173793 83879 -173749
rect 83971 -173793 83979 -173749
rect 84071 -173793 84079 -173749
rect 84171 -173793 84179 -173749
rect 84271 -173793 84279 -173749
rect 84371 -173793 84379 -173749
rect 84471 -173793 84479 -173749
rect 84571 -173793 84579 -173749
rect 84671 -173793 84679 -173749
rect 84771 -173793 84779 -173749
rect 84871 -173793 84879 -173749
rect 84971 -173793 84979 -173749
rect 85071 -173793 85079 -173749
rect 85171 -173793 85179 -173749
rect 85671 -173793 85679 -173749
rect 85771 -173793 85779 -173749
rect 85871 -173793 85879 -173749
rect 85971 -173793 85979 -173749
rect 86071 -173793 86079 -173749
rect 86171 -173793 86179 -173749
rect 86271 -173793 86279 -173749
rect 86371 -173793 86379 -173749
rect 86471 -173793 86479 -173749
rect 86571 -173793 86579 -173749
rect 86671 -173793 86679 -173749
rect 86771 -173793 86779 -173749
rect 86871 -173793 86879 -173749
rect 86971 -173793 86979 -173749
rect 87071 -173793 87079 -173749
rect 87171 -173793 87179 -173749
rect 87671 -173793 87679 -173749
rect 87771 -173793 87779 -173749
rect 87871 -173793 87879 -173749
rect 87971 -173793 87979 -173749
rect 88071 -173793 88079 -173749
rect 88171 -173793 88179 -173749
rect 88271 -173793 88279 -173749
rect 88371 -173793 88379 -173749
rect 88471 -173793 88479 -173749
rect 88571 -173793 88579 -173749
rect 88671 -173793 88679 -173749
rect 88771 -173793 88779 -173749
rect 88871 -173793 88879 -173749
rect 88971 -173793 88979 -173749
rect 89071 -173793 89079 -173749
rect 89171 -173793 89179 -173749
rect 165525 -173789 165569 -173781
rect 165625 -173789 165669 -173781
rect 165725 -173789 165769 -173781
rect 165825 -173789 165869 -173781
rect 165925 -173789 165969 -173781
rect 166025 -173789 166069 -173781
rect 166125 -173789 166169 -173781
rect 166225 -173789 166269 -173781
rect 166325 -173789 166369 -173781
rect 166425 -173789 166469 -173781
rect 166525 -173789 166569 -173781
rect 166625 -173789 166669 -173781
rect 166725 -173789 166769 -173781
rect 166825 -173789 166869 -173781
rect 166925 -173789 166969 -173781
rect 167025 -173789 167069 -173781
rect 167525 -173789 167569 -173781
rect 167625 -173789 167669 -173781
rect 167725 -173789 167769 -173781
rect 167825 -173789 167869 -173781
rect 167925 -173789 167969 -173781
rect 168025 -173789 168069 -173781
rect 168125 -173789 168169 -173781
rect 168225 -173789 168269 -173781
rect 168325 -173789 168369 -173781
rect 168425 -173789 168469 -173781
rect 168525 -173789 168569 -173781
rect 168625 -173789 168669 -173781
rect 168725 -173789 168769 -173781
rect 168825 -173789 168869 -173781
rect 168925 -173789 168969 -173781
rect 169025 -173789 169069 -173781
rect 169525 -173789 169569 -173781
rect 169625 -173789 169669 -173781
rect 169725 -173789 169769 -173781
rect 169825 -173789 169869 -173781
rect 169925 -173789 169969 -173781
rect 170025 -173789 170069 -173781
rect 170125 -173789 170169 -173781
rect 170225 -173789 170269 -173781
rect 170325 -173789 170369 -173781
rect 170425 -173789 170469 -173781
rect 170525 -173789 170569 -173781
rect 170625 -173789 170669 -173781
rect 170725 -173789 170769 -173781
rect 170825 -173789 170869 -173781
rect 170925 -173789 170969 -173781
rect 171025 -173789 171069 -173781
rect 171525 -173789 171569 -173781
rect 171625 -173789 171669 -173781
rect 171725 -173789 171769 -173781
rect 171825 -173789 171869 -173781
rect 171925 -173789 171969 -173781
rect 172025 -173789 172069 -173781
rect 172125 -173789 172169 -173781
rect 172225 -173789 172269 -173781
rect 172325 -173789 172369 -173781
rect 172425 -173789 172469 -173781
rect 172525 -173789 172569 -173781
rect 172625 -173789 172669 -173781
rect 172725 -173789 172769 -173781
rect 172825 -173789 172869 -173781
rect 172925 -173789 172969 -173781
rect 173025 -173789 173069 -173781
rect 165569 -173833 165577 -173789
rect 165669 -173833 165677 -173789
rect 165769 -173833 165777 -173789
rect 165869 -173833 165877 -173789
rect 165969 -173833 165977 -173789
rect 166069 -173833 166077 -173789
rect 166169 -173833 166177 -173789
rect 166269 -173833 166277 -173789
rect 166369 -173833 166377 -173789
rect 166469 -173833 166477 -173789
rect 166569 -173833 166577 -173789
rect 166669 -173833 166677 -173789
rect 166769 -173833 166777 -173789
rect 166869 -173833 166877 -173789
rect 166969 -173833 166977 -173789
rect 167069 -173833 167077 -173789
rect 167569 -173833 167577 -173789
rect 167669 -173833 167677 -173789
rect 167769 -173833 167777 -173789
rect 167869 -173833 167877 -173789
rect 167969 -173833 167977 -173789
rect 168069 -173833 168077 -173789
rect 168169 -173833 168177 -173789
rect 168269 -173833 168277 -173789
rect 168369 -173833 168377 -173789
rect 168469 -173833 168477 -173789
rect 168569 -173833 168577 -173789
rect 168669 -173833 168677 -173789
rect 168769 -173833 168777 -173789
rect 168869 -173833 168877 -173789
rect 168969 -173833 168977 -173789
rect 169069 -173833 169077 -173789
rect 169569 -173833 169577 -173789
rect 169669 -173833 169677 -173789
rect 169769 -173833 169777 -173789
rect 169869 -173833 169877 -173789
rect 169969 -173833 169977 -173789
rect 170069 -173833 170077 -173789
rect 170169 -173833 170177 -173789
rect 170269 -173833 170277 -173789
rect 170369 -173833 170377 -173789
rect 170469 -173833 170477 -173789
rect 170569 -173833 170577 -173789
rect 170669 -173833 170677 -173789
rect 170769 -173833 170777 -173789
rect 170869 -173833 170877 -173789
rect 170969 -173833 170977 -173789
rect 171069 -173833 171077 -173789
rect 171569 -173833 171577 -173789
rect 171669 -173833 171677 -173789
rect 171769 -173833 171777 -173789
rect 171869 -173833 171877 -173789
rect 171969 -173833 171977 -173789
rect 172069 -173833 172077 -173789
rect 172169 -173833 172177 -173789
rect 172269 -173833 172277 -173789
rect 172369 -173833 172377 -173789
rect 172469 -173833 172477 -173789
rect 172569 -173833 172577 -173789
rect 172669 -173833 172677 -173789
rect 172769 -173833 172777 -173789
rect 172869 -173833 172877 -173789
rect 172969 -173833 172977 -173789
rect 173069 -173833 173077 -173789
rect 81627 -173849 81671 -173841
rect 81727 -173849 81771 -173841
rect 81827 -173849 81871 -173841
rect 81927 -173849 81971 -173841
rect 82027 -173849 82071 -173841
rect 82127 -173849 82171 -173841
rect 82227 -173849 82271 -173841
rect 82327 -173849 82371 -173841
rect 82427 -173849 82471 -173841
rect 82527 -173849 82571 -173841
rect 82627 -173849 82671 -173841
rect 82727 -173849 82771 -173841
rect 82827 -173849 82871 -173841
rect 82927 -173849 82971 -173841
rect 83027 -173849 83071 -173841
rect 83127 -173849 83171 -173841
rect 83627 -173849 83671 -173841
rect 83727 -173849 83771 -173841
rect 83827 -173849 83871 -173841
rect 83927 -173849 83971 -173841
rect 84027 -173849 84071 -173841
rect 84127 -173849 84171 -173841
rect 84227 -173849 84271 -173841
rect 84327 -173849 84371 -173841
rect 84427 -173849 84471 -173841
rect 84527 -173849 84571 -173841
rect 84627 -173849 84671 -173841
rect 84727 -173849 84771 -173841
rect 84827 -173849 84871 -173841
rect 84927 -173849 84971 -173841
rect 85027 -173849 85071 -173841
rect 85127 -173849 85171 -173841
rect 85627 -173849 85671 -173841
rect 85727 -173849 85771 -173841
rect 85827 -173849 85871 -173841
rect 85927 -173849 85971 -173841
rect 86027 -173849 86071 -173841
rect 86127 -173849 86171 -173841
rect 86227 -173849 86271 -173841
rect 86327 -173849 86371 -173841
rect 86427 -173849 86471 -173841
rect 86527 -173849 86571 -173841
rect 86627 -173849 86671 -173841
rect 86727 -173849 86771 -173841
rect 86827 -173849 86871 -173841
rect 86927 -173849 86971 -173841
rect 87027 -173849 87071 -173841
rect 87127 -173849 87171 -173841
rect 87627 -173849 87671 -173841
rect 87727 -173849 87771 -173841
rect 87827 -173849 87871 -173841
rect 87927 -173849 87971 -173841
rect 88027 -173849 88071 -173841
rect 88127 -173849 88171 -173841
rect 88227 -173849 88271 -173841
rect 88327 -173849 88371 -173841
rect 88427 -173849 88471 -173841
rect 88527 -173849 88571 -173841
rect 88627 -173849 88671 -173841
rect 88727 -173849 88771 -173841
rect 88827 -173849 88871 -173841
rect 88927 -173849 88971 -173841
rect 89027 -173849 89071 -173841
rect 89127 -173849 89171 -173841
rect 81671 -173893 81679 -173849
rect 81771 -173893 81779 -173849
rect 81871 -173893 81879 -173849
rect 81971 -173893 81979 -173849
rect 82071 -173893 82079 -173849
rect 82171 -173893 82179 -173849
rect 82271 -173893 82279 -173849
rect 82371 -173893 82379 -173849
rect 82471 -173893 82479 -173849
rect 82571 -173893 82579 -173849
rect 82671 -173893 82679 -173849
rect 82771 -173893 82779 -173849
rect 82871 -173893 82879 -173849
rect 82971 -173893 82979 -173849
rect 83071 -173893 83079 -173849
rect 83171 -173893 83179 -173849
rect 83671 -173893 83679 -173849
rect 83771 -173893 83779 -173849
rect 83871 -173893 83879 -173849
rect 83971 -173893 83979 -173849
rect 84071 -173893 84079 -173849
rect 84171 -173893 84179 -173849
rect 84271 -173893 84279 -173849
rect 84371 -173893 84379 -173849
rect 84471 -173893 84479 -173849
rect 84571 -173893 84579 -173849
rect 84671 -173893 84679 -173849
rect 84771 -173893 84779 -173849
rect 84871 -173893 84879 -173849
rect 84971 -173893 84979 -173849
rect 85071 -173893 85079 -173849
rect 85171 -173893 85179 -173849
rect 85671 -173893 85679 -173849
rect 85771 -173893 85779 -173849
rect 85871 -173893 85879 -173849
rect 85971 -173893 85979 -173849
rect 86071 -173893 86079 -173849
rect 86171 -173893 86179 -173849
rect 86271 -173893 86279 -173849
rect 86371 -173893 86379 -173849
rect 86471 -173893 86479 -173849
rect 86571 -173893 86579 -173849
rect 86671 -173893 86679 -173849
rect 86771 -173893 86779 -173849
rect 86871 -173893 86879 -173849
rect 86971 -173893 86979 -173849
rect 87071 -173893 87079 -173849
rect 87171 -173893 87179 -173849
rect 87671 -173893 87679 -173849
rect 87771 -173893 87779 -173849
rect 87871 -173893 87879 -173849
rect 87971 -173893 87979 -173849
rect 88071 -173893 88079 -173849
rect 88171 -173893 88179 -173849
rect 88271 -173893 88279 -173849
rect 88371 -173893 88379 -173849
rect 88471 -173893 88479 -173849
rect 88571 -173893 88579 -173849
rect 88671 -173893 88679 -173849
rect 88771 -173893 88779 -173849
rect 88871 -173893 88879 -173849
rect 88971 -173893 88979 -173849
rect 89071 -173893 89079 -173849
rect 89171 -173893 89179 -173849
rect 165525 -173889 165569 -173881
rect 165625 -173889 165669 -173881
rect 165725 -173889 165769 -173881
rect 165825 -173889 165869 -173881
rect 165925 -173889 165969 -173881
rect 166025 -173889 166069 -173881
rect 166125 -173889 166169 -173881
rect 166225 -173889 166269 -173881
rect 166325 -173889 166369 -173881
rect 166425 -173889 166469 -173881
rect 166525 -173889 166569 -173881
rect 166625 -173889 166669 -173881
rect 166725 -173889 166769 -173881
rect 166825 -173889 166869 -173881
rect 166925 -173889 166969 -173881
rect 167025 -173889 167069 -173881
rect 167525 -173889 167569 -173881
rect 167625 -173889 167669 -173881
rect 167725 -173889 167769 -173881
rect 167825 -173889 167869 -173881
rect 167925 -173889 167969 -173881
rect 168025 -173889 168069 -173881
rect 168125 -173889 168169 -173881
rect 168225 -173889 168269 -173881
rect 168325 -173889 168369 -173881
rect 168425 -173889 168469 -173881
rect 168525 -173889 168569 -173881
rect 168625 -173889 168669 -173881
rect 168725 -173889 168769 -173881
rect 168825 -173889 168869 -173881
rect 168925 -173889 168969 -173881
rect 169025 -173889 169069 -173881
rect 169525 -173889 169569 -173881
rect 169625 -173889 169669 -173881
rect 169725 -173889 169769 -173881
rect 169825 -173889 169869 -173881
rect 169925 -173889 169969 -173881
rect 170025 -173889 170069 -173881
rect 170125 -173889 170169 -173881
rect 170225 -173889 170269 -173881
rect 170325 -173889 170369 -173881
rect 170425 -173889 170469 -173881
rect 170525 -173889 170569 -173881
rect 170625 -173889 170669 -173881
rect 170725 -173889 170769 -173881
rect 170825 -173889 170869 -173881
rect 170925 -173889 170969 -173881
rect 171025 -173889 171069 -173881
rect 171525 -173889 171569 -173881
rect 171625 -173889 171669 -173881
rect 171725 -173889 171769 -173881
rect 171825 -173889 171869 -173881
rect 171925 -173889 171969 -173881
rect 172025 -173889 172069 -173881
rect 172125 -173889 172169 -173881
rect 172225 -173889 172269 -173881
rect 172325 -173889 172369 -173881
rect 172425 -173889 172469 -173881
rect 172525 -173889 172569 -173881
rect 172625 -173889 172669 -173881
rect 172725 -173889 172769 -173881
rect 172825 -173889 172869 -173881
rect 172925 -173889 172969 -173881
rect 173025 -173889 173069 -173881
rect 165569 -173933 165577 -173889
rect 165669 -173933 165677 -173889
rect 165769 -173933 165777 -173889
rect 165869 -173933 165877 -173889
rect 165969 -173933 165977 -173889
rect 166069 -173933 166077 -173889
rect 166169 -173933 166177 -173889
rect 166269 -173933 166277 -173889
rect 166369 -173933 166377 -173889
rect 166469 -173933 166477 -173889
rect 166569 -173933 166577 -173889
rect 166669 -173933 166677 -173889
rect 166769 -173933 166777 -173889
rect 166869 -173933 166877 -173889
rect 166969 -173933 166977 -173889
rect 167069 -173933 167077 -173889
rect 167569 -173933 167577 -173889
rect 167669 -173933 167677 -173889
rect 167769 -173933 167777 -173889
rect 167869 -173933 167877 -173889
rect 167969 -173933 167977 -173889
rect 168069 -173933 168077 -173889
rect 168169 -173933 168177 -173889
rect 168269 -173933 168277 -173889
rect 168369 -173933 168377 -173889
rect 168469 -173933 168477 -173889
rect 168569 -173933 168577 -173889
rect 168669 -173933 168677 -173889
rect 168769 -173933 168777 -173889
rect 168869 -173933 168877 -173889
rect 168969 -173933 168977 -173889
rect 169069 -173933 169077 -173889
rect 169569 -173933 169577 -173889
rect 169669 -173933 169677 -173889
rect 169769 -173933 169777 -173889
rect 169869 -173933 169877 -173889
rect 169969 -173933 169977 -173889
rect 170069 -173933 170077 -173889
rect 170169 -173933 170177 -173889
rect 170269 -173933 170277 -173889
rect 170369 -173933 170377 -173889
rect 170469 -173933 170477 -173889
rect 170569 -173933 170577 -173889
rect 170669 -173933 170677 -173889
rect 170769 -173933 170777 -173889
rect 170869 -173933 170877 -173889
rect 170969 -173933 170977 -173889
rect 171069 -173933 171077 -173889
rect 171569 -173933 171577 -173889
rect 171669 -173933 171677 -173889
rect 171769 -173933 171777 -173889
rect 171869 -173933 171877 -173889
rect 171969 -173933 171977 -173889
rect 172069 -173933 172077 -173889
rect 172169 -173933 172177 -173889
rect 172269 -173933 172277 -173889
rect 172369 -173933 172377 -173889
rect 172469 -173933 172477 -173889
rect 172569 -173933 172577 -173889
rect 172669 -173933 172677 -173889
rect 172769 -173933 172777 -173889
rect 172869 -173933 172877 -173889
rect 172969 -173933 172977 -173889
rect 173069 -173933 173077 -173889
rect 81627 -173949 81671 -173941
rect 81727 -173949 81771 -173941
rect 81827 -173949 81871 -173941
rect 81927 -173949 81971 -173941
rect 82027 -173949 82071 -173941
rect 82127 -173949 82171 -173941
rect 82227 -173949 82271 -173941
rect 82327 -173949 82371 -173941
rect 82427 -173949 82471 -173941
rect 82527 -173949 82571 -173941
rect 82627 -173949 82671 -173941
rect 82727 -173949 82771 -173941
rect 82827 -173949 82871 -173941
rect 82927 -173949 82971 -173941
rect 83027 -173949 83071 -173941
rect 83127 -173949 83171 -173941
rect 83627 -173949 83671 -173941
rect 83727 -173949 83771 -173941
rect 83827 -173949 83871 -173941
rect 83927 -173949 83971 -173941
rect 84027 -173949 84071 -173941
rect 84127 -173949 84171 -173941
rect 84227 -173949 84271 -173941
rect 84327 -173949 84371 -173941
rect 84427 -173949 84471 -173941
rect 84527 -173949 84571 -173941
rect 84627 -173949 84671 -173941
rect 84727 -173949 84771 -173941
rect 84827 -173949 84871 -173941
rect 84927 -173949 84971 -173941
rect 85027 -173949 85071 -173941
rect 85127 -173949 85171 -173941
rect 85627 -173949 85671 -173941
rect 85727 -173949 85771 -173941
rect 85827 -173949 85871 -173941
rect 85927 -173949 85971 -173941
rect 86027 -173949 86071 -173941
rect 86127 -173949 86171 -173941
rect 86227 -173949 86271 -173941
rect 86327 -173949 86371 -173941
rect 86427 -173949 86471 -173941
rect 86527 -173949 86571 -173941
rect 86627 -173949 86671 -173941
rect 86727 -173949 86771 -173941
rect 86827 -173949 86871 -173941
rect 86927 -173949 86971 -173941
rect 87027 -173949 87071 -173941
rect 87127 -173949 87171 -173941
rect 87627 -173949 87671 -173941
rect 87727 -173949 87771 -173941
rect 87827 -173949 87871 -173941
rect 87927 -173949 87971 -173941
rect 88027 -173949 88071 -173941
rect 88127 -173949 88171 -173941
rect 88227 -173949 88271 -173941
rect 88327 -173949 88371 -173941
rect 88427 -173949 88471 -173941
rect 88527 -173949 88571 -173941
rect 88627 -173949 88671 -173941
rect 88727 -173949 88771 -173941
rect 88827 -173949 88871 -173941
rect 88927 -173949 88971 -173941
rect 89027 -173949 89071 -173941
rect 89127 -173949 89171 -173941
rect 81671 -173993 81679 -173949
rect 81771 -173993 81779 -173949
rect 81871 -173993 81879 -173949
rect 81971 -173993 81979 -173949
rect 82071 -173993 82079 -173949
rect 82171 -173993 82179 -173949
rect 82271 -173993 82279 -173949
rect 82371 -173993 82379 -173949
rect 82471 -173993 82479 -173949
rect 82571 -173993 82579 -173949
rect 82671 -173993 82679 -173949
rect 82771 -173993 82779 -173949
rect 82871 -173993 82879 -173949
rect 82971 -173993 82979 -173949
rect 83071 -173993 83079 -173949
rect 83171 -173993 83179 -173949
rect 83671 -173993 83679 -173949
rect 83771 -173993 83779 -173949
rect 83871 -173993 83879 -173949
rect 83971 -173993 83979 -173949
rect 84071 -173993 84079 -173949
rect 84171 -173993 84179 -173949
rect 84271 -173993 84279 -173949
rect 84371 -173993 84379 -173949
rect 84471 -173993 84479 -173949
rect 84571 -173993 84579 -173949
rect 84671 -173993 84679 -173949
rect 84771 -173993 84779 -173949
rect 84871 -173993 84879 -173949
rect 84971 -173993 84979 -173949
rect 85071 -173993 85079 -173949
rect 85171 -173993 85179 -173949
rect 85671 -173993 85679 -173949
rect 85771 -173993 85779 -173949
rect 85871 -173993 85879 -173949
rect 85971 -173993 85979 -173949
rect 86071 -173993 86079 -173949
rect 86171 -173993 86179 -173949
rect 86271 -173993 86279 -173949
rect 86371 -173993 86379 -173949
rect 86471 -173993 86479 -173949
rect 86571 -173993 86579 -173949
rect 86671 -173993 86679 -173949
rect 86771 -173993 86779 -173949
rect 86871 -173993 86879 -173949
rect 86971 -173993 86979 -173949
rect 87071 -173993 87079 -173949
rect 87171 -173993 87179 -173949
rect 87671 -173993 87679 -173949
rect 87771 -173993 87779 -173949
rect 87871 -173993 87879 -173949
rect 87971 -173993 87979 -173949
rect 88071 -173993 88079 -173949
rect 88171 -173993 88179 -173949
rect 88271 -173993 88279 -173949
rect 88371 -173993 88379 -173949
rect 88471 -173993 88479 -173949
rect 88571 -173993 88579 -173949
rect 88671 -173993 88679 -173949
rect 88771 -173993 88779 -173949
rect 88871 -173993 88879 -173949
rect 88971 -173993 88979 -173949
rect 89071 -173993 89079 -173949
rect 89171 -173993 89179 -173949
rect 165525 -173989 165569 -173981
rect 165625 -173989 165669 -173981
rect 165725 -173989 165769 -173981
rect 165825 -173989 165869 -173981
rect 165925 -173989 165969 -173981
rect 166025 -173989 166069 -173981
rect 166125 -173989 166169 -173981
rect 166225 -173989 166269 -173981
rect 166325 -173989 166369 -173981
rect 166425 -173989 166469 -173981
rect 166525 -173989 166569 -173981
rect 166625 -173989 166669 -173981
rect 166725 -173989 166769 -173981
rect 166825 -173989 166869 -173981
rect 166925 -173989 166969 -173981
rect 167025 -173989 167069 -173981
rect 167525 -173989 167569 -173981
rect 167625 -173989 167669 -173981
rect 167725 -173989 167769 -173981
rect 167825 -173989 167869 -173981
rect 167925 -173989 167969 -173981
rect 168025 -173989 168069 -173981
rect 168125 -173989 168169 -173981
rect 168225 -173989 168269 -173981
rect 168325 -173989 168369 -173981
rect 168425 -173989 168469 -173981
rect 168525 -173989 168569 -173981
rect 168625 -173989 168669 -173981
rect 168725 -173989 168769 -173981
rect 168825 -173989 168869 -173981
rect 168925 -173989 168969 -173981
rect 169025 -173989 169069 -173981
rect 169525 -173989 169569 -173981
rect 169625 -173989 169669 -173981
rect 169725 -173989 169769 -173981
rect 169825 -173989 169869 -173981
rect 169925 -173989 169969 -173981
rect 170025 -173989 170069 -173981
rect 170125 -173989 170169 -173981
rect 170225 -173989 170269 -173981
rect 170325 -173989 170369 -173981
rect 170425 -173989 170469 -173981
rect 170525 -173989 170569 -173981
rect 170625 -173989 170669 -173981
rect 170725 -173989 170769 -173981
rect 170825 -173989 170869 -173981
rect 170925 -173989 170969 -173981
rect 171025 -173989 171069 -173981
rect 171525 -173989 171569 -173981
rect 171625 -173989 171669 -173981
rect 171725 -173989 171769 -173981
rect 171825 -173989 171869 -173981
rect 171925 -173989 171969 -173981
rect 172025 -173989 172069 -173981
rect 172125 -173989 172169 -173981
rect 172225 -173989 172269 -173981
rect 172325 -173989 172369 -173981
rect 172425 -173989 172469 -173981
rect 172525 -173989 172569 -173981
rect 172625 -173989 172669 -173981
rect 172725 -173989 172769 -173981
rect 172825 -173989 172869 -173981
rect 172925 -173989 172969 -173981
rect 173025 -173989 173069 -173981
rect 165569 -174033 165577 -173989
rect 165669 -174033 165677 -173989
rect 165769 -174033 165777 -173989
rect 165869 -174033 165877 -173989
rect 165969 -174033 165977 -173989
rect 166069 -174033 166077 -173989
rect 166169 -174033 166177 -173989
rect 166269 -174033 166277 -173989
rect 166369 -174033 166377 -173989
rect 166469 -174033 166477 -173989
rect 166569 -174033 166577 -173989
rect 166669 -174033 166677 -173989
rect 166769 -174033 166777 -173989
rect 166869 -174033 166877 -173989
rect 166969 -174033 166977 -173989
rect 167069 -174033 167077 -173989
rect 167569 -174033 167577 -173989
rect 167669 -174033 167677 -173989
rect 167769 -174033 167777 -173989
rect 167869 -174033 167877 -173989
rect 167969 -174033 167977 -173989
rect 168069 -174033 168077 -173989
rect 168169 -174033 168177 -173989
rect 168269 -174033 168277 -173989
rect 168369 -174033 168377 -173989
rect 168469 -174033 168477 -173989
rect 168569 -174033 168577 -173989
rect 168669 -174033 168677 -173989
rect 168769 -174033 168777 -173989
rect 168869 -174033 168877 -173989
rect 168969 -174033 168977 -173989
rect 169069 -174033 169077 -173989
rect 169569 -174033 169577 -173989
rect 169669 -174033 169677 -173989
rect 169769 -174033 169777 -173989
rect 169869 -174033 169877 -173989
rect 169969 -174033 169977 -173989
rect 170069 -174033 170077 -173989
rect 170169 -174033 170177 -173989
rect 170269 -174033 170277 -173989
rect 170369 -174033 170377 -173989
rect 170469 -174033 170477 -173989
rect 170569 -174033 170577 -173989
rect 170669 -174033 170677 -173989
rect 170769 -174033 170777 -173989
rect 170869 -174033 170877 -173989
rect 170969 -174033 170977 -173989
rect 171069 -174033 171077 -173989
rect 171569 -174033 171577 -173989
rect 171669 -174033 171677 -173989
rect 171769 -174033 171777 -173989
rect 171869 -174033 171877 -173989
rect 171969 -174033 171977 -173989
rect 172069 -174033 172077 -173989
rect 172169 -174033 172177 -173989
rect 172269 -174033 172277 -173989
rect 172369 -174033 172377 -173989
rect 172469 -174033 172477 -173989
rect 172569 -174033 172577 -173989
rect 172669 -174033 172677 -173989
rect 172769 -174033 172777 -173989
rect 172869 -174033 172877 -173989
rect 172969 -174033 172977 -173989
rect 173069 -174033 173077 -173989
rect 81627 -174049 81671 -174041
rect 81727 -174049 81771 -174041
rect 81827 -174049 81871 -174041
rect 81927 -174049 81971 -174041
rect 82027 -174049 82071 -174041
rect 82127 -174049 82171 -174041
rect 82227 -174049 82271 -174041
rect 82327 -174049 82371 -174041
rect 82427 -174049 82471 -174041
rect 82527 -174049 82571 -174041
rect 82627 -174049 82671 -174041
rect 82727 -174049 82771 -174041
rect 82827 -174049 82871 -174041
rect 82927 -174049 82971 -174041
rect 83027 -174049 83071 -174041
rect 83127 -174049 83171 -174041
rect 83627 -174049 83671 -174041
rect 83727 -174049 83771 -174041
rect 83827 -174049 83871 -174041
rect 83927 -174049 83971 -174041
rect 84027 -174049 84071 -174041
rect 84127 -174049 84171 -174041
rect 84227 -174049 84271 -174041
rect 84327 -174049 84371 -174041
rect 84427 -174049 84471 -174041
rect 84527 -174049 84571 -174041
rect 84627 -174049 84671 -174041
rect 84727 -174049 84771 -174041
rect 84827 -174049 84871 -174041
rect 84927 -174049 84971 -174041
rect 85027 -174049 85071 -174041
rect 85127 -174049 85171 -174041
rect 85627 -174049 85671 -174041
rect 85727 -174049 85771 -174041
rect 85827 -174049 85871 -174041
rect 85927 -174049 85971 -174041
rect 86027 -174049 86071 -174041
rect 86127 -174049 86171 -174041
rect 86227 -174049 86271 -174041
rect 86327 -174049 86371 -174041
rect 86427 -174049 86471 -174041
rect 86527 -174049 86571 -174041
rect 86627 -174049 86671 -174041
rect 86727 -174049 86771 -174041
rect 86827 -174049 86871 -174041
rect 86927 -174049 86971 -174041
rect 87027 -174049 87071 -174041
rect 87127 -174049 87171 -174041
rect 87627 -174049 87671 -174041
rect 87727 -174049 87771 -174041
rect 87827 -174049 87871 -174041
rect 87927 -174049 87971 -174041
rect 88027 -174049 88071 -174041
rect 88127 -174049 88171 -174041
rect 88227 -174049 88271 -174041
rect 88327 -174049 88371 -174041
rect 88427 -174049 88471 -174041
rect 88527 -174049 88571 -174041
rect 88627 -174049 88671 -174041
rect 88727 -174049 88771 -174041
rect 88827 -174049 88871 -174041
rect 88927 -174049 88971 -174041
rect 89027 -174049 89071 -174041
rect 89127 -174049 89171 -174041
rect 81671 -174093 81679 -174049
rect 81771 -174093 81779 -174049
rect 81871 -174093 81879 -174049
rect 81971 -174093 81979 -174049
rect 82071 -174093 82079 -174049
rect 82171 -174093 82179 -174049
rect 82271 -174093 82279 -174049
rect 82371 -174093 82379 -174049
rect 82471 -174093 82479 -174049
rect 82571 -174093 82579 -174049
rect 82671 -174093 82679 -174049
rect 82771 -174093 82779 -174049
rect 82871 -174093 82879 -174049
rect 82971 -174093 82979 -174049
rect 83071 -174093 83079 -174049
rect 83171 -174093 83179 -174049
rect 83671 -174093 83679 -174049
rect 83771 -174093 83779 -174049
rect 83871 -174093 83879 -174049
rect 83971 -174093 83979 -174049
rect 84071 -174093 84079 -174049
rect 84171 -174093 84179 -174049
rect 84271 -174093 84279 -174049
rect 84371 -174093 84379 -174049
rect 84471 -174093 84479 -174049
rect 84571 -174093 84579 -174049
rect 84671 -174093 84679 -174049
rect 84771 -174093 84779 -174049
rect 84871 -174093 84879 -174049
rect 84971 -174093 84979 -174049
rect 85071 -174093 85079 -174049
rect 85171 -174093 85179 -174049
rect 85671 -174093 85679 -174049
rect 85771 -174093 85779 -174049
rect 85871 -174093 85879 -174049
rect 85971 -174093 85979 -174049
rect 86071 -174093 86079 -174049
rect 86171 -174093 86179 -174049
rect 86271 -174093 86279 -174049
rect 86371 -174093 86379 -174049
rect 86471 -174093 86479 -174049
rect 86571 -174093 86579 -174049
rect 86671 -174093 86679 -174049
rect 86771 -174093 86779 -174049
rect 86871 -174093 86879 -174049
rect 86971 -174093 86979 -174049
rect 87071 -174093 87079 -174049
rect 87171 -174093 87179 -174049
rect 87671 -174093 87679 -174049
rect 87771 -174093 87779 -174049
rect 87871 -174093 87879 -174049
rect 87971 -174093 87979 -174049
rect 88071 -174093 88079 -174049
rect 88171 -174093 88179 -174049
rect 88271 -174093 88279 -174049
rect 88371 -174093 88379 -174049
rect 88471 -174093 88479 -174049
rect 88571 -174093 88579 -174049
rect 88671 -174093 88679 -174049
rect 88771 -174093 88779 -174049
rect 88871 -174093 88879 -174049
rect 88971 -174093 88979 -174049
rect 89071 -174093 89079 -174049
rect 89171 -174093 89179 -174049
rect 165525 -174089 165569 -174081
rect 165625 -174089 165669 -174081
rect 165725 -174089 165769 -174081
rect 165825 -174089 165869 -174081
rect 165925 -174089 165969 -174081
rect 166025 -174089 166069 -174081
rect 166125 -174089 166169 -174081
rect 166225 -174089 166269 -174081
rect 166325 -174089 166369 -174081
rect 166425 -174089 166469 -174081
rect 166525 -174089 166569 -174081
rect 166625 -174089 166669 -174081
rect 166725 -174089 166769 -174081
rect 166825 -174089 166869 -174081
rect 166925 -174089 166969 -174081
rect 167025 -174089 167069 -174081
rect 167525 -174089 167569 -174081
rect 167625 -174089 167669 -174081
rect 167725 -174089 167769 -174081
rect 167825 -174089 167869 -174081
rect 167925 -174089 167969 -174081
rect 168025 -174089 168069 -174081
rect 168125 -174089 168169 -174081
rect 168225 -174089 168269 -174081
rect 168325 -174089 168369 -174081
rect 168425 -174089 168469 -174081
rect 168525 -174089 168569 -174081
rect 168625 -174089 168669 -174081
rect 168725 -174089 168769 -174081
rect 168825 -174089 168869 -174081
rect 168925 -174089 168969 -174081
rect 169025 -174089 169069 -174081
rect 169525 -174089 169569 -174081
rect 169625 -174089 169669 -174081
rect 169725 -174089 169769 -174081
rect 169825 -174089 169869 -174081
rect 169925 -174089 169969 -174081
rect 170025 -174089 170069 -174081
rect 170125 -174089 170169 -174081
rect 170225 -174089 170269 -174081
rect 170325 -174089 170369 -174081
rect 170425 -174089 170469 -174081
rect 170525 -174089 170569 -174081
rect 170625 -174089 170669 -174081
rect 170725 -174089 170769 -174081
rect 170825 -174089 170869 -174081
rect 170925 -174089 170969 -174081
rect 171025 -174089 171069 -174081
rect 171525 -174089 171569 -174081
rect 171625 -174089 171669 -174081
rect 171725 -174089 171769 -174081
rect 171825 -174089 171869 -174081
rect 171925 -174089 171969 -174081
rect 172025 -174089 172069 -174081
rect 172125 -174089 172169 -174081
rect 172225 -174089 172269 -174081
rect 172325 -174089 172369 -174081
rect 172425 -174089 172469 -174081
rect 172525 -174089 172569 -174081
rect 172625 -174089 172669 -174081
rect 172725 -174089 172769 -174081
rect 172825 -174089 172869 -174081
rect 172925 -174089 172969 -174081
rect 173025 -174089 173069 -174081
rect 165569 -174133 165577 -174089
rect 165669 -174133 165677 -174089
rect 165769 -174133 165777 -174089
rect 165869 -174133 165877 -174089
rect 165969 -174133 165977 -174089
rect 166069 -174133 166077 -174089
rect 166169 -174133 166177 -174089
rect 166269 -174133 166277 -174089
rect 166369 -174133 166377 -174089
rect 166469 -174133 166477 -174089
rect 166569 -174133 166577 -174089
rect 166669 -174133 166677 -174089
rect 166769 -174133 166777 -174089
rect 166869 -174133 166877 -174089
rect 166969 -174133 166977 -174089
rect 167069 -174133 167077 -174089
rect 167569 -174133 167577 -174089
rect 167669 -174133 167677 -174089
rect 167769 -174133 167777 -174089
rect 167869 -174133 167877 -174089
rect 167969 -174133 167977 -174089
rect 168069 -174133 168077 -174089
rect 168169 -174133 168177 -174089
rect 168269 -174133 168277 -174089
rect 168369 -174133 168377 -174089
rect 168469 -174133 168477 -174089
rect 168569 -174133 168577 -174089
rect 168669 -174133 168677 -174089
rect 168769 -174133 168777 -174089
rect 168869 -174133 168877 -174089
rect 168969 -174133 168977 -174089
rect 169069 -174133 169077 -174089
rect 169569 -174133 169577 -174089
rect 169669 -174133 169677 -174089
rect 169769 -174133 169777 -174089
rect 169869 -174133 169877 -174089
rect 169969 -174133 169977 -174089
rect 170069 -174133 170077 -174089
rect 170169 -174133 170177 -174089
rect 170269 -174133 170277 -174089
rect 170369 -174133 170377 -174089
rect 170469 -174133 170477 -174089
rect 170569 -174133 170577 -174089
rect 170669 -174133 170677 -174089
rect 170769 -174133 170777 -174089
rect 170869 -174133 170877 -174089
rect 170969 -174133 170977 -174089
rect 171069 -174133 171077 -174089
rect 171569 -174133 171577 -174089
rect 171669 -174133 171677 -174089
rect 171769 -174133 171777 -174089
rect 171869 -174133 171877 -174089
rect 171969 -174133 171977 -174089
rect 172069 -174133 172077 -174089
rect 172169 -174133 172177 -174089
rect 172269 -174133 172277 -174089
rect 172369 -174133 172377 -174089
rect 172469 -174133 172477 -174089
rect 172569 -174133 172577 -174089
rect 172669 -174133 172677 -174089
rect 172769 -174133 172777 -174089
rect 172869 -174133 172877 -174089
rect 172969 -174133 172977 -174089
rect 173069 -174133 173077 -174089
rect 81627 -174149 81671 -174141
rect 81727 -174149 81771 -174141
rect 81827 -174149 81871 -174141
rect 81927 -174149 81971 -174141
rect 82027 -174149 82071 -174141
rect 82127 -174149 82171 -174141
rect 82227 -174149 82271 -174141
rect 82327 -174149 82371 -174141
rect 82427 -174149 82471 -174141
rect 82527 -174149 82571 -174141
rect 82627 -174149 82671 -174141
rect 82727 -174149 82771 -174141
rect 82827 -174149 82871 -174141
rect 82927 -174149 82971 -174141
rect 83027 -174149 83071 -174141
rect 83127 -174149 83171 -174141
rect 83627 -174149 83671 -174141
rect 83727 -174149 83771 -174141
rect 83827 -174149 83871 -174141
rect 83927 -174149 83971 -174141
rect 84027 -174149 84071 -174141
rect 84127 -174149 84171 -174141
rect 84227 -174149 84271 -174141
rect 84327 -174149 84371 -174141
rect 84427 -174149 84471 -174141
rect 84527 -174149 84571 -174141
rect 84627 -174149 84671 -174141
rect 84727 -174149 84771 -174141
rect 84827 -174149 84871 -174141
rect 84927 -174149 84971 -174141
rect 85027 -174149 85071 -174141
rect 85127 -174149 85171 -174141
rect 85627 -174149 85671 -174141
rect 85727 -174149 85771 -174141
rect 85827 -174149 85871 -174141
rect 85927 -174149 85971 -174141
rect 86027 -174149 86071 -174141
rect 86127 -174149 86171 -174141
rect 86227 -174149 86271 -174141
rect 86327 -174149 86371 -174141
rect 86427 -174149 86471 -174141
rect 86527 -174149 86571 -174141
rect 86627 -174149 86671 -174141
rect 86727 -174149 86771 -174141
rect 86827 -174149 86871 -174141
rect 86927 -174149 86971 -174141
rect 87027 -174149 87071 -174141
rect 87127 -174149 87171 -174141
rect 87627 -174149 87671 -174141
rect 87727 -174149 87771 -174141
rect 87827 -174149 87871 -174141
rect 87927 -174149 87971 -174141
rect 88027 -174149 88071 -174141
rect 88127 -174149 88171 -174141
rect 88227 -174149 88271 -174141
rect 88327 -174149 88371 -174141
rect 88427 -174149 88471 -174141
rect 88527 -174149 88571 -174141
rect 88627 -174149 88671 -174141
rect 88727 -174149 88771 -174141
rect 88827 -174149 88871 -174141
rect 88927 -174149 88971 -174141
rect 89027 -174149 89071 -174141
rect 89127 -174149 89171 -174141
rect 81671 -174193 81679 -174149
rect 81771 -174193 81779 -174149
rect 81871 -174193 81879 -174149
rect 81971 -174193 81979 -174149
rect 82071 -174193 82079 -174149
rect 82171 -174193 82179 -174149
rect 82271 -174193 82279 -174149
rect 82371 -174193 82379 -174149
rect 82471 -174193 82479 -174149
rect 82571 -174193 82579 -174149
rect 82671 -174193 82679 -174149
rect 82771 -174193 82779 -174149
rect 82871 -174193 82879 -174149
rect 82971 -174193 82979 -174149
rect 83071 -174193 83079 -174149
rect 83171 -174193 83179 -174149
rect 83671 -174193 83679 -174149
rect 83771 -174193 83779 -174149
rect 83871 -174193 83879 -174149
rect 83971 -174193 83979 -174149
rect 84071 -174193 84079 -174149
rect 84171 -174193 84179 -174149
rect 84271 -174193 84279 -174149
rect 84371 -174193 84379 -174149
rect 84471 -174193 84479 -174149
rect 84571 -174193 84579 -174149
rect 84671 -174193 84679 -174149
rect 84771 -174193 84779 -174149
rect 84871 -174193 84879 -174149
rect 84971 -174193 84979 -174149
rect 85071 -174193 85079 -174149
rect 85171 -174193 85179 -174149
rect 85671 -174193 85679 -174149
rect 85771 -174193 85779 -174149
rect 85871 -174193 85879 -174149
rect 85971 -174193 85979 -174149
rect 86071 -174193 86079 -174149
rect 86171 -174193 86179 -174149
rect 86271 -174193 86279 -174149
rect 86371 -174193 86379 -174149
rect 86471 -174193 86479 -174149
rect 86571 -174193 86579 -174149
rect 86671 -174193 86679 -174149
rect 86771 -174193 86779 -174149
rect 86871 -174193 86879 -174149
rect 86971 -174193 86979 -174149
rect 87071 -174193 87079 -174149
rect 87171 -174193 87179 -174149
rect 87671 -174193 87679 -174149
rect 87771 -174193 87779 -174149
rect 87871 -174193 87879 -174149
rect 87971 -174193 87979 -174149
rect 88071 -174193 88079 -174149
rect 88171 -174193 88179 -174149
rect 88271 -174193 88279 -174149
rect 88371 -174193 88379 -174149
rect 88471 -174193 88479 -174149
rect 88571 -174193 88579 -174149
rect 88671 -174193 88679 -174149
rect 88771 -174193 88779 -174149
rect 88871 -174193 88879 -174149
rect 88971 -174193 88979 -174149
rect 89071 -174193 89079 -174149
rect 89171 -174193 89179 -174149
rect 165525 -174189 165569 -174181
rect 165625 -174189 165669 -174181
rect 165725 -174189 165769 -174181
rect 165825 -174189 165869 -174181
rect 165925 -174189 165969 -174181
rect 166025 -174189 166069 -174181
rect 166125 -174189 166169 -174181
rect 166225 -174189 166269 -174181
rect 166325 -174189 166369 -174181
rect 166425 -174189 166469 -174181
rect 166525 -174189 166569 -174181
rect 166625 -174189 166669 -174181
rect 166725 -174189 166769 -174181
rect 166825 -174189 166869 -174181
rect 166925 -174189 166969 -174181
rect 167025 -174189 167069 -174181
rect 167525 -174189 167569 -174181
rect 167625 -174189 167669 -174181
rect 167725 -174189 167769 -174181
rect 167825 -174189 167869 -174181
rect 167925 -174189 167969 -174181
rect 168025 -174189 168069 -174181
rect 168125 -174189 168169 -174181
rect 168225 -174189 168269 -174181
rect 168325 -174189 168369 -174181
rect 168425 -174189 168469 -174181
rect 168525 -174189 168569 -174181
rect 168625 -174189 168669 -174181
rect 168725 -174189 168769 -174181
rect 168825 -174189 168869 -174181
rect 168925 -174189 168969 -174181
rect 169025 -174189 169069 -174181
rect 169525 -174189 169569 -174181
rect 169625 -174189 169669 -174181
rect 169725 -174189 169769 -174181
rect 169825 -174189 169869 -174181
rect 169925 -174189 169969 -174181
rect 170025 -174189 170069 -174181
rect 170125 -174189 170169 -174181
rect 170225 -174189 170269 -174181
rect 170325 -174189 170369 -174181
rect 170425 -174189 170469 -174181
rect 170525 -174189 170569 -174181
rect 170625 -174189 170669 -174181
rect 170725 -174189 170769 -174181
rect 170825 -174189 170869 -174181
rect 170925 -174189 170969 -174181
rect 171025 -174189 171069 -174181
rect 171525 -174189 171569 -174181
rect 171625 -174189 171669 -174181
rect 171725 -174189 171769 -174181
rect 171825 -174189 171869 -174181
rect 171925 -174189 171969 -174181
rect 172025 -174189 172069 -174181
rect 172125 -174189 172169 -174181
rect 172225 -174189 172269 -174181
rect 172325 -174189 172369 -174181
rect 172425 -174189 172469 -174181
rect 172525 -174189 172569 -174181
rect 172625 -174189 172669 -174181
rect 172725 -174189 172769 -174181
rect 172825 -174189 172869 -174181
rect 172925 -174189 172969 -174181
rect 173025 -174189 173069 -174181
rect 165569 -174233 165577 -174189
rect 165669 -174233 165677 -174189
rect 165769 -174233 165777 -174189
rect 165869 -174233 165877 -174189
rect 165969 -174233 165977 -174189
rect 166069 -174233 166077 -174189
rect 166169 -174233 166177 -174189
rect 166269 -174233 166277 -174189
rect 166369 -174233 166377 -174189
rect 166469 -174233 166477 -174189
rect 166569 -174233 166577 -174189
rect 166669 -174233 166677 -174189
rect 166769 -174233 166777 -174189
rect 166869 -174233 166877 -174189
rect 166969 -174233 166977 -174189
rect 167069 -174233 167077 -174189
rect 167569 -174233 167577 -174189
rect 167669 -174233 167677 -174189
rect 167769 -174233 167777 -174189
rect 167869 -174233 167877 -174189
rect 167969 -174233 167977 -174189
rect 168069 -174233 168077 -174189
rect 168169 -174233 168177 -174189
rect 168269 -174233 168277 -174189
rect 168369 -174233 168377 -174189
rect 168469 -174233 168477 -174189
rect 168569 -174233 168577 -174189
rect 168669 -174233 168677 -174189
rect 168769 -174233 168777 -174189
rect 168869 -174233 168877 -174189
rect 168969 -174233 168977 -174189
rect 169069 -174233 169077 -174189
rect 169569 -174233 169577 -174189
rect 169669 -174233 169677 -174189
rect 169769 -174233 169777 -174189
rect 169869 -174233 169877 -174189
rect 169969 -174233 169977 -174189
rect 170069 -174233 170077 -174189
rect 170169 -174233 170177 -174189
rect 170269 -174233 170277 -174189
rect 170369 -174233 170377 -174189
rect 170469 -174233 170477 -174189
rect 170569 -174233 170577 -174189
rect 170669 -174233 170677 -174189
rect 170769 -174233 170777 -174189
rect 170869 -174233 170877 -174189
rect 170969 -174233 170977 -174189
rect 171069 -174233 171077 -174189
rect 171569 -174233 171577 -174189
rect 171669 -174233 171677 -174189
rect 171769 -174233 171777 -174189
rect 171869 -174233 171877 -174189
rect 171969 -174233 171977 -174189
rect 172069 -174233 172077 -174189
rect 172169 -174233 172177 -174189
rect 172269 -174233 172277 -174189
rect 172369 -174233 172377 -174189
rect 172469 -174233 172477 -174189
rect 172569 -174233 172577 -174189
rect 172669 -174233 172677 -174189
rect 172769 -174233 172777 -174189
rect 172869 -174233 172877 -174189
rect 172969 -174233 172977 -174189
rect 173069 -174233 173077 -174189
rect 81627 -174249 81671 -174241
rect 81727 -174249 81771 -174241
rect 81827 -174249 81871 -174241
rect 81927 -174249 81971 -174241
rect 82027 -174249 82071 -174241
rect 82127 -174249 82171 -174241
rect 82227 -174249 82271 -174241
rect 82327 -174249 82371 -174241
rect 82427 -174249 82471 -174241
rect 82527 -174249 82571 -174241
rect 82627 -174249 82671 -174241
rect 82727 -174249 82771 -174241
rect 82827 -174249 82871 -174241
rect 82927 -174249 82971 -174241
rect 83027 -174249 83071 -174241
rect 83127 -174249 83171 -174241
rect 83627 -174249 83671 -174241
rect 83727 -174249 83771 -174241
rect 83827 -174249 83871 -174241
rect 83927 -174249 83971 -174241
rect 84027 -174249 84071 -174241
rect 84127 -174249 84171 -174241
rect 84227 -174249 84271 -174241
rect 84327 -174249 84371 -174241
rect 84427 -174249 84471 -174241
rect 84527 -174249 84571 -174241
rect 84627 -174249 84671 -174241
rect 84727 -174249 84771 -174241
rect 84827 -174249 84871 -174241
rect 84927 -174249 84971 -174241
rect 85027 -174249 85071 -174241
rect 85127 -174249 85171 -174241
rect 85627 -174249 85671 -174241
rect 85727 -174249 85771 -174241
rect 85827 -174249 85871 -174241
rect 85927 -174249 85971 -174241
rect 86027 -174249 86071 -174241
rect 86127 -174249 86171 -174241
rect 86227 -174249 86271 -174241
rect 86327 -174249 86371 -174241
rect 86427 -174249 86471 -174241
rect 86527 -174249 86571 -174241
rect 86627 -174249 86671 -174241
rect 86727 -174249 86771 -174241
rect 86827 -174249 86871 -174241
rect 86927 -174249 86971 -174241
rect 87027 -174249 87071 -174241
rect 87127 -174249 87171 -174241
rect 87627 -174249 87671 -174241
rect 87727 -174249 87771 -174241
rect 87827 -174249 87871 -174241
rect 87927 -174249 87971 -174241
rect 88027 -174249 88071 -174241
rect 88127 -174249 88171 -174241
rect 88227 -174249 88271 -174241
rect 88327 -174249 88371 -174241
rect 88427 -174249 88471 -174241
rect 88527 -174249 88571 -174241
rect 88627 -174249 88671 -174241
rect 88727 -174249 88771 -174241
rect 88827 -174249 88871 -174241
rect 88927 -174249 88971 -174241
rect 89027 -174249 89071 -174241
rect 89127 -174249 89171 -174241
rect 81671 -174293 81679 -174249
rect 81771 -174293 81779 -174249
rect 81871 -174293 81879 -174249
rect 81971 -174293 81979 -174249
rect 82071 -174293 82079 -174249
rect 82171 -174293 82179 -174249
rect 82271 -174293 82279 -174249
rect 82371 -174293 82379 -174249
rect 82471 -174293 82479 -174249
rect 82571 -174293 82579 -174249
rect 82671 -174293 82679 -174249
rect 82771 -174293 82779 -174249
rect 82871 -174293 82879 -174249
rect 82971 -174293 82979 -174249
rect 83071 -174293 83079 -174249
rect 83171 -174293 83179 -174249
rect 83671 -174293 83679 -174249
rect 83771 -174293 83779 -174249
rect 83871 -174293 83879 -174249
rect 83971 -174293 83979 -174249
rect 84071 -174293 84079 -174249
rect 84171 -174293 84179 -174249
rect 84271 -174293 84279 -174249
rect 84371 -174293 84379 -174249
rect 84471 -174293 84479 -174249
rect 84571 -174293 84579 -174249
rect 84671 -174293 84679 -174249
rect 84771 -174293 84779 -174249
rect 84871 -174293 84879 -174249
rect 84971 -174293 84979 -174249
rect 85071 -174293 85079 -174249
rect 85171 -174293 85179 -174249
rect 85671 -174293 85679 -174249
rect 85771 -174293 85779 -174249
rect 85871 -174293 85879 -174249
rect 85971 -174293 85979 -174249
rect 86071 -174293 86079 -174249
rect 86171 -174293 86179 -174249
rect 86271 -174293 86279 -174249
rect 86371 -174293 86379 -174249
rect 86471 -174293 86479 -174249
rect 86571 -174293 86579 -174249
rect 86671 -174293 86679 -174249
rect 86771 -174293 86779 -174249
rect 86871 -174293 86879 -174249
rect 86971 -174293 86979 -174249
rect 87071 -174293 87079 -174249
rect 87171 -174293 87179 -174249
rect 87671 -174293 87679 -174249
rect 87771 -174293 87779 -174249
rect 87871 -174293 87879 -174249
rect 87971 -174293 87979 -174249
rect 88071 -174293 88079 -174249
rect 88171 -174293 88179 -174249
rect 88271 -174293 88279 -174249
rect 88371 -174293 88379 -174249
rect 88471 -174293 88479 -174249
rect 88571 -174293 88579 -174249
rect 88671 -174293 88679 -174249
rect 88771 -174293 88779 -174249
rect 88871 -174293 88879 -174249
rect 88971 -174293 88979 -174249
rect 89071 -174293 89079 -174249
rect 89171 -174293 89179 -174249
rect 165525 -174289 165569 -174281
rect 165625 -174289 165669 -174281
rect 165725 -174289 165769 -174281
rect 165825 -174289 165869 -174281
rect 165925 -174289 165969 -174281
rect 166025 -174289 166069 -174281
rect 166125 -174289 166169 -174281
rect 166225 -174289 166269 -174281
rect 166325 -174289 166369 -174281
rect 166425 -174289 166469 -174281
rect 166525 -174289 166569 -174281
rect 166625 -174289 166669 -174281
rect 166725 -174289 166769 -174281
rect 166825 -174289 166869 -174281
rect 166925 -174289 166969 -174281
rect 167025 -174289 167069 -174281
rect 167525 -174289 167569 -174281
rect 167625 -174289 167669 -174281
rect 167725 -174289 167769 -174281
rect 167825 -174289 167869 -174281
rect 167925 -174289 167969 -174281
rect 168025 -174289 168069 -174281
rect 168125 -174289 168169 -174281
rect 168225 -174289 168269 -174281
rect 168325 -174289 168369 -174281
rect 168425 -174289 168469 -174281
rect 168525 -174289 168569 -174281
rect 168625 -174289 168669 -174281
rect 168725 -174289 168769 -174281
rect 168825 -174289 168869 -174281
rect 168925 -174289 168969 -174281
rect 169025 -174289 169069 -174281
rect 169525 -174289 169569 -174281
rect 169625 -174289 169669 -174281
rect 169725 -174289 169769 -174281
rect 169825 -174289 169869 -174281
rect 169925 -174289 169969 -174281
rect 170025 -174289 170069 -174281
rect 170125 -174289 170169 -174281
rect 170225 -174289 170269 -174281
rect 170325 -174289 170369 -174281
rect 170425 -174289 170469 -174281
rect 170525 -174289 170569 -174281
rect 170625 -174289 170669 -174281
rect 170725 -174289 170769 -174281
rect 170825 -174289 170869 -174281
rect 170925 -174289 170969 -174281
rect 171025 -174289 171069 -174281
rect 171525 -174289 171569 -174281
rect 171625 -174289 171669 -174281
rect 171725 -174289 171769 -174281
rect 171825 -174289 171869 -174281
rect 171925 -174289 171969 -174281
rect 172025 -174289 172069 -174281
rect 172125 -174289 172169 -174281
rect 172225 -174289 172269 -174281
rect 172325 -174289 172369 -174281
rect 172425 -174289 172469 -174281
rect 172525 -174289 172569 -174281
rect 172625 -174289 172669 -174281
rect 172725 -174289 172769 -174281
rect 172825 -174289 172869 -174281
rect 172925 -174289 172969 -174281
rect 173025 -174289 173069 -174281
rect 165569 -174333 165577 -174289
rect 165669 -174333 165677 -174289
rect 165769 -174333 165777 -174289
rect 165869 -174333 165877 -174289
rect 165969 -174333 165977 -174289
rect 166069 -174333 166077 -174289
rect 166169 -174333 166177 -174289
rect 166269 -174333 166277 -174289
rect 166369 -174333 166377 -174289
rect 166469 -174333 166477 -174289
rect 166569 -174333 166577 -174289
rect 166669 -174333 166677 -174289
rect 166769 -174333 166777 -174289
rect 166869 -174333 166877 -174289
rect 166969 -174333 166977 -174289
rect 167069 -174333 167077 -174289
rect 167569 -174333 167577 -174289
rect 167669 -174333 167677 -174289
rect 167769 -174333 167777 -174289
rect 167869 -174333 167877 -174289
rect 167969 -174333 167977 -174289
rect 168069 -174333 168077 -174289
rect 168169 -174333 168177 -174289
rect 168269 -174333 168277 -174289
rect 168369 -174333 168377 -174289
rect 168469 -174333 168477 -174289
rect 168569 -174333 168577 -174289
rect 168669 -174333 168677 -174289
rect 168769 -174333 168777 -174289
rect 168869 -174333 168877 -174289
rect 168969 -174333 168977 -174289
rect 169069 -174333 169077 -174289
rect 169569 -174333 169577 -174289
rect 169669 -174333 169677 -174289
rect 169769 -174333 169777 -174289
rect 169869 -174333 169877 -174289
rect 169969 -174333 169977 -174289
rect 170069 -174333 170077 -174289
rect 170169 -174333 170177 -174289
rect 170269 -174333 170277 -174289
rect 170369 -174333 170377 -174289
rect 170469 -174333 170477 -174289
rect 170569 -174333 170577 -174289
rect 170669 -174333 170677 -174289
rect 170769 -174333 170777 -174289
rect 170869 -174333 170877 -174289
rect 170969 -174333 170977 -174289
rect 171069 -174333 171077 -174289
rect 171569 -174333 171577 -174289
rect 171669 -174333 171677 -174289
rect 171769 -174333 171777 -174289
rect 171869 -174333 171877 -174289
rect 171969 -174333 171977 -174289
rect 172069 -174333 172077 -174289
rect 172169 -174333 172177 -174289
rect 172269 -174333 172277 -174289
rect 172369 -174333 172377 -174289
rect 172469 -174333 172477 -174289
rect 172569 -174333 172577 -174289
rect 172669 -174333 172677 -174289
rect 172769 -174333 172777 -174289
rect 172869 -174333 172877 -174289
rect 172969 -174333 172977 -174289
rect 173069 -174333 173077 -174289
rect 81627 -174349 81671 -174341
rect 81727 -174349 81771 -174341
rect 81827 -174349 81871 -174341
rect 81927 -174349 81971 -174341
rect 82027 -174349 82071 -174341
rect 82127 -174349 82171 -174341
rect 82227 -174349 82271 -174341
rect 82327 -174349 82371 -174341
rect 82427 -174349 82471 -174341
rect 82527 -174349 82571 -174341
rect 82627 -174349 82671 -174341
rect 82727 -174349 82771 -174341
rect 82827 -174349 82871 -174341
rect 82927 -174349 82971 -174341
rect 83027 -174349 83071 -174341
rect 83127 -174349 83171 -174341
rect 83627 -174349 83671 -174341
rect 83727 -174349 83771 -174341
rect 83827 -174349 83871 -174341
rect 83927 -174349 83971 -174341
rect 84027 -174349 84071 -174341
rect 84127 -174349 84171 -174341
rect 84227 -174349 84271 -174341
rect 84327 -174349 84371 -174341
rect 84427 -174349 84471 -174341
rect 84527 -174349 84571 -174341
rect 84627 -174349 84671 -174341
rect 84727 -174349 84771 -174341
rect 84827 -174349 84871 -174341
rect 84927 -174349 84971 -174341
rect 85027 -174349 85071 -174341
rect 85127 -174349 85171 -174341
rect 85627 -174349 85671 -174341
rect 85727 -174349 85771 -174341
rect 85827 -174349 85871 -174341
rect 85927 -174349 85971 -174341
rect 86027 -174349 86071 -174341
rect 86127 -174349 86171 -174341
rect 86227 -174349 86271 -174341
rect 86327 -174349 86371 -174341
rect 86427 -174349 86471 -174341
rect 86527 -174349 86571 -174341
rect 86627 -174349 86671 -174341
rect 86727 -174349 86771 -174341
rect 86827 -174349 86871 -174341
rect 86927 -174349 86971 -174341
rect 87027 -174349 87071 -174341
rect 87127 -174349 87171 -174341
rect 87627 -174349 87671 -174341
rect 87727 -174349 87771 -174341
rect 87827 -174349 87871 -174341
rect 87927 -174349 87971 -174341
rect 88027 -174349 88071 -174341
rect 88127 -174349 88171 -174341
rect 88227 -174349 88271 -174341
rect 88327 -174349 88371 -174341
rect 88427 -174349 88471 -174341
rect 88527 -174349 88571 -174341
rect 88627 -174349 88671 -174341
rect 88727 -174349 88771 -174341
rect 88827 -174349 88871 -174341
rect 88927 -174349 88971 -174341
rect 89027 -174349 89071 -174341
rect 89127 -174349 89171 -174341
rect 81671 -174393 81679 -174349
rect 81771 -174393 81779 -174349
rect 81871 -174393 81879 -174349
rect 81971 -174393 81979 -174349
rect 82071 -174393 82079 -174349
rect 82171 -174393 82179 -174349
rect 82271 -174393 82279 -174349
rect 82371 -174393 82379 -174349
rect 82471 -174393 82479 -174349
rect 82571 -174393 82579 -174349
rect 82671 -174393 82679 -174349
rect 82771 -174393 82779 -174349
rect 82871 -174393 82879 -174349
rect 82971 -174393 82979 -174349
rect 83071 -174393 83079 -174349
rect 83171 -174393 83179 -174349
rect 83671 -174393 83679 -174349
rect 83771 -174393 83779 -174349
rect 83871 -174393 83879 -174349
rect 83971 -174393 83979 -174349
rect 84071 -174393 84079 -174349
rect 84171 -174393 84179 -174349
rect 84271 -174393 84279 -174349
rect 84371 -174393 84379 -174349
rect 84471 -174393 84479 -174349
rect 84571 -174393 84579 -174349
rect 84671 -174393 84679 -174349
rect 84771 -174393 84779 -174349
rect 84871 -174393 84879 -174349
rect 84971 -174393 84979 -174349
rect 85071 -174393 85079 -174349
rect 85171 -174393 85179 -174349
rect 85671 -174393 85679 -174349
rect 85771 -174393 85779 -174349
rect 85871 -174393 85879 -174349
rect 85971 -174393 85979 -174349
rect 86071 -174393 86079 -174349
rect 86171 -174393 86179 -174349
rect 86271 -174393 86279 -174349
rect 86371 -174393 86379 -174349
rect 86471 -174393 86479 -174349
rect 86571 -174393 86579 -174349
rect 86671 -174393 86679 -174349
rect 86771 -174393 86779 -174349
rect 86871 -174393 86879 -174349
rect 86971 -174393 86979 -174349
rect 87071 -174393 87079 -174349
rect 87171 -174393 87179 -174349
rect 87671 -174393 87679 -174349
rect 87771 -174393 87779 -174349
rect 87871 -174393 87879 -174349
rect 87971 -174393 87979 -174349
rect 88071 -174393 88079 -174349
rect 88171 -174393 88179 -174349
rect 88271 -174393 88279 -174349
rect 88371 -174393 88379 -174349
rect 88471 -174393 88479 -174349
rect 88571 -174393 88579 -174349
rect 88671 -174393 88679 -174349
rect 88771 -174393 88779 -174349
rect 88871 -174393 88879 -174349
rect 88971 -174393 88979 -174349
rect 89071 -174393 89079 -174349
rect 89171 -174393 89179 -174349
rect 165525 -174389 165569 -174381
rect 165625 -174389 165669 -174381
rect 165725 -174389 165769 -174381
rect 165825 -174389 165869 -174381
rect 165925 -174389 165969 -174381
rect 166025 -174389 166069 -174381
rect 166125 -174389 166169 -174381
rect 166225 -174389 166269 -174381
rect 166325 -174389 166369 -174381
rect 166425 -174389 166469 -174381
rect 166525 -174389 166569 -174381
rect 166625 -174389 166669 -174381
rect 166725 -174389 166769 -174381
rect 166825 -174389 166869 -174381
rect 166925 -174389 166969 -174381
rect 167025 -174389 167069 -174381
rect 167525 -174389 167569 -174381
rect 167625 -174389 167669 -174381
rect 167725 -174389 167769 -174381
rect 167825 -174389 167869 -174381
rect 167925 -174389 167969 -174381
rect 168025 -174389 168069 -174381
rect 168125 -174389 168169 -174381
rect 168225 -174389 168269 -174381
rect 168325 -174389 168369 -174381
rect 168425 -174389 168469 -174381
rect 168525 -174389 168569 -174381
rect 168625 -174389 168669 -174381
rect 168725 -174389 168769 -174381
rect 168825 -174389 168869 -174381
rect 168925 -174389 168969 -174381
rect 169025 -174389 169069 -174381
rect 169525 -174389 169569 -174381
rect 169625 -174389 169669 -174381
rect 169725 -174389 169769 -174381
rect 169825 -174389 169869 -174381
rect 169925 -174389 169969 -174381
rect 170025 -174389 170069 -174381
rect 170125 -174389 170169 -174381
rect 170225 -174389 170269 -174381
rect 170325 -174389 170369 -174381
rect 170425 -174389 170469 -174381
rect 170525 -174389 170569 -174381
rect 170625 -174389 170669 -174381
rect 170725 -174389 170769 -174381
rect 170825 -174389 170869 -174381
rect 170925 -174389 170969 -174381
rect 171025 -174389 171069 -174381
rect 171525 -174389 171569 -174381
rect 171625 -174389 171669 -174381
rect 171725 -174389 171769 -174381
rect 171825 -174389 171869 -174381
rect 171925 -174389 171969 -174381
rect 172025 -174389 172069 -174381
rect 172125 -174389 172169 -174381
rect 172225 -174389 172269 -174381
rect 172325 -174389 172369 -174381
rect 172425 -174389 172469 -174381
rect 172525 -174389 172569 -174381
rect 172625 -174389 172669 -174381
rect 172725 -174389 172769 -174381
rect 172825 -174389 172869 -174381
rect 172925 -174389 172969 -174381
rect 173025 -174389 173069 -174381
rect 165569 -174433 165577 -174389
rect 165669 -174433 165677 -174389
rect 165769 -174433 165777 -174389
rect 165869 -174433 165877 -174389
rect 165969 -174433 165977 -174389
rect 166069 -174433 166077 -174389
rect 166169 -174433 166177 -174389
rect 166269 -174433 166277 -174389
rect 166369 -174433 166377 -174389
rect 166469 -174433 166477 -174389
rect 166569 -174433 166577 -174389
rect 166669 -174433 166677 -174389
rect 166769 -174433 166777 -174389
rect 166869 -174433 166877 -174389
rect 166969 -174433 166977 -174389
rect 167069 -174433 167077 -174389
rect 167569 -174433 167577 -174389
rect 167669 -174433 167677 -174389
rect 167769 -174433 167777 -174389
rect 167869 -174433 167877 -174389
rect 167969 -174433 167977 -174389
rect 168069 -174433 168077 -174389
rect 168169 -174433 168177 -174389
rect 168269 -174433 168277 -174389
rect 168369 -174433 168377 -174389
rect 168469 -174433 168477 -174389
rect 168569 -174433 168577 -174389
rect 168669 -174433 168677 -174389
rect 168769 -174433 168777 -174389
rect 168869 -174433 168877 -174389
rect 168969 -174433 168977 -174389
rect 169069 -174433 169077 -174389
rect 169569 -174433 169577 -174389
rect 169669 -174433 169677 -174389
rect 169769 -174433 169777 -174389
rect 169869 -174433 169877 -174389
rect 169969 -174433 169977 -174389
rect 170069 -174433 170077 -174389
rect 170169 -174433 170177 -174389
rect 170269 -174433 170277 -174389
rect 170369 -174433 170377 -174389
rect 170469 -174433 170477 -174389
rect 170569 -174433 170577 -174389
rect 170669 -174433 170677 -174389
rect 170769 -174433 170777 -174389
rect 170869 -174433 170877 -174389
rect 170969 -174433 170977 -174389
rect 171069 -174433 171077 -174389
rect 171569 -174433 171577 -174389
rect 171669 -174433 171677 -174389
rect 171769 -174433 171777 -174389
rect 171869 -174433 171877 -174389
rect 171969 -174433 171977 -174389
rect 172069 -174433 172077 -174389
rect 172169 -174433 172177 -174389
rect 172269 -174433 172277 -174389
rect 172369 -174433 172377 -174389
rect 172469 -174433 172477 -174389
rect 172569 -174433 172577 -174389
rect 172669 -174433 172677 -174389
rect 172769 -174433 172777 -174389
rect 172869 -174433 172877 -174389
rect 172969 -174433 172977 -174389
rect 173069 -174433 173077 -174389
rect 81627 -174449 81671 -174441
rect 81727 -174449 81771 -174441
rect 81827 -174449 81871 -174441
rect 81927 -174449 81971 -174441
rect 82027 -174449 82071 -174441
rect 82127 -174449 82171 -174441
rect 82227 -174449 82271 -174441
rect 82327 -174449 82371 -174441
rect 82427 -174449 82471 -174441
rect 82527 -174449 82571 -174441
rect 82627 -174449 82671 -174441
rect 82727 -174449 82771 -174441
rect 82827 -174449 82871 -174441
rect 82927 -174449 82971 -174441
rect 83027 -174449 83071 -174441
rect 83127 -174449 83171 -174441
rect 83627 -174449 83671 -174441
rect 83727 -174449 83771 -174441
rect 83827 -174449 83871 -174441
rect 83927 -174449 83971 -174441
rect 84027 -174449 84071 -174441
rect 84127 -174449 84171 -174441
rect 84227 -174449 84271 -174441
rect 84327 -174449 84371 -174441
rect 84427 -174449 84471 -174441
rect 84527 -174449 84571 -174441
rect 84627 -174449 84671 -174441
rect 84727 -174449 84771 -174441
rect 84827 -174449 84871 -174441
rect 84927 -174449 84971 -174441
rect 85027 -174449 85071 -174441
rect 85127 -174449 85171 -174441
rect 85627 -174449 85671 -174441
rect 85727 -174449 85771 -174441
rect 85827 -174449 85871 -174441
rect 85927 -174449 85971 -174441
rect 86027 -174449 86071 -174441
rect 86127 -174449 86171 -174441
rect 86227 -174449 86271 -174441
rect 86327 -174449 86371 -174441
rect 86427 -174449 86471 -174441
rect 86527 -174449 86571 -174441
rect 86627 -174449 86671 -174441
rect 86727 -174449 86771 -174441
rect 86827 -174449 86871 -174441
rect 86927 -174449 86971 -174441
rect 87027 -174449 87071 -174441
rect 87127 -174449 87171 -174441
rect 87627 -174449 87671 -174441
rect 87727 -174449 87771 -174441
rect 87827 -174449 87871 -174441
rect 87927 -174449 87971 -174441
rect 88027 -174449 88071 -174441
rect 88127 -174449 88171 -174441
rect 88227 -174449 88271 -174441
rect 88327 -174449 88371 -174441
rect 88427 -174449 88471 -174441
rect 88527 -174449 88571 -174441
rect 88627 -174449 88671 -174441
rect 88727 -174449 88771 -174441
rect 88827 -174449 88871 -174441
rect 88927 -174449 88971 -174441
rect 89027 -174449 89071 -174441
rect 89127 -174449 89171 -174441
rect 81671 -174493 81679 -174449
rect 81771 -174493 81779 -174449
rect 81871 -174493 81879 -174449
rect 81971 -174493 81979 -174449
rect 82071 -174493 82079 -174449
rect 82171 -174493 82179 -174449
rect 82271 -174493 82279 -174449
rect 82371 -174493 82379 -174449
rect 82471 -174493 82479 -174449
rect 82571 -174493 82579 -174449
rect 82671 -174493 82679 -174449
rect 82771 -174493 82779 -174449
rect 82871 -174493 82879 -174449
rect 82971 -174493 82979 -174449
rect 83071 -174493 83079 -174449
rect 83171 -174493 83179 -174449
rect 83671 -174493 83679 -174449
rect 83771 -174493 83779 -174449
rect 83871 -174493 83879 -174449
rect 83971 -174493 83979 -174449
rect 84071 -174493 84079 -174449
rect 84171 -174493 84179 -174449
rect 84271 -174493 84279 -174449
rect 84371 -174493 84379 -174449
rect 84471 -174493 84479 -174449
rect 84571 -174493 84579 -174449
rect 84671 -174493 84679 -174449
rect 84771 -174493 84779 -174449
rect 84871 -174493 84879 -174449
rect 84971 -174493 84979 -174449
rect 85071 -174493 85079 -174449
rect 85171 -174493 85179 -174449
rect 85671 -174493 85679 -174449
rect 85771 -174493 85779 -174449
rect 85871 -174493 85879 -174449
rect 85971 -174493 85979 -174449
rect 86071 -174493 86079 -174449
rect 86171 -174493 86179 -174449
rect 86271 -174493 86279 -174449
rect 86371 -174493 86379 -174449
rect 86471 -174493 86479 -174449
rect 86571 -174493 86579 -174449
rect 86671 -174493 86679 -174449
rect 86771 -174493 86779 -174449
rect 86871 -174493 86879 -174449
rect 86971 -174493 86979 -174449
rect 87071 -174493 87079 -174449
rect 87171 -174493 87179 -174449
rect 87671 -174493 87679 -174449
rect 87771 -174493 87779 -174449
rect 87871 -174493 87879 -174449
rect 87971 -174493 87979 -174449
rect 88071 -174493 88079 -174449
rect 88171 -174493 88179 -174449
rect 88271 -174493 88279 -174449
rect 88371 -174493 88379 -174449
rect 88471 -174493 88479 -174449
rect 88571 -174493 88579 -174449
rect 88671 -174493 88679 -174449
rect 88771 -174493 88779 -174449
rect 88871 -174493 88879 -174449
rect 88971 -174493 88979 -174449
rect 89071 -174493 89079 -174449
rect 89171 -174493 89179 -174449
rect 165525 -174489 165569 -174481
rect 165625 -174489 165669 -174481
rect 165725 -174489 165769 -174481
rect 165825 -174489 165869 -174481
rect 165925 -174489 165969 -174481
rect 166025 -174489 166069 -174481
rect 166125 -174489 166169 -174481
rect 166225 -174489 166269 -174481
rect 166325 -174489 166369 -174481
rect 166425 -174489 166469 -174481
rect 166525 -174489 166569 -174481
rect 166625 -174489 166669 -174481
rect 166725 -174489 166769 -174481
rect 166825 -174489 166869 -174481
rect 166925 -174489 166969 -174481
rect 167025 -174489 167069 -174481
rect 167525 -174489 167569 -174481
rect 167625 -174489 167669 -174481
rect 167725 -174489 167769 -174481
rect 167825 -174489 167869 -174481
rect 167925 -174489 167969 -174481
rect 168025 -174489 168069 -174481
rect 168125 -174489 168169 -174481
rect 168225 -174489 168269 -174481
rect 168325 -174489 168369 -174481
rect 168425 -174489 168469 -174481
rect 168525 -174489 168569 -174481
rect 168625 -174489 168669 -174481
rect 168725 -174489 168769 -174481
rect 168825 -174489 168869 -174481
rect 168925 -174489 168969 -174481
rect 169025 -174489 169069 -174481
rect 169525 -174489 169569 -174481
rect 169625 -174489 169669 -174481
rect 169725 -174489 169769 -174481
rect 169825 -174489 169869 -174481
rect 169925 -174489 169969 -174481
rect 170025 -174489 170069 -174481
rect 170125 -174489 170169 -174481
rect 170225 -174489 170269 -174481
rect 170325 -174489 170369 -174481
rect 170425 -174489 170469 -174481
rect 170525 -174489 170569 -174481
rect 170625 -174489 170669 -174481
rect 170725 -174489 170769 -174481
rect 170825 -174489 170869 -174481
rect 170925 -174489 170969 -174481
rect 171025 -174489 171069 -174481
rect 171525 -174489 171569 -174481
rect 171625 -174489 171669 -174481
rect 171725 -174489 171769 -174481
rect 171825 -174489 171869 -174481
rect 171925 -174489 171969 -174481
rect 172025 -174489 172069 -174481
rect 172125 -174489 172169 -174481
rect 172225 -174489 172269 -174481
rect 172325 -174489 172369 -174481
rect 172425 -174489 172469 -174481
rect 172525 -174489 172569 -174481
rect 172625 -174489 172669 -174481
rect 172725 -174489 172769 -174481
rect 172825 -174489 172869 -174481
rect 172925 -174489 172969 -174481
rect 173025 -174489 173069 -174481
rect 165569 -174533 165577 -174489
rect 165669 -174533 165677 -174489
rect 165769 -174533 165777 -174489
rect 165869 -174533 165877 -174489
rect 165969 -174533 165977 -174489
rect 166069 -174533 166077 -174489
rect 166169 -174533 166177 -174489
rect 166269 -174533 166277 -174489
rect 166369 -174533 166377 -174489
rect 166469 -174533 166477 -174489
rect 166569 -174533 166577 -174489
rect 166669 -174533 166677 -174489
rect 166769 -174533 166777 -174489
rect 166869 -174533 166877 -174489
rect 166969 -174533 166977 -174489
rect 167069 -174533 167077 -174489
rect 167569 -174533 167577 -174489
rect 167669 -174533 167677 -174489
rect 167769 -174533 167777 -174489
rect 167869 -174533 167877 -174489
rect 167969 -174533 167977 -174489
rect 168069 -174533 168077 -174489
rect 168169 -174533 168177 -174489
rect 168269 -174533 168277 -174489
rect 168369 -174533 168377 -174489
rect 168469 -174533 168477 -174489
rect 168569 -174533 168577 -174489
rect 168669 -174533 168677 -174489
rect 168769 -174533 168777 -174489
rect 168869 -174533 168877 -174489
rect 168969 -174533 168977 -174489
rect 169069 -174533 169077 -174489
rect 169569 -174533 169577 -174489
rect 169669 -174533 169677 -174489
rect 169769 -174533 169777 -174489
rect 169869 -174533 169877 -174489
rect 169969 -174533 169977 -174489
rect 170069 -174533 170077 -174489
rect 170169 -174533 170177 -174489
rect 170269 -174533 170277 -174489
rect 170369 -174533 170377 -174489
rect 170469 -174533 170477 -174489
rect 170569 -174533 170577 -174489
rect 170669 -174533 170677 -174489
rect 170769 -174533 170777 -174489
rect 170869 -174533 170877 -174489
rect 170969 -174533 170977 -174489
rect 171069 -174533 171077 -174489
rect 171569 -174533 171577 -174489
rect 171669 -174533 171677 -174489
rect 171769 -174533 171777 -174489
rect 171869 -174533 171877 -174489
rect 171969 -174533 171977 -174489
rect 172069 -174533 172077 -174489
rect 172169 -174533 172177 -174489
rect 172269 -174533 172277 -174489
rect 172369 -174533 172377 -174489
rect 172469 -174533 172477 -174489
rect 172569 -174533 172577 -174489
rect 172669 -174533 172677 -174489
rect 172769 -174533 172777 -174489
rect 172869 -174533 172877 -174489
rect 172969 -174533 172977 -174489
rect 173069 -174533 173077 -174489
rect 81627 -174549 81671 -174541
rect 81727 -174549 81771 -174541
rect 81827 -174549 81871 -174541
rect 81927 -174549 81971 -174541
rect 82027 -174549 82071 -174541
rect 82127 -174549 82171 -174541
rect 82227 -174549 82271 -174541
rect 82327 -174549 82371 -174541
rect 82427 -174549 82471 -174541
rect 82527 -174549 82571 -174541
rect 82627 -174549 82671 -174541
rect 82727 -174549 82771 -174541
rect 82827 -174549 82871 -174541
rect 82927 -174549 82971 -174541
rect 83027 -174549 83071 -174541
rect 83127 -174549 83171 -174541
rect 83627 -174549 83671 -174541
rect 83727 -174549 83771 -174541
rect 83827 -174549 83871 -174541
rect 83927 -174549 83971 -174541
rect 84027 -174549 84071 -174541
rect 84127 -174549 84171 -174541
rect 84227 -174549 84271 -174541
rect 84327 -174549 84371 -174541
rect 84427 -174549 84471 -174541
rect 84527 -174549 84571 -174541
rect 84627 -174549 84671 -174541
rect 84727 -174549 84771 -174541
rect 84827 -174549 84871 -174541
rect 84927 -174549 84971 -174541
rect 85027 -174549 85071 -174541
rect 85127 -174549 85171 -174541
rect 85627 -174549 85671 -174541
rect 85727 -174549 85771 -174541
rect 85827 -174549 85871 -174541
rect 85927 -174549 85971 -174541
rect 86027 -174549 86071 -174541
rect 86127 -174549 86171 -174541
rect 86227 -174549 86271 -174541
rect 86327 -174549 86371 -174541
rect 86427 -174549 86471 -174541
rect 86527 -174549 86571 -174541
rect 86627 -174549 86671 -174541
rect 86727 -174549 86771 -174541
rect 86827 -174549 86871 -174541
rect 86927 -174549 86971 -174541
rect 87027 -174549 87071 -174541
rect 87127 -174549 87171 -174541
rect 87627 -174549 87671 -174541
rect 87727 -174549 87771 -174541
rect 87827 -174549 87871 -174541
rect 87927 -174549 87971 -174541
rect 88027 -174549 88071 -174541
rect 88127 -174549 88171 -174541
rect 88227 -174549 88271 -174541
rect 88327 -174549 88371 -174541
rect 88427 -174549 88471 -174541
rect 88527 -174549 88571 -174541
rect 88627 -174549 88671 -174541
rect 88727 -174549 88771 -174541
rect 88827 -174549 88871 -174541
rect 88927 -174549 88971 -174541
rect 89027 -174549 89071 -174541
rect 89127 -174549 89171 -174541
rect 81671 -174593 81679 -174549
rect 81771 -174593 81779 -174549
rect 81871 -174593 81879 -174549
rect 81971 -174593 81979 -174549
rect 82071 -174593 82079 -174549
rect 82171 -174593 82179 -174549
rect 82271 -174593 82279 -174549
rect 82371 -174593 82379 -174549
rect 82471 -174593 82479 -174549
rect 82571 -174593 82579 -174549
rect 82671 -174593 82679 -174549
rect 82771 -174593 82779 -174549
rect 82871 -174593 82879 -174549
rect 82971 -174593 82979 -174549
rect 83071 -174593 83079 -174549
rect 83171 -174593 83179 -174549
rect 83671 -174593 83679 -174549
rect 83771 -174593 83779 -174549
rect 83871 -174593 83879 -174549
rect 83971 -174593 83979 -174549
rect 84071 -174593 84079 -174549
rect 84171 -174593 84179 -174549
rect 84271 -174593 84279 -174549
rect 84371 -174593 84379 -174549
rect 84471 -174593 84479 -174549
rect 84571 -174593 84579 -174549
rect 84671 -174593 84679 -174549
rect 84771 -174593 84779 -174549
rect 84871 -174593 84879 -174549
rect 84971 -174593 84979 -174549
rect 85071 -174593 85079 -174549
rect 85171 -174593 85179 -174549
rect 85671 -174593 85679 -174549
rect 85771 -174593 85779 -174549
rect 85871 -174593 85879 -174549
rect 85971 -174593 85979 -174549
rect 86071 -174593 86079 -174549
rect 86171 -174593 86179 -174549
rect 86271 -174593 86279 -174549
rect 86371 -174593 86379 -174549
rect 86471 -174593 86479 -174549
rect 86571 -174593 86579 -174549
rect 86671 -174593 86679 -174549
rect 86771 -174593 86779 -174549
rect 86871 -174593 86879 -174549
rect 86971 -174593 86979 -174549
rect 87071 -174593 87079 -174549
rect 87171 -174593 87179 -174549
rect 87671 -174593 87679 -174549
rect 87771 -174593 87779 -174549
rect 87871 -174593 87879 -174549
rect 87971 -174593 87979 -174549
rect 88071 -174593 88079 -174549
rect 88171 -174593 88179 -174549
rect 88271 -174593 88279 -174549
rect 88371 -174593 88379 -174549
rect 88471 -174593 88479 -174549
rect 88571 -174593 88579 -174549
rect 88671 -174593 88679 -174549
rect 88771 -174593 88779 -174549
rect 88871 -174593 88879 -174549
rect 88971 -174593 88979 -174549
rect 89071 -174593 89079 -174549
rect 89171 -174593 89179 -174549
<< error_s >>
rect -6848 4066 -6846 6066
rect -6782 4066 -6780 6066
rect -172 -46 -170 9954
rect -106 -46 -104 9954
rect 27828 -46 27830 9954
rect 27894 -46 27896 9954
rect 57950 5307 57952 25307
rect 58016 5307 58018 25307
rect 84950 5307 84952 25307
rect 85016 5307 85018 25307
rect 37223 -9638 37267 -9630
rect 37323 -9638 37367 -9630
rect 37423 -9638 37467 -9630
rect 37523 -9638 37567 -9630
rect 37623 -9638 37667 -9630
rect 37723 -9638 37767 -9630
rect 37823 -9638 37867 -9630
rect 37923 -9638 37967 -9630
rect 38023 -9638 38067 -9630
rect 38123 -9638 38167 -9630
rect 38223 -9638 38267 -9630
rect 38323 -9638 38367 -9630
rect 38423 -9638 38467 -9630
rect 38523 -9638 38567 -9630
rect 38623 -9638 38667 -9630
rect 38723 -9638 38767 -9630
rect 39223 -9638 39267 -9630
rect 39323 -9638 39367 -9630
rect 39423 -9638 39467 -9630
rect 39523 -9638 39567 -9630
rect 39623 -9638 39667 -9630
rect 39723 -9638 39767 -9630
rect 39823 -9638 39867 -9630
rect 39923 -9638 39967 -9630
rect 40023 -9638 40067 -9630
rect 40123 -9638 40167 -9630
rect 40223 -9638 40267 -9630
rect 40323 -9638 40367 -9630
rect 40423 -9638 40467 -9630
rect 40523 -9638 40567 -9630
rect 40623 -9638 40667 -9630
rect 40723 -9638 40767 -9630
rect 41223 -9638 41267 -9630
rect 41323 -9638 41367 -9630
rect 41423 -9638 41467 -9630
rect 41523 -9638 41567 -9630
rect 41623 -9638 41667 -9630
rect 41723 -9638 41767 -9630
rect 41823 -9638 41867 -9630
rect 41923 -9638 41967 -9630
rect 42023 -9638 42067 -9630
rect 42123 -9638 42167 -9630
rect 42223 -9638 42267 -9630
rect 42323 -9638 42367 -9630
rect 42423 -9638 42467 -9630
rect 42523 -9638 42567 -9630
rect 42623 -9638 42667 -9630
rect 42723 -9638 42767 -9630
rect 43223 -9638 43267 -9630
rect 43323 -9638 43367 -9630
rect 43423 -9638 43467 -9630
rect 43523 -9638 43567 -9630
rect 43623 -9638 43667 -9630
rect 43723 -9638 43767 -9630
rect 43823 -9638 43867 -9630
rect 43923 -9638 43967 -9630
rect 44023 -9638 44067 -9630
rect 44123 -9638 44167 -9630
rect 44223 -9638 44267 -9630
rect 44323 -9638 44367 -9630
rect 44423 -9638 44467 -9630
rect 44523 -9638 44567 -9630
rect 44623 -9638 44667 -9630
rect 44723 -9638 44767 -9630
rect 37267 -9682 37275 -9638
rect 37367 -9682 37375 -9638
rect 37467 -9682 37475 -9638
rect 37567 -9682 37575 -9638
rect 37667 -9682 37675 -9638
rect 37767 -9682 37775 -9638
rect 37867 -9682 37875 -9638
rect 37967 -9682 37975 -9638
rect 38067 -9682 38075 -9638
rect 38167 -9682 38175 -9638
rect 38267 -9682 38275 -9638
rect 38367 -9682 38375 -9638
rect 38467 -9682 38475 -9638
rect 38567 -9682 38575 -9638
rect 38667 -9682 38675 -9638
rect 38767 -9682 38775 -9638
rect 39267 -9682 39275 -9638
rect 39367 -9682 39375 -9638
rect 39467 -9682 39475 -9638
rect 39567 -9682 39575 -9638
rect 39667 -9682 39675 -9638
rect 39767 -9682 39775 -9638
rect 39867 -9682 39875 -9638
rect 39967 -9682 39975 -9638
rect 40067 -9682 40075 -9638
rect 40167 -9682 40175 -9638
rect 40267 -9682 40275 -9638
rect 40367 -9682 40375 -9638
rect 40467 -9682 40475 -9638
rect 40567 -9682 40575 -9638
rect 40667 -9682 40675 -9638
rect 40767 -9682 40775 -9638
rect 41267 -9682 41275 -9638
rect 41367 -9682 41375 -9638
rect 41467 -9682 41475 -9638
rect 41567 -9682 41575 -9638
rect 41667 -9682 41675 -9638
rect 41767 -9682 41775 -9638
rect 41867 -9682 41875 -9638
rect 41967 -9682 41975 -9638
rect 42067 -9682 42075 -9638
rect 42167 -9682 42175 -9638
rect 42267 -9682 42275 -9638
rect 42367 -9682 42375 -9638
rect 42467 -9682 42475 -9638
rect 42567 -9682 42575 -9638
rect 42667 -9682 42675 -9638
rect 42767 -9682 42775 -9638
rect 43267 -9682 43275 -9638
rect 43367 -9682 43375 -9638
rect 43467 -9682 43475 -9638
rect 43567 -9682 43575 -9638
rect 43667 -9682 43675 -9638
rect 43767 -9682 43775 -9638
rect 43867 -9682 43875 -9638
rect 43967 -9682 43975 -9638
rect 44067 -9682 44075 -9638
rect 44167 -9682 44175 -9638
rect 44267 -9682 44275 -9638
rect 44367 -9682 44375 -9638
rect 44467 -9682 44475 -9638
rect 44567 -9682 44575 -9638
rect 44667 -9682 44675 -9638
rect 44767 -9682 44775 -9638
rect 37223 -9738 37267 -9730
rect 37323 -9738 37367 -9730
rect 37423 -9738 37467 -9730
rect 37523 -9738 37567 -9730
rect 37623 -9738 37667 -9730
rect 37723 -9738 37767 -9730
rect 37823 -9738 37867 -9730
rect 37923 -9738 37967 -9730
rect 38023 -9738 38067 -9730
rect 38123 -9738 38167 -9730
rect 38223 -9738 38267 -9730
rect 38323 -9738 38367 -9730
rect 38423 -9738 38467 -9730
rect 38523 -9738 38567 -9730
rect 38623 -9738 38667 -9730
rect 38723 -9738 38767 -9730
rect 39223 -9738 39267 -9730
rect 39323 -9738 39367 -9730
rect 39423 -9738 39467 -9730
rect 39523 -9738 39567 -9730
rect 39623 -9738 39667 -9730
rect 39723 -9738 39767 -9730
rect 39823 -9738 39867 -9730
rect 39923 -9738 39967 -9730
rect 40023 -9738 40067 -9730
rect 40123 -9738 40167 -9730
rect 40223 -9738 40267 -9730
rect 40323 -9738 40367 -9730
rect 40423 -9738 40467 -9730
rect 40523 -9738 40567 -9730
rect 40623 -9738 40667 -9730
rect 40723 -9738 40767 -9730
rect 41223 -9738 41267 -9730
rect 41323 -9738 41367 -9730
rect 41423 -9738 41467 -9730
rect 41523 -9738 41567 -9730
rect 41623 -9738 41667 -9730
rect 41723 -9738 41767 -9730
rect 41823 -9738 41867 -9730
rect 41923 -9738 41967 -9730
rect 42023 -9738 42067 -9730
rect 42123 -9738 42167 -9730
rect 42223 -9738 42267 -9730
rect 42323 -9738 42367 -9730
rect 42423 -9738 42467 -9730
rect 42523 -9738 42567 -9730
rect 42623 -9738 42667 -9730
rect 42723 -9738 42767 -9730
rect 43223 -9738 43267 -9730
rect 43323 -9738 43367 -9730
rect 43423 -9738 43467 -9730
rect 43523 -9738 43567 -9730
rect 43623 -9738 43667 -9730
rect 43723 -9738 43767 -9730
rect 43823 -9738 43867 -9730
rect 43923 -9738 43967 -9730
rect 44023 -9738 44067 -9730
rect 44123 -9738 44167 -9730
rect 44223 -9738 44267 -9730
rect 44323 -9738 44367 -9730
rect 44423 -9738 44467 -9730
rect 44523 -9738 44567 -9730
rect 44623 -9738 44667 -9730
rect 44723 -9738 44767 -9730
rect 9195 -9756 9239 -9748
rect 9295 -9756 9339 -9748
rect 9395 -9756 9439 -9748
rect 9495 -9756 9539 -9748
rect 9595 -9756 9639 -9748
rect 9695 -9756 9739 -9748
rect 9795 -9756 9839 -9748
rect 9895 -9756 9939 -9748
rect 9995 -9756 10039 -9748
rect 10095 -9756 10139 -9748
rect 10195 -9756 10239 -9748
rect 10295 -9756 10339 -9748
rect 10395 -9756 10439 -9748
rect 10495 -9756 10539 -9748
rect 10595 -9756 10639 -9748
rect 10695 -9756 10739 -9748
rect 11195 -9756 11239 -9748
rect 11295 -9756 11339 -9748
rect 11395 -9756 11439 -9748
rect 11495 -9756 11539 -9748
rect 11595 -9756 11639 -9748
rect 11695 -9756 11739 -9748
rect 11795 -9756 11839 -9748
rect 11895 -9756 11939 -9748
rect 11995 -9756 12039 -9748
rect 12095 -9756 12139 -9748
rect 12195 -9756 12239 -9748
rect 12295 -9756 12339 -9748
rect 12395 -9756 12439 -9748
rect 12495 -9756 12539 -9748
rect 12595 -9756 12639 -9748
rect 12695 -9756 12739 -9748
rect 13195 -9756 13239 -9748
rect 13295 -9756 13339 -9748
rect 13395 -9756 13439 -9748
rect 13495 -9756 13539 -9748
rect 13595 -9756 13639 -9748
rect 13695 -9756 13739 -9748
rect 13795 -9756 13839 -9748
rect 13895 -9756 13939 -9748
rect 13995 -9756 14039 -9748
rect 14095 -9756 14139 -9748
rect 14195 -9756 14239 -9748
rect 14295 -9756 14339 -9748
rect 14395 -9756 14439 -9748
rect 14495 -9756 14539 -9748
rect 14595 -9756 14639 -9748
rect 14695 -9756 14739 -9748
rect 15195 -9756 15239 -9748
rect 15295 -9756 15339 -9748
rect 15395 -9756 15439 -9748
rect 15495 -9756 15539 -9748
rect 15595 -9756 15639 -9748
rect 15695 -9756 15739 -9748
rect 15795 -9756 15839 -9748
rect 15895 -9756 15939 -9748
rect 15995 -9756 16039 -9748
rect 16095 -9756 16139 -9748
rect 16195 -9756 16239 -9748
rect 16295 -9756 16339 -9748
rect 16395 -9756 16439 -9748
rect 16495 -9756 16539 -9748
rect 16595 -9756 16639 -9748
rect 16695 -9756 16739 -9748
rect 9239 -9800 9247 -9756
rect 9339 -9800 9347 -9756
rect 9439 -9800 9447 -9756
rect 9539 -9800 9547 -9756
rect 9639 -9800 9647 -9756
rect 9739 -9800 9747 -9756
rect 9839 -9800 9847 -9756
rect 9939 -9800 9947 -9756
rect 10039 -9800 10047 -9756
rect 10139 -9800 10147 -9756
rect 10239 -9800 10247 -9756
rect 10339 -9800 10347 -9756
rect 10439 -9800 10447 -9756
rect 10539 -9800 10547 -9756
rect 10639 -9800 10647 -9756
rect 10739 -9800 10747 -9756
rect 11239 -9800 11247 -9756
rect 11339 -9800 11347 -9756
rect 11439 -9800 11447 -9756
rect 11539 -9800 11547 -9756
rect 11639 -9800 11647 -9756
rect 11739 -9800 11747 -9756
rect 11839 -9800 11847 -9756
rect 11939 -9800 11947 -9756
rect 12039 -9800 12047 -9756
rect 12139 -9800 12147 -9756
rect 12239 -9800 12247 -9756
rect 12339 -9800 12347 -9756
rect 12439 -9800 12447 -9756
rect 12539 -9800 12547 -9756
rect 12639 -9800 12647 -9756
rect 12739 -9800 12747 -9756
rect 13239 -9800 13247 -9756
rect 13339 -9800 13347 -9756
rect 13439 -9800 13447 -9756
rect 13539 -9800 13547 -9756
rect 13639 -9800 13647 -9756
rect 13739 -9800 13747 -9756
rect 13839 -9800 13847 -9756
rect 13939 -9800 13947 -9756
rect 14039 -9800 14047 -9756
rect 14139 -9800 14147 -9756
rect 14239 -9800 14247 -9756
rect 14339 -9800 14347 -9756
rect 14439 -9800 14447 -9756
rect 14539 -9800 14547 -9756
rect 14639 -9800 14647 -9756
rect 14739 -9800 14747 -9756
rect 15239 -9800 15247 -9756
rect 15339 -9800 15347 -9756
rect 15439 -9800 15447 -9756
rect 15539 -9800 15547 -9756
rect 15639 -9800 15647 -9756
rect 15739 -9800 15747 -9756
rect 15839 -9800 15847 -9756
rect 15939 -9800 15947 -9756
rect 16039 -9800 16047 -9756
rect 16139 -9800 16147 -9756
rect 16239 -9800 16247 -9756
rect 16339 -9800 16347 -9756
rect 16439 -9800 16447 -9756
rect 16539 -9800 16547 -9756
rect 16639 -9800 16647 -9756
rect 16739 -9800 16747 -9756
rect 37267 -9782 37275 -9738
rect 37367 -9782 37375 -9738
rect 37467 -9782 37475 -9738
rect 37567 -9782 37575 -9738
rect 37667 -9782 37675 -9738
rect 37767 -9782 37775 -9738
rect 37867 -9782 37875 -9738
rect 37967 -9782 37975 -9738
rect 38067 -9782 38075 -9738
rect 38167 -9782 38175 -9738
rect 38267 -9782 38275 -9738
rect 38367 -9782 38375 -9738
rect 38467 -9782 38475 -9738
rect 38567 -9782 38575 -9738
rect 38667 -9782 38675 -9738
rect 38767 -9782 38775 -9738
rect 39267 -9782 39275 -9738
rect 39367 -9782 39375 -9738
rect 39467 -9782 39475 -9738
rect 39567 -9782 39575 -9738
rect 39667 -9782 39675 -9738
rect 39767 -9782 39775 -9738
rect 39867 -9782 39875 -9738
rect 39967 -9782 39975 -9738
rect 40067 -9782 40075 -9738
rect 40167 -9782 40175 -9738
rect 40267 -9782 40275 -9738
rect 40367 -9782 40375 -9738
rect 40467 -9782 40475 -9738
rect 40567 -9782 40575 -9738
rect 40667 -9782 40675 -9738
rect 40767 -9782 40775 -9738
rect 41267 -9782 41275 -9738
rect 41367 -9782 41375 -9738
rect 41467 -9782 41475 -9738
rect 41567 -9782 41575 -9738
rect 41667 -9782 41675 -9738
rect 41767 -9782 41775 -9738
rect 41867 -9782 41875 -9738
rect 41967 -9782 41975 -9738
rect 42067 -9782 42075 -9738
rect 42167 -9782 42175 -9738
rect 42267 -9782 42275 -9738
rect 42367 -9782 42375 -9738
rect 42467 -9782 42475 -9738
rect 42567 -9782 42575 -9738
rect 42667 -9782 42675 -9738
rect 42767 -9782 42775 -9738
rect 43267 -9782 43275 -9738
rect 43367 -9782 43375 -9738
rect 43467 -9782 43475 -9738
rect 43567 -9782 43575 -9738
rect 43667 -9782 43675 -9738
rect 43767 -9782 43775 -9738
rect 43867 -9782 43875 -9738
rect 43967 -9782 43975 -9738
rect 44067 -9782 44075 -9738
rect 44167 -9782 44175 -9738
rect 44267 -9782 44275 -9738
rect 44367 -9782 44375 -9738
rect 44467 -9782 44475 -9738
rect 44567 -9782 44575 -9738
rect 44667 -9782 44675 -9738
rect 44767 -9782 44775 -9738
rect 37223 -9838 37267 -9830
rect 37323 -9838 37367 -9830
rect 37423 -9838 37467 -9830
rect 37523 -9838 37567 -9830
rect 37623 -9838 37667 -9830
rect 37723 -9838 37767 -9830
rect 37823 -9838 37867 -9830
rect 37923 -9838 37967 -9830
rect 38023 -9838 38067 -9830
rect 38123 -9838 38167 -9830
rect 38223 -9838 38267 -9830
rect 38323 -9838 38367 -9830
rect 38423 -9838 38467 -9830
rect 38523 -9838 38567 -9830
rect 38623 -9838 38667 -9830
rect 38723 -9838 38767 -9830
rect 39223 -9838 39267 -9830
rect 39323 -9838 39367 -9830
rect 39423 -9838 39467 -9830
rect 39523 -9838 39567 -9830
rect 39623 -9838 39667 -9830
rect 39723 -9838 39767 -9830
rect 39823 -9838 39867 -9830
rect 39923 -9838 39967 -9830
rect 40023 -9838 40067 -9830
rect 40123 -9838 40167 -9830
rect 40223 -9838 40267 -9830
rect 40323 -9838 40367 -9830
rect 40423 -9838 40467 -9830
rect 40523 -9838 40567 -9830
rect 40623 -9838 40667 -9830
rect 40723 -9838 40767 -9830
rect 41223 -9838 41267 -9830
rect 41323 -9838 41367 -9830
rect 41423 -9838 41467 -9830
rect 41523 -9838 41567 -9830
rect 41623 -9838 41667 -9830
rect 41723 -9838 41767 -9830
rect 41823 -9838 41867 -9830
rect 41923 -9838 41967 -9830
rect 42023 -9838 42067 -9830
rect 42123 -9838 42167 -9830
rect 42223 -9838 42267 -9830
rect 42323 -9838 42367 -9830
rect 42423 -9838 42467 -9830
rect 42523 -9838 42567 -9830
rect 42623 -9838 42667 -9830
rect 42723 -9838 42767 -9830
rect 43223 -9838 43267 -9830
rect 43323 -9838 43367 -9830
rect 43423 -9838 43467 -9830
rect 43523 -9838 43567 -9830
rect 43623 -9838 43667 -9830
rect 43723 -9838 43767 -9830
rect 43823 -9838 43867 -9830
rect 43923 -9838 43967 -9830
rect 44023 -9838 44067 -9830
rect 44123 -9838 44167 -9830
rect 44223 -9838 44267 -9830
rect 44323 -9838 44367 -9830
rect 44423 -9838 44467 -9830
rect 44523 -9838 44567 -9830
rect 44623 -9838 44667 -9830
rect 44723 -9838 44767 -9830
rect 9195 -9856 9239 -9848
rect 9295 -9856 9339 -9848
rect 9395 -9856 9439 -9848
rect 9495 -9856 9539 -9848
rect 9595 -9856 9639 -9848
rect 9695 -9856 9739 -9848
rect 9795 -9856 9839 -9848
rect 9895 -9856 9939 -9848
rect 9995 -9856 10039 -9848
rect 10095 -9856 10139 -9848
rect 10195 -9856 10239 -9848
rect 10295 -9856 10339 -9848
rect 10395 -9856 10439 -9848
rect 10495 -9856 10539 -9848
rect 10595 -9856 10639 -9848
rect 10695 -9856 10739 -9848
rect 11195 -9856 11239 -9848
rect 11295 -9856 11339 -9848
rect 11395 -9856 11439 -9848
rect 11495 -9856 11539 -9848
rect 11595 -9856 11639 -9848
rect 11695 -9856 11739 -9848
rect 11795 -9856 11839 -9848
rect 11895 -9856 11939 -9848
rect 11995 -9856 12039 -9848
rect 12095 -9856 12139 -9848
rect 12195 -9856 12239 -9848
rect 12295 -9856 12339 -9848
rect 12395 -9856 12439 -9848
rect 12495 -9856 12539 -9848
rect 12595 -9856 12639 -9848
rect 12695 -9856 12739 -9848
rect 13195 -9856 13239 -9848
rect 13295 -9856 13339 -9848
rect 13395 -9856 13439 -9848
rect 13495 -9856 13539 -9848
rect 13595 -9856 13639 -9848
rect 13695 -9856 13739 -9848
rect 13795 -9856 13839 -9848
rect 13895 -9856 13939 -9848
rect 13995 -9856 14039 -9848
rect 14095 -9856 14139 -9848
rect 14195 -9856 14239 -9848
rect 14295 -9856 14339 -9848
rect 14395 -9856 14439 -9848
rect 14495 -9856 14539 -9848
rect 14595 -9856 14639 -9848
rect 14695 -9856 14739 -9848
rect 15195 -9856 15239 -9848
rect 15295 -9856 15339 -9848
rect 15395 -9856 15439 -9848
rect 15495 -9856 15539 -9848
rect 15595 -9856 15639 -9848
rect 15695 -9856 15739 -9848
rect 15795 -9856 15839 -9848
rect 15895 -9856 15939 -9848
rect 15995 -9856 16039 -9848
rect 16095 -9856 16139 -9848
rect 16195 -9856 16239 -9848
rect 16295 -9856 16339 -9848
rect 16395 -9856 16439 -9848
rect 16495 -9856 16539 -9848
rect 16595 -9856 16639 -9848
rect 16695 -9856 16739 -9848
rect 9239 -9900 9247 -9856
rect 9339 -9900 9347 -9856
rect 9439 -9900 9447 -9856
rect 9539 -9900 9547 -9856
rect 9639 -9900 9647 -9856
rect 9739 -9900 9747 -9856
rect 9839 -9900 9847 -9856
rect 9939 -9900 9947 -9856
rect 10039 -9900 10047 -9856
rect 10139 -9900 10147 -9856
rect 10239 -9900 10247 -9856
rect 10339 -9900 10347 -9856
rect 10439 -9900 10447 -9856
rect 10539 -9900 10547 -9856
rect 10639 -9900 10647 -9856
rect 10739 -9900 10747 -9856
rect 11239 -9900 11247 -9856
rect 11339 -9900 11347 -9856
rect 11439 -9900 11447 -9856
rect 11539 -9900 11547 -9856
rect 11639 -9900 11647 -9856
rect 11739 -9900 11747 -9856
rect 11839 -9900 11847 -9856
rect 11939 -9900 11947 -9856
rect 12039 -9900 12047 -9856
rect 12139 -9900 12147 -9856
rect 12239 -9900 12247 -9856
rect 12339 -9900 12347 -9856
rect 12439 -9900 12447 -9856
rect 12539 -9900 12547 -9856
rect 12639 -9900 12647 -9856
rect 12739 -9900 12747 -9856
rect 13239 -9900 13247 -9856
rect 13339 -9900 13347 -9856
rect 13439 -9900 13447 -9856
rect 13539 -9900 13547 -9856
rect 13639 -9900 13647 -9856
rect 13739 -9900 13747 -9856
rect 13839 -9900 13847 -9856
rect 13939 -9900 13947 -9856
rect 14039 -9900 14047 -9856
rect 14139 -9900 14147 -9856
rect 14239 -9900 14247 -9856
rect 14339 -9900 14347 -9856
rect 14439 -9900 14447 -9856
rect 14539 -9900 14547 -9856
rect 14639 -9900 14647 -9856
rect 14739 -9900 14747 -9856
rect 15239 -9900 15247 -9856
rect 15339 -9900 15347 -9856
rect 15439 -9900 15447 -9856
rect 15539 -9900 15547 -9856
rect 15639 -9900 15647 -9856
rect 15739 -9900 15747 -9856
rect 15839 -9900 15847 -9856
rect 15939 -9900 15947 -9856
rect 16039 -9900 16047 -9856
rect 16139 -9900 16147 -9856
rect 16239 -9900 16247 -9856
rect 16339 -9900 16347 -9856
rect 16439 -9900 16447 -9856
rect 16539 -9900 16547 -9856
rect 16639 -9900 16647 -9856
rect 16739 -9900 16747 -9856
rect 37267 -9882 37275 -9838
rect 37367 -9882 37375 -9838
rect 37467 -9882 37475 -9838
rect 37567 -9882 37575 -9838
rect 37667 -9882 37675 -9838
rect 37767 -9882 37775 -9838
rect 37867 -9882 37875 -9838
rect 37967 -9882 37975 -9838
rect 38067 -9882 38075 -9838
rect 38167 -9882 38175 -9838
rect 38267 -9882 38275 -9838
rect 38367 -9882 38375 -9838
rect 38467 -9882 38475 -9838
rect 38567 -9882 38575 -9838
rect 38667 -9882 38675 -9838
rect 38767 -9882 38775 -9838
rect 39267 -9882 39275 -9838
rect 39367 -9882 39375 -9838
rect 39467 -9882 39475 -9838
rect 39567 -9882 39575 -9838
rect 39667 -9882 39675 -9838
rect 39767 -9882 39775 -9838
rect 39867 -9882 39875 -9838
rect 39967 -9882 39975 -9838
rect 40067 -9882 40075 -9838
rect 40167 -9882 40175 -9838
rect 40267 -9882 40275 -9838
rect 40367 -9882 40375 -9838
rect 40467 -9882 40475 -9838
rect 40567 -9882 40575 -9838
rect 40667 -9882 40675 -9838
rect 40767 -9882 40775 -9838
rect 41267 -9882 41275 -9838
rect 41367 -9882 41375 -9838
rect 41467 -9882 41475 -9838
rect 41567 -9882 41575 -9838
rect 41667 -9882 41675 -9838
rect 41767 -9882 41775 -9838
rect 41867 -9882 41875 -9838
rect 41967 -9882 41975 -9838
rect 42067 -9882 42075 -9838
rect 42167 -9882 42175 -9838
rect 42267 -9882 42275 -9838
rect 42367 -9882 42375 -9838
rect 42467 -9882 42475 -9838
rect 42567 -9882 42575 -9838
rect 42667 -9882 42675 -9838
rect 42767 -9882 42775 -9838
rect 43267 -9882 43275 -9838
rect 43367 -9882 43375 -9838
rect 43467 -9882 43475 -9838
rect 43567 -9882 43575 -9838
rect 43667 -9882 43675 -9838
rect 43767 -9882 43775 -9838
rect 43867 -9882 43875 -9838
rect 43967 -9882 43975 -9838
rect 44067 -9882 44075 -9838
rect 44167 -9882 44175 -9838
rect 44267 -9882 44275 -9838
rect 44367 -9882 44375 -9838
rect 44467 -9882 44475 -9838
rect 44567 -9882 44575 -9838
rect 44667 -9882 44675 -9838
rect 44767 -9882 44775 -9838
rect 37223 -9938 37267 -9930
rect 37323 -9938 37367 -9930
rect 37423 -9938 37467 -9930
rect 37523 -9938 37567 -9930
rect 37623 -9938 37667 -9930
rect 37723 -9938 37767 -9930
rect 37823 -9938 37867 -9930
rect 37923 -9938 37967 -9930
rect 38023 -9938 38067 -9930
rect 38123 -9938 38167 -9930
rect 38223 -9938 38267 -9930
rect 38323 -9938 38367 -9930
rect 38423 -9938 38467 -9930
rect 38523 -9938 38567 -9930
rect 38623 -9938 38667 -9930
rect 38723 -9938 38767 -9930
rect 39223 -9938 39267 -9930
rect 39323 -9938 39367 -9930
rect 39423 -9938 39467 -9930
rect 39523 -9938 39567 -9930
rect 39623 -9938 39667 -9930
rect 39723 -9938 39767 -9930
rect 39823 -9938 39867 -9930
rect 39923 -9938 39967 -9930
rect 40023 -9938 40067 -9930
rect 40123 -9938 40167 -9930
rect 40223 -9938 40267 -9930
rect 40323 -9938 40367 -9930
rect 40423 -9938 40467 -9930
rect 40523 -9938 40567 -9930
rect 40623 -9938 40667 -9930
rect 40723 -9938 40767 -9930
rect 41223 -9938 41267 -9930
rect 41323 -9938 41367 -9930
rect 41423 -9938 41467 -9930
rect 41523 -9938 41567 -9930
rect 41623 -9938 41667 -9930
rect 41723 -9938 41767 -9930
rect 41823 -9938 41867 -9930
rect 41923 -9938 41967 -9930
rect 42023 -9938 42067 -9930
rect 42123 -9938 42167 -9930
rect 42223 -9938 42267 -9930
rect 42323 -9938 42367 -9930
rect 42423 -9938 42467 -9930
rect 42523 -9938 42567 -9930
rect 42623 -9938 42667 -9930
rect 42723 -9938 42767 -9930
rect 43223 -9938 43267 -9930
rect 43323 -9938 43367 -9930
rect 43423 -9938 43467 -9930
rect 43523 -9938 43567 -9930
rect 43623 -9938 43667 -9930
rect 43723 -9938 43767 -9930
rect 43823 -9938 43867 -9930
rect 43923 -9938 43967 -9930
rect 44023 -9938 44067 -9930
rect 44123 -9938 44167 -9930
rect 44223 -9938 44267 -9930
rect 44323 -9938 44367 -9930
rect 44423 -9938 44467 -9930
rect 44523 -9938 44567 -9930
rect 44623 -9938 44667 -9930
rect 44723 -9938 44767 -9930
rect 9195 -9956 9239 -9948
rect 9295 -9956 9339 -9948
rect 9395 -9956 9439 -9948
rect 9495 -9956 9539 -9948
rect 9595 -9956 9639 -9948
rect 9695 -9956 9739 -9948
rect 9795 -9956 9839 -9948
rect 9895 -9956 9939 -9948
rect 9995 -9956 10039 -9948
rect 10095 -9956 10139 -9948
rect 10195 -9956 10239 -9948
rect 10295 -9956 10339 -9948
rect 10395 -9956 10439 -9948
rect 10495 -9956 10539 -9948
rect 10595 -9956 10639 -9948
rect 10695 -9956 10739 -9948
rect 11195 -9956 11239 -9948
rect 11295 -9956 11339 -9948
rect 11395 -9956 11439 -9948
rect 11495 -9956 11539 -9948
rect 11595 -9956 11639 -9948
rect 11695 -9956 11739 -9948
rect 11795 -9956 11839 -9948
rect 11895 -9956 11939 -9948
rect 11995 -9956 12039 -9948
rect 12095 -9956 12139 -9948
rect 12195 -9956 12239 -9948
rect 12295 -9956 12339 -9948
rect 12395 -9956 12439 -9948
rect 12495 -9956 12539 -9948
rect 12595 -9956 12639 -9948
rect 12695 -9956 12739 -9948
rect 13195 -9956 13239 -9948
rect 13295 -9956 13339 -9948
rect 13395 -9956 13439 -9948
rect 13495 -9956 13539 -9948
rect 13595 -9956 13639 -9948
rect 13695 -9956 13739 -9948
rect 13795 -9956 13839 -9948
rect 13895 -9956 13939 -9948
rect 13995 -9956 14039 -9948
rect 14095 -9956 14139 -9948
rect 14195 -9956 14239 -9948
rect 14295 -9956 14339 -9948
rect 14395 -9956 14439 -9948
rect 14495 -9956 14539 -9948
rect 14595 -9956 14639 -9948
rect 14695 -9956 14739 -9948
rect 15195 -9956 15239 -9948
rect 15295 -9956 15339 -9948
rect 15395 -9956 15439 -9948
rect 15495 -9956 15539 -9948
rect 15595 -9956 15639 -9948
rect 15695 -9956 15739 -9948
rect 15795 -9956 15839 -9948
rect 15895 -9956 15939 -9948
rect 15995 -9956 16039 -9948
rect 16095 -9956 16139 -9948
rect 16195 -9956 16239 -9948
rect 16295 -9956 16339 -9948
rect 16395 -9956 16439 -9948
rect 16495 -9956 16539 -9948
rect 16595 -9956 16639 -9948
rect 16695 -9956 16739 -9948
rect 9239 -10000 9247 -9956
rect 9339 -10000 9347 -9956
rect 9439 -10000 9447 -9956
rect 9539 -10000 9547 -9956
rect 9639 -10000 9647 -9956
rect 9739 -10000 9747 -9956
rect 9839 -10000 9847 -9956
rect 9939 -10000 9947 -9956
rect 10039 -10000 10047 -9956
rect 10139 -10000 10147 -9956
rect 10239 -10000 10247 -9956
rect 10339 -10000 10347 -9956
rect 10439 -10000 10447 -9956
rect 10539 -10000 10547 -9956
rect 10639 -10000 10647 -9956
rect 10739 -10000 10747 -9956
rect 11239 -10000 11247 -9956
rect 11339 -10000 11347 -9956
rect 11439 -10000 11447 -9956
rect 11539 -10000 11547 -9956
rect 11639 -10000 11647 -9956
rect 11739 -10000 11747 -9956
rect 11839 -10000 11847 -9956
rect 11939 -10000 11947 -9956
rect 12039 -10000 12047 -9956
rect 12139 -10000 12147 -9956
rect 12239 -10000 12247 -9956
rect 12339 -10000 12347 -9956
rect 12439 -10000 12447 -9956
rect 12539 -10000 12547 -9956
rect 12639 -10000 12647 -9956
rect 12739 -10000 12747 -9956
rect 13239 -10000 13247 -9956
rect 13339 -10000 13347 -9956
rect 13439 -10000 13447 -9956
rect 13539 -10000 13547 -9956
rect 13639 -10000 13647 -9956
rect 13739 -10000 13747 -9956
rect 13839 -10000 13847 -9956
rect 13939 -10000 13947 -9956
rect 14039 -10000 14047 -9956
rect 14139 -10000 14147 -9956
rect 14239 -10000 14247 -9956
rect 14339 -10000 14347 -9956
rect 14439 -10000 14447 -9956
rect 14539 -10000 14547 -9956
rect 14639 -10000 14647 -9956
rect 14739 -10000 14747 -9956
rect 15239 -10000 15247 -9956
rect 15339 -10000 15347 -9956
rect 15439 -10000 15447 -9956
rect 15539 -10000 15547 -9956
rect 15639 -10000 15647 -9956
rect 15739 -10000 15747 -9956
rect 15839 -10000 15847 -9956
rect 15939 -10000 15947 -9956
rect 16039 -10000 16047 -9956
rect 16139 -10000 16147 -9956
rect 16239 -10000 16247 -9956
rect 16339 -10000 16347 -9956
rect 16439 -10000 16447 -9956
rect 16539 -10000 16547 -9956
rect 16639 -10000 16647 -9956
rect 16739 -10000 16747 -9956
rect 37267 -9982 37275 -9938
rect 37367 -9982 37375 -9938
rect 37467 -9982 37475 -9938
rect 37567 -9982 37575 -9938
rect 37667 -9982 37675 -9938
rect 37767 -9982 37775 -9938
rect 37867 -9982 37875 -9938
rect 37967 -9982 37975 -9938
rect 38067 -9982 38075 -9938
rect 38167 -9982 38175 -9938
rect 38267 -9982 38275 -9938
rect 38367 -9982 38375 -9938
rect 38467 -9982 38475 -9938
rect 38567 -9982 38575 -9938
rect 38667 -9982 38675 -9938
rect 38767 -9982 38775 -9938
rect 39267 -9982 39275 -9938
rect 39367 -9982 39375 -9938
rect 39467 -9982 39475 -9938
rect 39567 -9982 39575 -9938
rect 39667 -9982 39675 -9938
rect 39767 -9982 39775 -9938
rect 39867 -9982 39875 -9938
rect 39967 -9982 39975 -9938
rect 40067 -9982 40075 -9938
rect 40167 -9982 40175 -9938
rect 40267 -9982 40275 -9938
rect 40367 -9982 40375 -9938
rect 40467 -9982 40475 -9938
rect 40567 -9982 40575 -9938
rect 40667 -9982 40675 -9938
rect 40767 -9982 40775 -9938
rect 41267 -9982 41275 -9938
rect 41367 -9982 41375 -9938
rect 41467 -9982 41475 -9938
rect 41567 -9982 41575 -9938
rect 41667 -9982 41675 -9938
rect 41767 -9982 41775 -9938
rect 41867 -9982 41875 -9938
rect 41967 -9982 41975 -9938
rect 42067 -9982 42075 -9938
rect 42167 -9982 42175 -9938
rect 42267 -9982 42275 -9938
rect 42367 -9982 42375 -9938
rect 42467 -9982 42475 -9938
rect 42567 -9982 42575 -9938
rect 42667 -9982 42675 -9938
rect 42767 -9982 42775 -9938
rect 43267 -9982 43275 -9938
rect 43367 -9982 43375 -9938
rect 43467 -9982 43475 -9938
rect 43567 -9982 43575 -9938
rect 43667 -9982 43675 -9938
rect 43767 -9982 43775 -9938
rect 43867 -9982 43875 -9938
rect 43967 -9982 43975 -9938
rect 44067 -9982 44075 -9938
rect 44167 -9982 44175 -9938
rect 44267 -9982 44275 -9938
rect 44367 -9982 44375 -9938
rect 44467 -9982 44475 -9938
rect 44567 -9982 44575 -9938
rect 44667 -9982 44675 -9938
rect 44767 -9982 44775 -9938
rect 37223 -10038 37267 -10030
rect 37323 -10038 37367 -10030
rect 37423 -10038 37467 -10030
rect 37523 -10038 37567 -10030
rect 37623 -10038 37667 -10030
rect 37723 -10038 37767 -10030
rect 37823 -10038 37867 -10030
rect 37923 -10038 37967 -10030
rect 38023 -10038 38067 -10030
rect 38123 -10038 38167 -10030
rect 38223 -10038 38267 -10030
rect 38323 -10038 38367 -10030
rect 38423 -10038 38467 -10030
rect 38523 -10038 38567 -10030
rect 38623 -10038 38667 -10030
rect 38723 -10038 38767 -10030
rect 39223 -10038 39267 -10030
rect 39323 -10038 39367 -10030
rect 39423 -10038 39467 -10030
rect 39523 -10038 39567 -10030
rect 39623 -10038 39667 -10030
rect 39723 -10038 39767 -10030
rect 39823 -10038 39867 -10030
rect 39923 -10038 39967 -10030
rect 40023 -10038 40067 -10030
rect 40123 -10038 40167 -10030
rect 40223 -10038 40267 -10030
rect 40323 -10038 40367 -10030
rect 40423 -10038 40467 -10030
rect 40523 -10038 40567 -10030
rect 40623 -10038 40667 -10030
rect 40723 -10038 40767 -10030
rect 41223 -10038 41267 -10030
rect 41323 -10038 41367 -10030
rect 41423 -10038 41467 -10030
rect 41523 -10038 41567 -10030
rect 41623 -10038 41667 -10030
rect 41723 -10038 41767 -10030
rect 41823 -10038 41867 -10030
rect 41923 -10038 41967 -10030
rect 42023 -10038 42067 -10030
rect 42123 -10038 42167 -10030
rect 42223 -10038 42267 -10030
rect 42323 -10038 42367 -10030
rect 42423 -10038 42467 -10030
rect 42523 -10038 42567 -10030
rect 42623 -10038 42667 -10030
rect 42723 -10038 42767 -10030
rect 43223 -10038 43267 -10030
rect 43323 -10038 43367 -10030
rect 43423 -10038 43467 -10030
rect 43523 -10038 43567 -10030
rect 43623 -10038 43667 -10030
rect 43723 -10038 43767 -10030
rect 43823 -10038 43867 -10030
rect 43923 -10038 43967 -10030
rect 44023 -10038 44067 -10030
rect 44123 -10038 44167 -10030
rect 44223 -10038 44267 -10030
rect 44323 -10038 44367 -10030
rect 44423 -10038 44467 -10030
rect 44523 -10038 44567 -10030
rect 44623 -10038 44667 -10030
rect 44723 -10038 44767 -10030
rect 9195 -10056 9239 -10048
rect 9295 -10056 9339 -10048
rect 9395 -10056 9439 -10048
rect 9495 -10056 9539 -10048
rect 9595 -10056 9639 -10048
rect 9695 -10056 9739 -10048
rect 9795 -10056 9839 -10048
rect 9895 -10056 9939 -10048
rect 9995 -10056 10039 -10048
rect 10095 -10056 10139 -10048
rect 10195 -10056 10239 -10048
rect 10295 -10056 10339 -10048
rect 10395 -10056 10439 -10048
rect 10495 -10056 10539 -10048
rect 10595 -10056 10639 -10048
rect 10695 -10056 10739 -10048
rect 11195 -10056 11239 -10048
rect 11295 -10056 11339 -10048
rect 11395 -10056 11439 -10048
rect 11495 -10056 11539 -10048
rect 11595 -10056 11639 -10048
rect 11695 -10056 11739 -10048
rect 11795 -10056 11839 -10048
rect 11895 -10056 11939 -10048
rect 11995 -10056 12039 -10048
rect 12095 -10056 12139 -10048
rect 12195 -10056 12239 -10048
rect 12295 -10056 12339 -10048
rect 12395 -10056 12439 -10048
rect 12495 -10056 12539 -10048
rect 12595 -10056 12639 -10048
rect 12695 -10056 12739 -10048
rect 13195 -10056 13239 -10048
rect 13295 -10056 13339 -10048
rect 13395 -10056 13439 -10048
rect 13495 -10056 13539 -10048
rect 13595 -10056 13639 -10048
rect 13695 -10056 13739 -10048
rect 13795 -10056 13839 -10048
rect 13895 -10056 13939 -10048
rect 13995 -10056 14039 -10048
rect 14095 -10056 14139 -10048
rect 14195 -10056 14239 -10048
rect 14295 -10056 14339 -10048
rect 14395 -10056 14439 -10048
rect 14495 -10056 14539 -10048
rect 14595 -10056 14639 -10048
rect 14695 -10056 14739 -10048
rect 15195 -10056 15239 -10048
rect 15295 -10056 15339 -10048
rect 15395 -10056 15439 -10048
rect 15495 -10056 15539 -10048
rect 15595 -10056 15639 -10048
rect 15695 -10056 15739 -10048
rect 15795 -10056 15839 -10048
rect 15895 -10056 15939 -10048
rect 15995 -10056 16039 -10048
rect 16095 -10056 16139 -10048
rect 16195 -10056 16239 -10048
rect 16295 -10056 16339 -10048
rect 16395 -10056 16439 -10048
rect 16495 -10056 16539 -10048
rect 16595 -10056 16639 -10048
rect 16695 -10056 16739 -10048
rect 9239 -10100 9247 -10056
rect 9339 -10100 9347 -10056
rect 9439 -10100 9447 -10056
rect 9539 -10100 9547 -10056
rect 9639 -10100 9647 -10056
rect 9739 -10100 9747 -10056
rect 9839 -10100 9847 -10056
rect 9939 -10100 9947 -10056
rect 10039 -10100 10047 -10056
rect 10139 -10100 10147 -10056
rect 10239 -10100 10247 -10056
rect 10339 -10100 10347 -10056
rect 10439 -10100 10447 -10056
rect 10539 -10100 10547 -10056
rect 10639 -10100 10647 -10056
rect 10739 -10100 10747 -10056
rect 11239 -10100 11247 -10056
rect 11339 -10100 11347 -10056
rect 11439 -10100 11447 -10056
rect 11539 -10100 11547 -10056
rect 11639 -10100 11647 -10056
rect 11739 -10100 11747 -10056
rect 11839 -10100 11847 -10056
rect 11939 -10100 11947 -10056
rect 12039 -10100 12047 -10056
rect 12139 -10100 12147 -10056
rect 12239 -10100 12247 -10056
rect 12339 -10100 12347 -10056
rect 12439 -10100 12447 -10056
rect 12539 -10100 12547 -10056
rect 12639 -10100 12647 -10056
rect 12739 -10100 12747 -10056
rect 13239 -10100 13247 -10056
rect 13339 -10100 13347 -10056
rect 13439 -10100 13447 -10056
rect 13539 -10100 13547 -10056
rect 13639 -10100 13647 -10056
rect 13739 -10100 13747 -10056
rect 13839 -10100 13847 -10056
rect 13939 -10100 13947 -10056
rect 14039 -10100 14047 -10056
rect 14139 -10100 14147 -10056
rect 14239 -10100 14247 -10056
rect 14339 -10100 14347 -10056
rect 14439 -10100 14447 -10056
rect 14539 -10100 14547 -10056
rect 14639 -10100 14647 -10056
rect 14739 -10100 14747 -10056
rect 15239 -10100 15247 -10056
rect 15339 -10100 15347 -10056
rect 15439 -10100 15447 -10056
rect 15539 -10100 15547 -10056
rect 15639 -10100 15647 -10056
rect 15739 -10100 15747 -10056
rect 15839 -10100 15847 -10056
rect 15939 -10100 15947 -10056
rect 16039 -10100 16047 -10056
rect 16139 -10100 16147 -10056
rect 16239 -10100 16247 -10056
rect 16339 -10100 16347 -10056
rect 16439 -10100 16447 -10056
rect 16539 -10100 16547 -10056
rect 16639 -10100 16647 -10056
rect 16739 -10100 16747 -10056
rect 37267 -10082 37275 -10038
rect 37367 -10082 37375 -10038
rect 37467 -10082 37475 -10038
rect 37567 -10082 37575 -10038
rect 37667 -10082 37675 -10038
rect 37767 -10082 37775 -10038
rect 37867 -10082 37875 -10038
rect 37967 -10082 37975 -10038
rect 38067 -10082 38075 -10038
rect 38167 -10082 38175 -10038
rect 38267 -10082 38275 -10038
rect 38367 -10082 38375 -10038
rect 38467 -10082 38475 -10038
rect 38567 -10082 38575 -10038
rect 38667 -10082 38675 -10038
rect 38767 -10082 38775 -10038
rect 39267 -10082 39275 -10038
rect 39367 -10082 39375 -10038
rect 39467 -10082 39475 -10038
rect 39567 -10082 39575 -10038
rect 39667 -10082 39675 -10038
rect 39767 -10082 39775 -10038
rect 39867 -10082 39875 -10038
rect 39967 -10082 39975 -10038
rect 40067 -10082 40075 -10038
rect 40167 -10082 40175 -10038
rect 40267 -10082 40275 -10038
rect 40367 -10082 40375 -10038
rect 40467 -10082 40475 -10038
rect 40567 -10082 40575 -10038
rect 40667 -10082 40675 -10038
rect 40767 -10082 40775 -10038
rect 41267 -10082 41275 -10038
rect 41367 -10082 41375 -10038
rect 41467 -10082 41475 -10038
rect 41567 -10082 41575 -10038
rect 41667 -10082 41675 -10038
rect 41767 -10082 41775 -10038
rect 41867 -10082 41875 -10038
rect 41967 -10082 41975 -10038
rect 42067 -10082 42075 -10038
rect 42167 -10082 42175 -10038
rect 42267 -10082 42275 -10038
rect 42367 -10082 42375 -10038
rect 42467 -10082 42475 -10038
rect 42567 -10082 42575 -10038
rect 42667 -10082 42675 -10038
rect 42767 -10082 42775 -10038
rect 43267 -10082 43275 -10038
rect 43367 -10082 43375 -10038
rect 43467 -10082 43475 -10038
rect 43567 -10082 43575 -10038
rect 43667 -10082 43675 -10038
rect 43767 -10082 43775 -10038
rect 43867 -10082 43875 -10038
rect 43967 -10082 43975 -10038
rect 44067 -10082 44075 -10038
rect 44167 -10082 44175 -10038
rect 44267 -10082 44275 -10038
rect 44367 -10082 44375 -10038
rect 44467 -10082 44475 -10038
rect 44567 -10082 44575 -10038
rect 44667 -10082 44675 -10038
rect 44767 -10082 44775 -10038
rect 37223 -10138 37267 -10130
rect 37323 -10138 37367 -10130
rect 37423 -10138 37467 -10130
rect 37523 -10138 37567 -10130
rect 37623 -10138 37667 -10130
rect 37723 -10138 37767 -10130
rect 37823 -10138 37867 -10130
rect 37923 -10138 37967 -10130
rect 38023 -10138 38067 -10130
rect 38123 -10138 38167 -10130
rect 38223 -10138 38267 -10130
rect 38323 -10138 38367 -10130
rect 38423 -10138 38467 -10130
rect 38523 -10138 38567 -10130
rect 38623 -10138 38667 -10130
rect 38723 -10138 38767 -10130
rect 39223 -10138 39267 -10130
rect 39323 -10138 39367 -10130
rect 39423 -10138 39467 -10130
rect 39523 -10138 39567 -10130
rect 39623 -10138 39667 -10130
rect 39723 -10138 39767 -10130
rect 39823 -10138 39867 -10130
rect 39923 -10138 39967 -10130
rect 40023 -10138 40067 -10130
rect 40123 -10138 40167 -10130
rect 40223 -10138 40267 -10130
rect 40323 -10138 40367 -10130
rect 40423 -10138 40467 -10130
rect 40523 -10138 40567 -10130
rect 40623 -10138 40667 -10130
rect 40723 -10138 40767 -10130
rect 41223 -10138 41267 -10130
rect 41323 -10138 41367 -10130
rect 41423 -10138 41467 -10130
rect 41523 -10138 41567 -10130
rect 41623 -10138 41667 -10130
rect 41723 -10138 41767 -10130
rect 41823 -10138 41867 -10130
rect 41923 -10138 41967 -10130
rect 42023 -10138 42067 -10130
rect 42123 -10138 42167 -10130
rect 42223 -10138 42267 -10130
rect 42323 -10138 42367 -10130
rect 42423 -10138 42467 -10130
rect 42523 -10138 42567 -10130
rect 42623 -10138 42667 -10130
rect 42723 -10138 42767 -10130
rect 43223 -10138 43267 -10130
rect 43323 -10138 43367 -10130
rect 43423 -10138 43467 -10130
rect 43523 -10138 43567 -10130
rect 43623 -10138 43667 -10130
rect 43723 -10138 43767 -10130
rect 43823 -10138 43867 -10130
rect 43923 -10138 43967 -10130
rect 44023 -10138 44067 -10130
rect 44123 -10138 44167 -10130
rect 44223 -10138 44267 -10130
rect 44323 -10138 44367 -10130
rect 44423 -10138 44467 -10130
rect 44523 -10138 44567 -10130
rect 44623 -10138 44667 -10130
rect 44723 -10138 44767 -10130
rect 9195 -10156 9239 -10148
rect 9295 -10156 9339 -10148
rect 9395 -10156 9439 -10148
rect 9495 -10156 9539 -10148
rect 9595 -10156 9639 -10148
rect 9695 -10156 9739 -10148
rect 9795 -10156 9839 -10148
rect 9895 -10156 9939 -10148
rect 9995 -10156 10039 -10148
rect 10095 -10156 10139 -10148
rect 10195 -10156 10239 -10148
rect 10295 -10156 10339 -10148
rect 10395 -10156 10439 -10148
rect 10495 -10156 10539 -10148
rect 10595 -10156 10639 -10148
rect 10695 -10156 10739 -10148
rect 11195 -10156 11239 -10148
rect 11295 -10156 11339 -10148
rect 11395 -10156 11439 -10148
rect 11495 -10156 11539 -10148
rect 11595 -10156 11639 -10148
rect 11695 -10156 11739 -10148
rect 11795 -10156 11839 -10148
rect 11895 -10156 11939 -10148
rect 11995 -10156 12039 -10148
rect 12095 -10156 12139 -10148
rect 12195 -10156 12239 -10148
rect 12295 -10156 12339 -10148
rect 12395 -10156 12439 -10148
rect 12495 -10156 12539 -10148
rect 12595 -10156 12639 -10148
rect 12695 -10156 12739 -10148
rect 13195 -10156 13239 -10148
rect 13295 -10156 13339 -10148
rect 13395 -10156 13439 -10148
rect 13495 -10156 13539 -10148
rect 13595 -10156 13639 -10148
rect 13695 -10156 13739 -10148
rect 13795 -10156 13839 -10148
rect 13895 -10156 13939 -10148
rect 13995 -10156 14039 -10148
rect 14095 -10156 14139 -10148
rect 14195 -10156 14239 -10148
rect 14295 -10156 14339 -10148
rect 14395 -10156 14439 -10148
rect 14495 -10156 14539 -10148
rect 14595 -10156 14639 -10148
rect 14695 -10156 14739 -10148
rect 15195 -10156 15239 -10148
rect 15295 -10156 15339 -10148
rect 15395 -10156 15439 -10148
rect 15495 -10156 15539 -10148
rect 15595 -10156 15639 -10148
rect 15695 -10156 15739 -10148
rect 15795 -10156 15839 -10148
rect 15895 -10156 15939 -10148
rect 15995 -10156 16039 -10148
rect 16095 -10156 16139 -10148
rect 16195 -10156 16239 -10148
rect 16295 -10156 16339 -10148
rect 16395 -10156 16439 -10148
rect 16495 -10156 16539 -10148
rect 16595 -10156 16639 -10148
rect 16695 -10156 16739 -10148
rect 9239 -10200 9247 -10156
rect 9339 -10200 9347 -10156
rect 9439 -10200 9447 -10156
rect 9539 -10200 9547 -10156
rect 9639 -10200 9647 -10156
rect 9739 -10200 9747 -10156
rect 9839 -10200 9847 -10156
rect 9939 -10200 9947 -10156
rect 10039 -10200 10047 -10156
rect 10139 -10200 10147 -10156
rect 10239 -10200 10247 -10156
rect 10339 -10200 10347 -10156
rect 10439 -10200 10447 -10156
rect 10539 -10200 10547 -10156
rect 10639 -10200 10647 -10156
rect 10739 -10200 10747 -10156
rect 11239 -10200 11247 -10156
rect 11339 -10200 11347 -10156
rect 11439 -10200 11447 -10156
rect 11539 -10200 11547 -10156
rect 11639 -10200 11647 -10156
rect 11739 -10200 11747 -10156
rect 11839 -10200 11847 -10156
rect 11939 -10200 11947 -10156
rect 12039 -10200 12047 -10156
rect 12139 -10200 12147 -10156
rect 12239 -10200 12247 -10156
rect 12339 -10200 12347 -10156
rect 12439 -10200 12447 -10156
rect 12539 -10200 12547 -10156
rect 12639 -10200 12647 -10156
rect 12739 -10200 12747 -10156
rect 13239 -10200 13247 -10156
rect 13339 -10200 13347 -10156
rect 13439 -10200 13447 -10156
rect 13539 -10200 13547 -10156
rect 13639 -10200 13647 -10156
rect 13739 -10200 13747 -10156
rect 13839 -10200 13847 -10156
rect 13939 -10200 13947 -10156
rect 14039 -10200 14047 -10156
rect 14139 -10200 14147 -10156
rect 14239 -10200 14247 -10156
rect 14339 -10200 14347 -10156
rect 14439 -10200 14447 -10156
rect 14539 -10200 14547 -10156
rect 14639 -10200 14647 -10156
rect 14739 -10200 14747 -10156
rect 15239 -10200 15247 -10156
rect 15339 -10200 15347 -10156
rect 15439 -10200 15447 -10156
rect 15539 -10200 15547 -10156
rect 15639 -10200 15647 -10156
rect 15739 -10200 15747 -10156
rect 15839 -10200 15847 -10156
rect 15939 -10200 15947 -10156
rect 16039 -10200 16047 -10156
rect 16139 -10200 16147 -10156
rect 16239 -10200 16247 -10156
rect 16339 -10200 16347 -10156
rect 16439 -10200 16447 -10156
rect 16539 -10200 16547 -10156
rect 16639 -10200 16647 -10156
rect 16739 -10200 16747 -10156
rect 37267 -10182 37275 -10138
rect 37367 -10182 37375 -10138
rect 37467 -10182 37475 -10138
rect 37567 -10182 37575 -10138
rect 37667 -10182 37675 -10138
rect 37767 -10182 37775 -10138
rect 37867 -10182 37875 -10138
rect 37967 -10182 37975 -10138
rect 38067 -10182 38075 -10138
rect 38167 -10182 38175 -10138
rect 38267 -10182 38275 -10138
rect 38367 -10182 38375 -10138
rect 38467 -10182 38475 -10138
rect 38567 -10182 38575 -10138
rect 38667 -10182 38675 -10138
rect 38767 -10182 38775 -10138
rect 39267 -10182 39275 -10138
rect 39367 -10182 39375 -10138
rect 39467 -10182 39475 -10138
rect 39567 -10182 39575 -10138
rect 39667 -10182 39675 -10138
rect 39767 -10182 39775 -10138
rect 39867 -10182 39875 -10138
rect 39967 -10182 39975 -10138
rect 40067 -10182 40075 -10138
rect 40167 -10182 40175 -10138
rect 40267 -10182 40275 -10138
rect 40367 -10182 40375 -10138
rect 40467 -10182 40475 -10138
rect 40567 -10182 40575 -10138
rect 40667 -10182 40675 -10138
rect 40767 -10182 40775 -10138
rect 41267 -10182 41275 -10138
rect 41367 -10182 41375 -10138
rect 41467 -10182 41475 -10138
rect 41567 -10182 41575 -10138
rect 41667 -10182 41675 -10138
rect 41767 -10182 41775 -10138
rect 41867 -10182 41875 -10138
rect 41967 -10182 41975 -10138
rect 42067 -10182 42075 -10138
rect 42167 -10182 42175 -10138
rect 42267 -10182 42275 -10138
rect 42367 -10182 42375 -10138
rect 42467 -10182 42475 -10138
rect 42567 -10182 42575 -10138
rect 42667 -10182 42675 -10138
rect 42767 -10182 42775 -10138
rect 43267 -10182 43275 -10138
rect 43367 -10182 43375 -10138
rect 43467 -10182 43475 -10138
rect 43567 -10182 43575 -10138
rect 43667 -10182 43675 -10138
rect 43767 -10182 43775 -10138
rect 43867 -10182 43875 -10138
rect 43967 -10182 43975 -10138
rect 44067 -10182 44075 -10138
rect 44167 -10182 44175 -10138
rect 44267 -10182 44275 -10138
rect 44367 -10182 44375 -10138
rect 44467 -10182 44475 -10138
rect 44567 -10182 44575 -10138
rect 44667 -10182 44675 -10138
rect 44767 -10182 44775 -10138
rect 37223 -10238 37267 -10230
rect 37323 -10238 37367 -10230
rect 37423 -10238 37467 -10230
rect 37523 -10238 37567 -10230
rect 37623 -10238 37667 -10230
rect 37723 -10238 37767 -10230
rect 37823 -10238 37867 -10230
rect 37923 -10238 37967 -10230
rect 38023 -10238 38067 -10230
rect 38123 -10238 38167 -10230
rect 38223 -10238 38267 -10230
rect 38323 -10238 38367 -10230
rect 38423 -10238 38467 -10230
rect 38523 -10238 38567 -10230
rect 38623 -10238 38667 -10230
rect 38723 -10238 38767 -10230
rect 39223 -10238 39267 -10230
rect 39323 -10238 39367 -10230
rect 39423 -10238 39467 -10230
rect 39523 -10238 39567 -10230
rect 39623 -10238 39667 -10230
rect 39723 -10238 39767 -10230
rect 39823 -10238 39867 -10230
rect 39923 -10238 39967 -10230
rect 40023 -10238 40067 -10230
rect 40123 -10238 40167 -10230
rect 40223 -10238 40267 -10230
rect 40323 -10238 40367 -10230
rect 40423 -10238 40467 -10230
rect 40523 -10238 40567 -10230
rect 40623 -10238 40667 -10230
rect 40723 -10238 40767 -10230
rect 41223 -10238 41267 -10230
rect 41323 -10238 41367 -10230
rect 41423 -10238 41467 -10230
rect 41523 -10238 41567 -10230
rect 41623 -10238 41667 -10230
rect 41723 -10238 41767 -10230
rect 41823 -10238 41867 -10230
rect 41923 -10238 41967 -10230
rect 42023 -10238 42067 -10230
rect 42123 -10238 42167 -10230
rect 42223 -10238 42267 -10230
rect 42323 -10238 42367 -10230
rect 42423 -10238 42467 -10230
rect 42523 -10238 42567 -10230
rect 42623 -10238 42667 -10230
rect 42723 -10238 42767 -10230
rect 43223 -10238 43267 -10230
rect 43323 -10238 43367 -10230
rect 43423 -10238 43467 -10230
rect 43523 -10238 43567 -10230
rect 43623 -10238 43667 -10230
rect 43723 -10238 43767 -10230
rect 43823 -10238 43867 -10230
rect 43923 -10238 43967 -10230
rect 44023 -10238 44067 -10230
rect 44123 -10238 44167 -10230
rect 44223 -10238 44267 -10230
rect 44323 -10238 44367 -10230
rect 44423 -10238 44467 -10230
rect 44523 -10238 44567 -10230
rect 44623 -10238 44667 -10230
rect 44723 -10238 44767 -10230
rect 9195 -10256 9239 -10248
rect 9295 -10256 9339 -10248
rect 9395 -10256 9439 -10248
rect 9495 -10256 9539 -10248
rect 9595 -10256 9639 -10248
rect 9695 -10256 9739 -10248
rect 9795 -10256 9839 -10248
rect 9895 -10256 9939 -10248
rect 9995 -10256 10039 -10248
rect 10095 -10256 10139 -10248
rect 10195 -10256 10239 -10248
rect 10295 -10256 10339 -10248
rect 10395 -10256 10439 -10248
rect 10495 -10256 10539 -10248
rect 10595 -10256 10639 -10248
rect 10695 -10256 10739 -10248
rect 11195 -10256 11239 -10248
rect 11295 -10256 11339 -10248
rect 11395 -10256 11439 -10248
rect 11495 -10256 11539 -10248
rect 11595 -10256 11639 -10248
rect 11695 -10256 11739 -10248
rect 11795 -10256 11839 -10248
rect 11895 -10256 11939 -10248
rect 11995 -10256 12039 -10248
rect 12095 -10256 12139 -10248
rect 12195 -10256 12239 -10248
rect 12295 -10256 12339 -10248
rect 12395 -10256 12439 -10248
rect 12495 -10256 12539 -10248
rect 12595 -10256 12639 -10248
rect 12695 -10256 12739 -10248
rect 13195 -10256 13239 -10248
rect 13295 -10256 13339 -10248
rect 13395 -10256 13439 -10248
rect 13495 -10256 13539 -10248
rect 13595 -10256 13639 -10248
rect 13695 -10256 13739 -10248
rect 13795 -10256 13839 -10248
rect 13895 -10256 13939 -10248
rect 13995 -10256 14039 -10248
rect 14095 -10256 14139 -10248
rect 14195 -10256 14239 -10248
rect 14295 -10256 14339 -10248
rect 14395 -10256 14439 -10248
rect 14495 -10256 14539 -10248
rect 14595 -10256 14639 -10248
rect 14695 -10256 14739 -10248
rect 15195 -10256 15239 -10248
rect 15295 -10256 15339 -10248
rect 15395 -10256 15439 -10248
rect 15495 -10256 15539 -10248
rect 15595 -10256 15639 -10248
rect 15695 -10256 15739 -10248
rect 15795 -10256 15839 -10248
rect 15895 -10256 15939 -10248
rect 15995 -10256 16039 -10248
rect 16095 -10256 16139 -10248
rect 16195 -10256 16239 -10248
rect 16295 -10256 16339 -10248
rect 16395 -10256 16439 -10248
rect 16495 -10256 16539 -10248
rect 16595 -10256 16639 -10248
rect 16695 -10256 16739 -10248
rect 9239 -10300 9247 -10256
rect 9339 -10300 9347 -10256
rect 9439 -10300 9447 -10256
rect 9539 -10300 9547 -10256
rect 9639 -10300 9647 -10256
rect 9739 -10300 9747 -10256
rect 9839 -10300 9847 -10256
rect 9939 -10300 9947 -10256
rect 10039 -10300 10047 -10256
rect 10139 -10300 10147 -10256
rect 10239 -10300 10247 -10256
rect 10339 -10300 10347 -10256
rect 10439 -10300 10447 -10256
rect 10539 -10300 10547 -10256
rect 10639 -10300 10647 -10256
rect 10739 -10300 10747 -10256
rect 11239 -10300 11247 -10256
rect 11339 -10300 11347 -10256
rect 11439 -10300 11447 -10256
rect 11539 -10300 11547 -10256
rect 11639 -10300 11647 -10256
rect 11739 -10300 11747 -10256
rect 11839 -10300 11847 -10256
rect 11939 -10300 11947 -10256
rect 12039 -10300 12047 -10256
rect 12139 -10300 12147 -10256
rect 12239 -10300 12247 -10256
rect 12339 -10300 12347 -10256
rect 12439 -10300 12447 -10256
rect 12539 -10300 12547 -10256
rect 12639 -10300 12647 -10256
rect 12739 -10300 12747 -10256
rect 13239 -10300 13247 -10256
rect 13339 -10300 13347 -10256
rect 13439 -10300 13447 -10256
rect 13539 -10300 13547 -10256
rect 13639 -10300 13647 -10256
rect 13739 -10300 13747 -10256
rect 13839 -10300 13847 -10256
rect 13939 -10300 13947 -10256
rect 14039 -10300 14047 -10256
rect 14139 -10300 14147 -10256
rect 14239 -10300 14247 -10256
rect 14339 -10300 14347 -10256
rect 14439 -10300 14447 -10256
rect 14539 -10300 14547 -10256
rect 14639 -10300 14647 -10256
rect 14739 -10300 14747 -10256
rect 15239 -10300 15247 -10256
rect 15339 -10300 15347 -10256
rect 15439 -10300 15447 -10256
rect 15539 -10300 15547 -10256
rect 15639 -10300 15647 -10256
rect 15739 -10300 15747 -10256
rect 15839 -10300 15847 -10256
rect 15939 -10300 15947 -10256
rect 16039 -10300 16047 -10256
rect 16139 -10300 16147 -10256
rect 16239 -10300 16247 -10256
rect 16339 -10300 16347 -10256
rect 16439 -10300 16447 -10256
rect 16539 -10300 16547 -10256
rect 16639 -10300 16647 -10256
rect 16739 -10300 16747 -10256
rect 37267 -10282 37275 -10238
rect 37367 -10282 37375 -10238
rect 37467 -10282 37475 -10238
rect 37567 -10282 37575 -10238
rect 37667 -10282 37675 -10238
rect 37767 -10282 37775 -10238
rect 37867 -10282 37875 -10238
rect 37967 -10282 37975 -10238
rect 38067 -10282 38075 -10238
rect 38167 -10282 38175 -10238
rect 38267 -10282 38275 -10238
rect 38367 -10282 38375 -10238
rect 38467 -10282 38475 -10238
rect 38567 -10282 38575 -10238
rect 38667 -10282 38675 -10238
rect 38767 -10282 38775 -10238
rect 39267 -10282 39275 -10238
rect 39367 -10282 39375 -10238
rect 39467 -10282 39475 -10238
rect 39567 -10282 39575 -10238
rect 39667 -10282 39675 -10238
rect 39767 -10282 39775 -10238
rect 39867 -10282 39875 -10238
rect 39967 -10282 39975 -10238
rect 40067 -10282 40075 -10238
rect 40167 -10282 40175 -10238
rect 40267 -10282 40275 -10238
rect 40367 -10282 40375 -10238
rect 40467 -10282 40475 -10238
rect 40567 -10282 40575 -10238
rect 40667 -10282 40675 -10238
rect 40767 -10282 40775 -10238
rect 41267 -10282 41275 -10238
rect 41367 -10282 41375 -10238
rect 41467 -10282 41475 -10238
rect 41567 -10282 41575 -10238
rect 41667 -10282 41675 -10238
rect 41767 -10282 41775 -10238
rect 41867 -10282 41875 -10238
rect 41967 -10282 41975 -10238
rect 42067 -10282 42075 -10238
rect 42167 -10282 42175 -10238
rect 42267 -10282 42275 -10238
rect 42367 -10282 42375 -10238
rect 42467 -10282 42475 -10238
rect 42567 -10282 42575 -10238
rect 42667 -10282 42675 -10238
rect 42767 -10282 42775 -10238
rect 43267 -10282 43275 -10238
rect 43367 -10282 43375 -10238
rect 43467 -10282 43475 -10238
rect 43567 -10282 43575 -10238
rect 43667 -10282 43675 -10238
rect 43767 -10282 43775 -10238
rect 43867 -10282 43875 -10238
rect 43967 -10282 43975 -10238
rect 44067 -10282 44075 -10238
rect 44167 -10282 44175 -10238
rect 44267 -10282 44275 -10238
rect 44367 -10282 44375 -10238
rect 44467 -10282 44475 -10238
rect 44567 -10282 44575 -10238
rect 44667 -10282 44675 -10238
rect 44767 -10282 44775 -10238
rect 37223 -10338 37267 -10330
rect 37323 -10338 37367 -10330
rect 37423 -10338 37467 -10330
rect 37523 -10338 37567 -10330
rect 37623 -10338 37667 -10330
rect 37723 -10338 37767 -10330
rect 37823 -10338 37867 -10330
rect 37923 -10338 37967 -10330
rect 38023 -10338 38067 -10330
rect 38123 -10338 38167 -10330
rect 38223 -10338 38267 -10330
rect 38323 -10338 38367 -10330
rect 38423 -10338 38467 -10330
rect 38523 -10338 38567 -10330
rect 38623 -10338 38667 -10330
rect 38723 -10338 38767 -10330
rect 39223 -10338 39267 -10330
rect 39323 -10338 39367 -10330
rect 39423 -10338 39467 -10330
rect 39523 -10338 39567 -10330
rect 39623 -10338 39667 -10330
rect 39723 -10338 39767 -10330
rect 39823 -10338 39867 -10330
rect 39923 -10338 39967 -10330
rect 40023 -10338 40067 -10330
rect 40123 -10338 40167 -10330
rect 40223 -10338 40267 -10330
rect 40323 -10338 40367 -10330
rect 40423 -10338 40467 -10330
rect 40523 -10338 40567 -10330
rect 40623 -10338 40667 -10330
rect 40723 -10338 40767 -10330
rect 41223 -10338 41267 -10330
rect 41323 -10338 41367 -10330
rect 41423 -10338 41467 -10330
rect 41523 -10338 41567 -10330
rect 41623 -10338 41667 -10330
rect 41723 -10338 41767 -10330
rect 41823 -10338 41867 -10330
rect 41923 -10338 41967 -10330
rect 42023 -10338 42067 -10330
rect 42123 -10338 42167 -10330
rect 42223 -10338 42267 -10330
rect 42323 -10338 42367 -10330
rect 42423 -10338 42467 -10330
rect 42523 -10338 42567 -10330
rect 42623 -10338 42667 -10330
rect 42723 -10338 42767 -10330
rect 43223 -10338 43267 -10330
rect 43323 -10338 43367 -10330
rect 43423 -10338 43467 -10330
rect 43523 -10338 43567 -10330
rect 43623 -10338 43667 -10330
rect 43723 -10338 43767 -10330
rect 43823 -10338 43867 -10330
rect 43923 -10338 43967 -10330
rect 44023 -10338 44067 -10330
rect 44123 -10338 44167 -10330
rect 44223 -10338 44267 -10330
rect 44323 -10338 44367 -10330
rect 44423 -10338 44467 -10330
rect 44523 -10338 44567 -10330
rect 44623 -10338 44667 -10330
rect 44723 -10338 44767 -10330
rect 9195 -10356 9239 -10348
rect 9295 -10356 9339 -10348
rect 9395 -10356 9439 -10348
rect 9495 -10356 9539 -10348
rect 9595 -10356 9639 -10348
rect 9695 -10356 9739 -10348
rect 9795 -10356 9839 -10348
rect 9895 -10356 9939 -10348
rect 9995 -10356 10039 -10348
rect 10095 -10356 10139 -10348
rect 10195 -10356 10239 -10348
rect 10295 -10356 10339 -10348
rect 10395 -10356 10439 -10348
rect 10495 -10356 10539 -10348
rect 10595 -10356 10639 -10348
rect 10695 -10356 10739 -10348
rect 11195 -10356 11239 -10348
rect 11295 -10356 11339 -10348
rect 11395 -10356 11439 -10348
rect 11495 -10356 11539 -10348
rect 11595 -10356 11639 -10348
rect 11695 -10356 11739 -10348
rect 11795 -10356 11839 -10348
rect 11895 -10356 11939 -10348
rect 11995 -10356 12039 -10348
rect 12095 -10356 12139 -10348
rect 12195 -10356 12239 -10348
rect 12295 -10356 12339 -10348
rect 12395 -10356 12439 -10348
rect 12495 -10356 12539 -10348
rect 12595 -10356 12639 -10348
rect 12695 -10356 12739 -10348
rect 13195 -10356 13239 -10348
rect 13295 -10356 13339 -10348
rect 13395 -10356 13439 -10348
rect 13495 -10356 13539 -10348
rect 13595 -10356 13639 -10348
rect 13695 -10356 13739 -10348
rect 13795 -10356 13839 -10348
rect 13895 -10356 13939 -10348
rect 13995 -10356 14039 -10348
rect 14095 -10356 14139 -10348
rect 14195 -10356 14239 -10348
rect 14295 -10356 14339 -10348
rect 14395 -10356 14439 -10348
rect 14495 -10356 14539 -10348
rect 14595 -10356 14639 -10348
rect 14695 -10356 14739 -10348
rect 15195 -10356 15239 -10348
rect 15295 -10356 15339 -10348
rect 15395 -10356 15439 -10348
rect 15495 -10356 15539 -10348
rect 15595 -10356 15639 -10348
rect 15695 -10356 15739 -10348
rect 15795 -10356 15839 -10348
rect 15895 -10356 15939 -10348
rect 15995 -10356 16039 -10348
rect 16095 -10356 16139 -10348
rect 16195 -10356 16239 -10348
rect 16295 -10356 16339 -10348
rect 16395 -10356 16439 -10348
rect 16495 -10356 16539 -10348
rect 16595 -10356 16639 -10348
rect 16695 -10356 16739 -10348
rect 9239 -10400 9247 -10356
rect 9339 -10400 9347 -10356
rect 9439 -10400 9447 -10356
rect 9539 -10400 9547 -10356
rect 9639 -10400 9647 -10356
rect 9739 -10400 9747 -10356
rect 9839 -10400 9847 -10356
rect 9939 -10400 9947 -10356
rect 10039 -10400 10047 -10356
rect 10139 -10400 10147 -10356
rect 10239 -10400 10247 -10356
rect 10339 -10400 10347 -10356
rect 10439 -10400 10447 -10356
rect 10539 -10400 10547 -10356
rect 10639 -10400 10647 -10356
rect 10739 -10400 10747 -10356
rect 11239 -10400 11247 -10356
rect 11339 -10400 11347 -10356
rect 11439 -10400 11447 -10356
rect 11539 -10400 11547 -10356
rect 11639 -10400 11647 -10356
rect 11739 -10400 11747 -10356
rect 11839 -10400 11847 -10356
rect 11939 -10400 11947 -10356
rect 12039 -10400 12047 -10356
rect 12139 -10400 12147 -10356
rect 12239 -10400 12247 -10356
rect 12339 -10400 12347 -10356
rect 12439 -10400 12447 -10356
rect 12539 -10400 12547 -10356
rect 12639 -10400 12647 -10356
rect 12739 -10400 12747 -10356
rect 13239 -10400 13247 -10356
rect 13339 -10400 13347 -10356
rect 13439 -10400 13447 -10356
rect 13539 -10400 13547 -10356
rect 13639 -10400 13647 -10356
rect 13739 -10400 13747 -10356
rect 13839 -10400 13847 -10356
rect 13939 -10400 13947 -10356
rect 14039 -10400 14047 -10356
rect 14139 -10400 14147 -10356
rect 14239 -10400 14247 -10356
rect 14339 -10400 14347 -10356
rect 14439 -10400 14447 -10356
rect 14539 -10400 14547 -10356
rect 14639 -10400 14647 -10356
rect 14739 -10400 14747 -10356
rect 15239 -10400 15247 -10356
rect 15339 -10400 15347 -10356
rect 15439 -10400 15447 -10356
rect 15539 -10400 15547 -10356
rect 15639 -10400 15647 -10356
rect 15739 -10400 15747 -10356
rect 15839 -10400 15847 -10356
rect 15939 -10400 15947 -10356
rect 16039 -10400 16047 -10356
rect 16139 -10400 16147 -10356
rect 16239 -10400 16247 -10356
rect 16339 -10400 16347 -10356
rect 16439 -10400 16447 -10356
rect 16539 -10400 16547 -10356
rect 16639 -10400 16647 -10356
rect 16739 -10400 16747 -10356
rect 37267 -10382 37275 -10338
rect 37367 -10382 37375 -10338
rect 37467 -10382 37475 -10338
rect 37567 -10382 37575 -10338
rect 37667 -10382 37675 -10338
rect 37767 -10382 37775 -10338
rect 37867 -10382 37875 -10338
rect 37967 -10382 37975 -10338
rect 38067 -10382 38075 -10338
rect 38167 -10382 38175 -10338
rect 38267 -10382 38275 -10338
rect 38367 -10382 38375 -10338
rect 38467 -10382 38475 -10338
rect 38567 -10382 38575 -10338
rect 38667 -10382 38675 -10338
rect 38767 -10382 38775 -10338
rect 39267 -10382 39275 -10338
rect 39367 -10382 39375 -10338
rect 39467 -10382 39475 -10338
rect 39567 -10382 39575 -10338
rect 39667 -10382 39675 -10338
rect 39767 -10382 39775 -10338
rect 39867 -10382 39875 -10338
rect 39967 -10382 39975 -10338
rect 40067 -10382 40075 -10338
rect 40167 -10382 40175 -10338
rect 40267 -10382 40275 -10338
rect 40367 -10382 40375 -10338
rect 40467 -10382 40475 -10338
rect 40567 -10382 40575 -10338
rect 40667 -10382 40675 -10338
rect 40767 -10382 40775 -10338
rect 41267 -10382 41275 -10338
rect 41367 -10382 41375 -10338
rect 41467 -10382 41475 -10338
rect 41567 -10382 41575 -10338
rect 41667 -10382 41675 -10338
rect 41767 -10382 41775 -10338
rect 41867 -10382 41875 -10338
rect 41967 -10382 41975 -10338
rect 42067 -10382 42075 -10338
rect 42167 -10382 42175 -10338
rect 42267 -10382 42275 -10338
rect 42367 -10382 42375 -10338
rect 42467 -10382 42475 -10338
rect 42567 -10382 42575 -10338
rect 42667 -10382 42675 -10338
rect 42767 -10382 42775 -10338
rect 43267 -10382 43275 -10338
rect 43367 -10382 43375 -10338
rect 43467 -10382 43475 -10338
rect 43567 -10382 43575 -10338
rect 43667 -10382 43675 -10338
rect 43767 -10382 43775 -10338
rect 43867 -10382 43875 -10338
rect 43967 -10382 43975 -10338
rect 44067 -10382 44075 -10338
rect 44167 -10382 44175 -10338
rect 44267 -10382 44275 -10338
rect 44367 -10382 44375 -10338
rect 44467 -10382 44475 -10338
rect 44567 -10382 44575 -10338
rect 44667 -10382 44675 -10338
rect 44767 -10382 44775 -10338
rect 37223 -10438 37267 -10430
rect 37323 -10438 37367 -10430
rect 37423 -10438 37467 -10430
rect 37523 -10438 37567 -10430
rect 37623 -10438 37667 -10430
rect 37723 -10438 37767 -10430
rect 37823 -10438 37867 -10430
rect 37923 -10438 37967 -10430
rect 38023 -10438 38067 -10430
rect 38123 -10438 38167 -10430
rect 38223 -10438 38267 -10430
rect 38323 -10438 38367 -10430
rect 38423 -10438 38467 -10430
rect 38523 -10438 38567 -10430
rect 38623 -10438 38667 -10430
rect 38723 -10438 38767 -10430
rect 39223 -10438 39267 -10430
rect 39323 -10438 39367 -10430
rect 39423 -10438 39467 -10430
rect 39523 -10438 39567 -10430
rect 39623 -10438 39667 -10430
rect 39723 -10438 39767 -10430
rect 39823 -10438 39867 -10430
rect 39923 -10438 39967 -10430
rect 40023 -10438 40067 -10430
rect 40123 -10438 40167 -10430
rect 40223 -10438 40267 -10430
rect 40323 -10438 40367 -10430
rect 40423 -10438 40467 -10430
rect 40523 -10438 40567 -10430
rect 40623 -10438 40667 -10430
rect 40723 -10438 40767 -10430
rect 41223 -10438 41267 -10430
rect 41323 -10438 41367 -10430
rect 41423 -10438 41467 -10430
rect 41523 -10438 41567 -10430
rect 41623 -10438 41667 -10430
rect 41723 -10438 41767 -10430
rect 41823 -10438 41867 -10430
rect 41923 -10438 41967 -10430
rect 42023 -10438 42067 -10430
rect 42123 -10438 42167 -10430
rect 42223 -10438 42267 -10430
rect 42323 -10438 42367 -10430
rect 42423 -10438 42467 -10430
rect 42523 -10438 42567 -10430
rect 42623 -10438 42667 -10430
rect 42723 -10438 42767 -10430
rect 43223 -10438 43267 -10430
rect 43323 -10438 43367 -10430
rect 43423 -10438 43467 -10430
rect 43523 -10438 43567 -10430
rect 43623 -10438 43667 -10430
rect 43723 -10438 43767 -10430
rect 43823 -10438 43867 -10430
rect 43923 -10438 43967 -10430
rect 44023 -10438 44067 -10430
rect 44123 -10438 44167 -10430
rect 44223 -10438 44267 -10430
rect 44323 -10438 44367 -10430
rect 44423 -10438 44467 -10430
rect 44523 -10438 44567 -10430
rect 44623 -10438 44667 -10430
rect 44723 -10438 44767 -10430
rect 9195 -10456 9239 -10448
rect 9295 -10456 9339 -10448
rect 9395 -10456 9439 -10448
rect 9495 -10456 9539 -10448
rect 9595 -10456 9639 -10448
rect 9695 -10456 9739 -10448
rect 9795 -10456 9839 -10448
rect 9895 -10456 9939 -10448
rect 9995 -10456 10039 -10448
rect 10095 -10456 10139 -10448
rect 10195 -10456 10239 -10448
rect 10295 -10456 10339 -10448
rect 10395 -10456 10439 -10448
rect 10495 -10456 10539 -10448
rect 10595 -10456 10639 -10448
rect 10695 -10456 10739 -10448
rect 11195 -10456 11239 -10448
rect 11295 -10456 11339 -10448
rect 11395 -10456 11439 -10448
rect 11495 -10456 11539 -10448
rect 11595 -10456 11639 -10448
rect 11695 -10456 11739 -10448
rect 11795 -10456 11839 -10448
rect 11895 -10456 11939 -10448
rect 11995 -10456 12039 -10448
rect 12095 -10456 12139 -10448
rect 12195 -10456 12239 -10448
rect 12295 -10456 12339 -10448
rect 12395 -10456 12439 -10448
rect 12495 -10456 12539 -10448
rect 12595 -10456 12639 -10448
rect 12695 -10456 12739 -10448
rect 13195 -10456 13239 -10448
rect 13295 -10456 13339 -10448
rect 13395 -10456 13439 -10448
rect 13495 -10456 13539 -10448
rect 13595 -10456 13639 -10448
rect 13695 -10456 13739 -10448
rect 13795 -10456 13839 -10448
rect 13895 -10456 13939 -10448
rect 13995 -10456 14039 -10448
rect 14095 -10456 14139 -10448
rect 14195 -10456 14239 -10448
rect 14295 -10456 14339 -10448
rect 14395 -10456 14439 -10448
rect 14495 -10456 14539 -10448
rect 14595 -10456 14639 -10448
rect 14695 -10456 14739 -10448
rect 15195 -10456 15239 -10448
rect 15295 -10456 15339 -10448
rect 15395 -10456 15439 -10448
rect 15495 -10456 15539 -10448
rect 15595 -10456 15639 -10448
rect 15695 -10456 15739 -10448
rect 15795 -10456 15839 -10448
rect 15895 -10456 15939 -10448
rect 15995 -10456 16039 -10448
rect 16095 -10456 16139 -10448
rect 16195 -10456 16239 -10448
rect 16295 -10456 16339 -10448
rect 16395 -10456 16439 -10448
rect 16495 -10456 16539 -10448
rect 16595 -10456 16639 -10448
rect 16695 -10456 16739 -10448
rect 9239 -10500 9247 -10456
rect 9339 -10500 9347 -10456
rect 9439 -10500 9447 -10456
rect 9539 -10500 9547 -10456
rect 9639 -10500 9647 -10456
rect 9739 -10500 9747 -10456
rect 9839 -10500 9847 -10456
rect 9939 -10500 9947 -10456
rect 10039 -10500 10047 -10456
rect 10139 -10500 10147 -10456
rect 10239 -10500 10247 -10456
rect 10339 -10500 10347 -10456
rect 10439 -10500 10447 -10456
rect 10539 -10500 10547 -10456
rect 10639 -10500 10647 -10456
rect 10739 -10500 10747 -10456
rect 11239 -10500 11247 -10456
rect 11339 -10500 11347 -10456
rect 11439 -10500 11447 -10456
rect 11539 -10500 11547 -10456
rect 11639 -10500 11647 -10456
rect 11739 -10500 11747 -10456
rect 11839 -10500 11847 -10456
rect 11939 -10500 11947 -10456
rect 12039 -10500 12047 -10456
rect 12139 -10500 12147 -10456
rect 12239 -10500 12247 -10456
rect 12339 -10500 12347 -10456
rect 12439 -10500 12447 -10456
rect 12539 -10500 12547 -10456
rect 12639 -10500 12647 -10456
rect 12739 -10500 12747 -10456
rect 13239 -10500 13247 -10456
rect 13339 -10500 13347 -10456
rect 13439 -10500 13447 -10456
rect 13539 -10500 13547 -10456
rect 13639 -10500 13647 -10456
rect 13739 -10500 13747 -10456
rect 13839 -10500 13847 -10456
rect 13939 -10500 13947 -10456
rect 14039 -10500 14047 -10456
rect 14139 -10500 14147 -10456
rect 14239 -10500 14247 -10456
rect 14339 -10500 14347 -10456
rect 14439 -10500 14447 -10456
rect 14539 -10500 14547 -10456
rect 14639 -10500 14647 -10456
rect 14739 -10500 14747 -10456
rect 15239 -10500 15247 -10456
rect 15339 -10500 15347 -10456
rect 15439 -10500 15447 -10456
rect 15539 -10500 15547 -10456
rect 15639 -10500 15647 -10456
rect 15739 -10500 15747 -10456
rect 15839 -10500 15847 -10456
rect 15939 -10500 15947 -10456
rect 16039 -10500 16047 -10456
rect 16139 -10500 16147 -10456
rect 16239 -10500 16247 -10456
rect 16339 -10500 16347 -10456
rect 16439 -10500 16447 -10456
rect 16539 -10500 16547 -10456
rect 16639 -10500 16647 -10456
rect 16739 -10500 16747 -10456
rect 37267 -10482 37275 -10438
rect 37367 -10482 37375 -10438
rect 37467 -10482 37475 -10438
rect 37567 -10482 37575 -10438
rect 37667 -10482 37675 -10438
rect 37767 -10482 37775 -10438
rect 37867 -10482 37875 -10438
rect 37967 -10482 37975 -10438
rect 38067 -10482 38075 -10438
rect 38167 -10482 38175 -10438
rect 38267 -10482 38275 -10438
rect 38367 -10482 38375 -10438
rect 38467 -10482 38475 -10438
rect 38567 -10482 38575 -10438
rect 38667 -10482 38675 -10438
rect 38767 -10482 38775 -10438
rect 39267 -10482 39275 -10438
rect 39367 -10482 39375 -10438
rect 39467 -10482 39475 -10438
rect 39567 -10482 39575 -10438
rect 39667 -10482 39675 -10438
rect 39767 -10482 39775 -10438
rect 39867 -10482 39875 -10438
rect 39967 -10482 39975 -10438
rect 40067 -10482 40075 -10438
rect 40167 -10482 40175 -10438
rect 40267 -10482 40275 -10438
rect 40367 -10482 40375 -10438
rect 40467 -10482 40475 -10438
rect 40567 -10482 40575 -10438
rect 40667 -10482 40675 -10438
rect 40767 -10482 40775 -10438
rect 41267 -10482 41275 -10438
rect 41367 -10482 41375 -10438
rect 41467 -10482 41475 -10438
rect 41567 -10482 41575 -10438
rect 41667 -10482 41675 -10438
rect 41767 -10482 41775 -10438
rect 41867 -10482 41875 -10438
rect 41967 -10482 41975 -10438
rect 42067 -10482 42075 -10438
rect 42167 -10482 42175 -10438
rect 42267 -10482 42275 -10438
rect 42367 -10482 42375 -10438
rect 42467 -10482 42475 -10438
rect 42567 -10482 42575 -10438
rect 42667 -10482 42675 -10438
rect 42767 -10482 42775 -10438
rect 43267 -10482 43275 -10438
rect 43367 -10482 43375 -10438
rect 43467 -10482 43475 -10438
rect 43567 -10482 43575 -10438
rect 43667 -10482 43675 -10438
rect 43767 -10482 43775 -10438
rect 43867 -10482 43875 -10438
rect 43967 -10482 43975 -10438
rect 44067 -10482 44075 -10438
rect 44167 -10482 44175 -10438
rect 44267 -10482 44275 -10438
rect 44367 -10482 44375 -10438
rect 44467 -10482 44475 -10438
rect 44567 -10482 44575 -10438
rect 44667 -10482 44675 -10438
rect 44767 -10482 44775 -10438
rect 37223 -10538 37267 -10530
rect 37323 -10538 37367 -10530
rect 37423 -10538 37467 -10530
rect 37523 -10538 37567 -10530
rect 37623 -10538 37667 -10530
rect 37723 -10538 37767 -10530
rect 37823 -10538 37867 -10530
rect 37923 -10538 37967 -10530
rect 38023 -10538 38067 -10530
rect 38123 -10538 38167 -10530
rect 38223 -10538 38267 -10530
rect 38323 -10538 38367 -10530
rect 38423 -10538 38467 -10530
rect 38523 -10538 38567 -10530
rect 38623 -10538 38667 -10530
rect 38723 -10538 38767 -10530
rect 39223 -10538 39267 -10530
rect 39323 -10538 39367 -10530
rect 39423 -10538 39467 -10530
rect 39523 -10538 39567 -10530
rect 39623 -10538 39667 -10530
rect 39723 -10538 39767 -10530
rect 39823 -10538 39867 -10530
rect 39923 -10538 39967 -10530
rect 40023 -10538 40067 -10530
rect 40123 -10538 40167 -10530
rect 40223 -10538 40267 -10530
rect 40323 -10538 40367 -10530
rect 40423 -10538 40467 -10530
rect 40523 -10538 40567 -10530
rect 40623 -10538 40667 -10530
rect 40723 -10538 40767 -10530
rect 41223 -10538 41267 -10530
rect 41323 -10538 41367 -10530
rect 41423 -10538 41467 -10530
rect 41523 -10538 41567 -10530
rect 41623 -10538 41667 -10530
rect 41723 -10538 41767 -10530
rect 41823 -10538 41867 -10530
rect 41923 -10538 41967 -10530
rect 42023 -10538 42067 -10530
rect 42123 -10538 42167 -10530
rect 42223 -10538 42267 -10530
rect 42323 -10538 42367 -10530
rect 42423 -10538 42467 -10530
rect 42523 -10538 42567 -10530
rect 42623 -10538 42667 -10530
rect 42723 -10538 42767 -10530
rect 43223 -10538 43267 -10530
rect 43323 -10538 43367 -10530
rect 43423 -10538 43467 -10530
rect 43523 -10538 43567 -10530
rect 43623 -10538 43667 -10530
rect 43723 -10538 43767 -10530
rect 43823 -10538 43867 -10530
rect 43923 -10538 43967 -10530
rect 44023 -10538 44067 -10530
rect 44123 -10538 44167 -10530
rect 44223 -10538 44267 -10530
rect 44323 -10538 44367 -10530
rect 44423 -10538 44467 -10530
rect 44523 -10538 44567 -10530
rect 44623 -10538 44667 -10530
rect 44723 -10538 44767 -10530
rect 9195 -10556 9239 -10548
rect 9295 -10556 9339 -10548
rect 9395 -10556 9439 -10548
rect 9495 -10556 9539 -10548
rect 9595 -10556 9639 -10548
rect 9695 -10556 9739 -10548
rect 9795 -10556 9839 -10548
rect 9895 -10556 9939 -10548
rect 9995 -10556 10039 -10548
rect 10095 -10556 10139 -10548
rect 10195 -10556 10239 -10548
rect 10295 -10556 10339 -10548
rect 10395 -10556 10439 -10548
rect 10495 -10556 10539 -10548
rect 10595 -10556 10639 -10548
rect 10695 -10556 10739 -10548
rect 11195 -10556 11239 -10548
rect 11295 -10556 11339 -10548
rect 11395 -10556 11439 -10548
rect 11495 -10556 11539 -10548
rect 11595 -10556 11639 -10548
rect 11695 -10556 11739 -10548
rect 11795 -10556 11839 -10548
rect 11895 -10556 11939 -10548
rect 11995 -10556 12039 -10548
rect 12095 -10556 12139 -10548
rect 12195 -10556 12239 -10548
rect 12295 -10556 12339 -10548
rect 12395 -10556 12439 -10548
rect 12495 -10556 12539 -10548
rect 12595 -10556 12639 -10548
rect 12695 -10556 12739 -10548
rect 13195 -10556 13239 -10548
rect 13295 -10556 13339 -10548
rect 13395 -10556 13439 -10548
rect 13495 -10556 13539 -10548
rect 13595 -10556 13639 -10548
rect 13695 -10556 13739 -10548
rect 13795 -10556 13839 -10548
rect 13895 -10556 13939 -10548
rect 13995 -10556 14039 -10548
rect 14095 -10556 14139 -10548
rect 14195 -10556 14239 -10548
rect 14295 -10556 14339 -10548
rect 14395 -10556 14439 -10548
rect 14495 -10556 14539 -10548
rect 14595 -10556 14639 -10548
rect 14695 -10556 14739 -10548
rect 15195 -10556 15239 -10548
rect 15295 -10556 15339 -10548
rect 15395 -10556 15439 -10548
rect 15495 -10556 15539 -10548
rect 15595 -10556 15639 -10548
rect 15695 -10556 15739 -10548
rect 15795 -10556 15839 -10548
rect 15895 -10556 15939 -10548
rect 15995 -10556 16039 -10548
rect 16095 -10556 16139 -10548
rect 16195 -10556 16239 -10548
rect 16295 -10556 16339 -10548
rect 16395 -10556 16439 -10548
rect 16495 -10556 16539 -10548
rect 16595 -10556 16639 -10548
rect 16695 -10556 16739 -10548
rect 9239 -10600 9247 -10556
rect 9339 -10600 9347 -10556
rect 9439 -10600 9447 -10556
rect 9539 -10600 9547 -10556
rect 9639 -10600 9647 -10556
rect 9739 -10600 9747 -10556
rect 9839 -10600 9847 -10556
rect 9939 -10600 9947 -10556
rect 10039 -10600 10047 -10556
rect 10139 -10600 10147 -10556
rect 10239 -10600 10247 -10556
rect 10339 -10600 10347 -10556
rect 10439 -10600 10447 -10556
rect 10539 -10600 10547 -10556
rect 10639 -10600 10647 -10556
rect 10739 -10600 10747 -10556
rect 11239 -10600 11247 -10556
rect 11339 -10600 11347 -10556
rect 11439 -10600 11447 -10556
rect 11539 -10600 11547 -10556
rect 11639 -10600 11647 -10556
rect 11739 -10600 11747 -10556
rect 11839 -10600 11847 -10556
rect 11939 -10600 11947 -10556
rect 12039 -10600 12047 -10556
rect 12139 -10600 12147 -10556
rect 12239 -10600 12247 -10556
rect 12339 -10600 12347 -10556
rect 12439 -10600 12447 -10556
rect 12539 -10600 12547 -10556
rect 12639 -10600 12647 -10556
rect 12739 -10600 12747 -10556
rect 13239 -10600 13247 -10556
rect 13339 -10600 13347 -10556
rect 13439 -10600 13447 -10556
rect 13539 -10600 13547 -10556
rect 13639 -10600 13647 -10556
rect 13739 -10600 13747 -10556
rect 13839 -10600 13847 -10556
rect 13939 -10600 13947 -10556
rect 14039 -10600 14047 -10556
rect 14139 -10600 14147 -10556
rect 14239 -10600 14247 -10556
rect 14339 -10600 14347 -10556
rect 14439 -10600 14447 -10556
rect 14539 -10600 14547 -10556
rect 14639 -10600 14647 -10556
rect 14739 -10600 14747 -10556
rect 15239 -10600 15247 -10556
rect 15339 -10600 15347 -10556
rect 15439 -10600 15447 -10556
rect 15539 -10600 15547 -10556
rect 15639 -10600 15647 -10556
rect 15739 -10600 15747 -10556
rect 15839 -10600 15847 -10556
rect 15939 -10600 15947 -10556
rect 16039 -10600 16047 -10556
rect 16139 -10600 16147 -10556
rect 16239 -10600 16247 -10556
rect 16339 -10600 16347 -10556
rect 16439 -10600 16447 -10556
rect 16539 -10600 16547 -10556
rect 16639 -10600 16647 -10556
rect 16739 -10600 16747 -10556
rect 37267 -10582 37275 -10538
rect 37367 -10582 37375 -10538
rect 37467 -10582 37475 -10538
rect 37567 -10582 37575 -10538
rect 37667 -10582 37675 -10538
rect 37767 -10582 37775 -10538
rect 37867 -10582 37875 -10538
rect 37967 -10582 37975 -10538
rect 38067 -10582 38075 -10538
rect 38167 -10582 38175 -10538
rect 38267 -10582 38275 -10538
rect 38367 -10582 38375 -10538
rect 38467 -10582 38475 -10538
rect 38567 -10582 38575 -10538
rect 38667 -10582 38675 -10538
rect 38767 -10582 38775 -10538
rect 39267 -10582 39275 -10538
rect 39367 -10582 39375 -10538
rect 39467 -10582 39475 -10538
rect 39567 -10582 39575 -10538
rect 39667 -10582 39675 -10538
rect 39767 -10582 39775 -10538
rect 39867 -10582 39875 -10538
rect 39967 -10582 39975 -10538
rect 40067 -10582 40075 -10538
rect 40167 -10582 40175 -10538
rect 40267 -10582 40275 -10538
rect 40367 -10582 40375 -10538
rect 40467 -10582 40475 -10538
rect 40567 -10582 40575 -10538
rect 40667 -10582 40675 -10538
rect 40767 -10582 40775 -10538
rect 41267 -10582 41275 -10538
rect 41367 -10582 41375 -10538
rect 41467 -10582 41475 -10538
rect 41567 -10582 41575 -10538
rect 41667 -10582 41675 -10538
rect 41767 -10582 41775 -10538
rect 41867 -10582 41875 -10538
rect 41967 -10582 41975 -10538
rect 42067 -10582 42075 -10538
rect 42167 -10582 42175 -10538
rect 42267 -10582 42275 -10538
rect 42367 -10582 42375 -10538
rect 42467 -10582 42475 -10538
rect 42567 -10582 42575 -10538
rect 42667 -10582 42675 -10538
rect 42767 -10582 42775 -10538
rect 43267 -10582 43275 -10538
rect 43367 -10582 43375 -10538
rect 43467 -10582 43475 -10538
rect 43567 -10582 43575 -10538
rect 43667 -10582 43675 -10538
rect 43767 -10582 43775 -10538
rect 43867 -10582 43875 -10538
rect 43967 -10582 43975 -10538
rect 44067 -10582 44075 -10538
rect 44167 -10582 44175 -10538
rect 44267 -10582 44275 -10538
rect 44367 -10582 44375 -10538
rect 44467 -10582 44475 -10538
rect 44567 -10582 44575 -10538
rect 44667 -10582 44675 -10538
rect 44767 -10582 44775 -10538
rect 37223 -10638 37267 -10630
rect 37323 -10638 37367 -10630
rect 37423 -10638 37467 -10630
rect 37523 -10638 37567 -10630
rect 37623 -10638 37667 -10630
rect 37723 -10638 37767 -10630
rect 37823 -10638 37867 -10630
rect 37923 -10638 37967 -10630
rect 38023 -10638 38067 -10630
rect 38123 -10638 38167 -10630
rect 38223 -10638 38267 -10630
rect 38323 -10638 38367 -10630
rect 38423 -10638 38467 -10630
rect 38523 -10638 38567 -10630
rect 38623 -10638 38667 -10630
rect 38723 -10638 38767 -10630
rect 39223 -10638 39267 -10630
rect 39323 -10638 39367 -10630
rect 39423 -10638 39467 -10630
rect 39523 -10638 39567 -10630
rect 39623 -10638 39667 -10630
rect 39723 -10638 39767 -10630
rect 39823 -10638 39867 -10630
rect 39923 -10638 39967 -10630
rect 40023 -10638 40067 -10630
rect 40123 -10638 40167 -10630
rect 40223 -10638 40267 -10630
rect 40323 -10638 40367 -10630
rect 40423 -10638 40467 -10630
rect 40523 -10638 40567 -10630
rect 40623 -10638 40667 -10630
rect 40723 -10638 40767 -10630
rect 41223 -10638 41267 -10630
rect 41323 -10638 41367 -10630
rect 41423 -10638 41467 -10630
rect 41523 -10638 41567 -10630
rect 41623 -10638 41667 -10630
rect 41723 -10638 41767 -10630
rect 41823 -10638 41867 -10630
rect 41923 -10638 41967 -10630
rect 42023 -10638 42067 -10630
rect 42123 -10638 42167 -10630
rect 42223 -10638 42267 -10630
rect 42323 -10638 42367 -10630
rect 42423 -10638 42467 -10630
rect 42523 -10638 42567 -10630
rect 42623 -10638 42667 -10630
rect 42723 -10638 42767 -10630
rect 43223 -10638 43267 -10630
rect 43323 -10638 43367 -10630
rect 43423 -10638 43467 -10630
rect 43523 -10638 43567 -10630
rect 43623 -10638 43667 -10630
rect 43723 -10638 43767 -10630
rect 43823 -10638 43867 -10630
rect 43923 -10638 43967 -10630
rect 44023 -10638 44067 -10630
rect 44123 -10638 44167 -10630
rect 44223 -10638 44267 -10630
rect 44323 -10638 44367 -10630
rect 44423 -10638 44467 -10630
rect 44523 -10638 44567 -10630
rect 44623 -10638 44667 -10630
rect 44723 -10638 44767 -10630
rect 9195 -10656 9239 -10648
rect 9295 -10656 9339 -10648
rect 9395 -10656 9439 -10648
rect 9495 -10656 9539 -10648
rect 9595 -10656 9639 -10648
rect 9695 -10656 9739 -10648
rect 9795 -10656 9839 -10648
rect 9895 -10656 9939 -10648
rect 9995 -10656 10039 -10648
rect 10095 -10656 10139 -10648
rect 10195 -10656 10239 -10648
rect 10295 -10656 10339 -10648
rect 10395 -10656 10439 -10648
rect 10495 -10656 10539 -10648
rect 10595 -10656 10639 -10648
rect 10695 -10656 10739 -10648
rect 11195 -10656 11239 -10648
rect 11295 -10656 11339 -10648
rect 11395 -10656 11439 -10648
rect 11495 -10656 11539 -10648
rect 11595 -10656 11639 -10648
rect 11695 -10656 11739 -10648
rect 11795 -10656 11839 -10648
rect 11895 -10656 11939 -10648
rect 11995 -10656 12039 -10648
rect 12095 -10656 12139 -10648
rect 12195 -10656 12239 -10648
rect 12295 -10656 12339 -10648
rect 12395 -10656 12439 -10648
rect 12495 -10656 12539 -10648
rect 12595 -10656 12639 -10648
rect 12695 -10656 12739 -10648
rect 13195 -10656 13239 -10648
rect 13295 -10656 13339 -10648
rect 13395 -10656 13439 -10648
rect 13495 -10656 13539 -10648
rect 13595 -10656 13639 -10648
rect 13695 -10656 13739 -10648
rect 13795 -10656 13839 -10648
rect 13895 -10656 13939 -10648
rect 13995 -10656 14039 -10648
rect 14095 -10656 14139 -10648
rect 14195 -10656 14239 -10648
rect 14295 -10656 14339 -10648
rect 14395 -10656 14439 -10648
rect 14495 -10656 14539 -10648
rect 14595 -10656 14639 -10648
rect 14695 -10656 14739 -10648
rect 15195 -10656 15239 -10648
rect 15295 -10656 15339 -10648
rect 15395 -10656 15439 -10648
rect 15495 -10656 15539 -10648
rect 15595 -10656 15639 -10648
rect 15695 -10656 15739 -10648
rect 15795 -10656 15839 -10648
rect 15895 -10656 15939 -10648
rect 15995 -10656 16039 -10648
rect 16095 -10656 16139 -10648
rect 16195 -10656 16239 -10648
rect 16295 -10656 16339 -10648
rect 16395 -10656 16439 -10648
rect 16495 -10656 16539 -10648
rect 16595 -10656 16639 -10648
rect 16695 -10656 16739 -10648
rect 9239 -10700 9247 -10656
rect 9339 -10700 9347 -10656
rect 9439 -10700 9447 -10656
rect 9539 -10700 9547 -10656
rect 9639 -10700 9647 -10656
rect 9739 -10700 9747 -10656
rect 9839 -10700 9847 -10656
rect 9939 -10700 9947 -10656
rect 10039 -10700 10047 -10656
rect 10139 -10700 10147 -10656
rect 10239 -10700 10247 -10656
rect 10339 -10700 10347 -10656
rect 10439 -10700 10447 -10656
rect 10539 -10700 10547 -10656
rect 10639 -10700 10647 -10656
rect 10739 -10700 10747 -10656
rect 11239 -10700 11247 -10656
rect 11339 -10700 11347 -10656
rect 11439 -10700 11447 -10656
rect 11539 -10700 11547 -10656
rect 11639 -10700 11647 -10656
rect 11739 -10700 11747 -10656
rect 11839 -10700 11847 -10656
rect 11939 -10700 11947 -10656
rect 12039 -10700 12047 -10656
rect 12139 -10700 12147 -10656
rect 12239 -10700 12247 -10656
rect 12339 -10700 12347 -10656
rect 12439 -10700 12447 -10656
rect 12539 -10700 12547 -10656
rect 12639 -10700 12647 -10656
rect 12739 -10700 12747 -10656
rect 13239 -10700 13247 -10656
rect 13339 -10700 13347 -10656
rect 13439 -10700 13447 -10656
rect 13539 -10700 13547 -10656
rect 13639 -10700 13647 -10656
rect 13739 -10700 13747 -10656
rect 13839 -10700 13847 -10656
rect 13939 -10700 13947 -10656
rect 14039 -10700 14047 -10656
rect 14139 -10700 14147 -10656
rect 14239 -10700 14247 -10656
rect 14339 -10700 14347 -10656
rect 14439 -10700 14447 -10656
rect 14539 -10700 14547 -10656
rect 14639 -10700 14647 -10656
rect 14739 -10700 14747 -10656
rect 15239 -10700 15247 -10656
rect 15339 -10700 15347 -10656
rect 15439 -10700 15447 -10656
rect 15539 -10700 15547 -10656
rect 15639 -10700 15647 -10656
rect 15739 -10700 15747 -10656
rect 15839 -10700 15847 -10656
rect 15939 -10700 15947 -10656
rect 16039 -10700 16047 -10656
rect 16139 -10700 16147 -10656
rect 16239 -10700 16247 -10656
rect 16339 -10700 16347 -10656
rect 16439 -10700 16447 -10656
rect 16539 -10700 16547 -10656
rect 16639 -10700 16647 -10656
rect 16739 -10700 16747 -10656
rect 37267 -10682 37275 -10638
rect 37367 -10682 37375 -10638
rect 37467 -10682 37475 -10638
rect 37567 -10682 37575 -10638
rect 37667 -10682 37675 -10638
rect 37767 -10682 37775 -10638
rect 37867 -10682 37875 -10638
rect 37967 -10682 37975 -10638
rect 38067 -10682 38075 -10638
rect 38167 -10682 38175 -10638
rect 38267 -10682 38275 -10638
rect 38367 -10682 38375 -10638
rect 38467 -10682 38475 -10638
rect 38567 -10682 38575 -10638
rect 38667 -10682 38675 -10638
rect 38767 -10682 38775 -10638
rect 39267 -10682 39275 -10638
rect 39367 -10682 39375 -10638
rect 39467 -10682 39475 -10638
rect 39567 -10682 39575 -10638
rect 39667 -10682 39675 -10638
rect 39767 -10682 39775 -10638
rect 39867 -10682 39875 -10638
rect 39967 -10682 39975 -10638
rect 40067 -10682 40075 -10638
rect 40167 -10682 40175 -10638
rect 40267 -10682 40275 -10638
rect 40367 -10682 40375 -10638
rect 40467 -10682 40475 -10638
rect 40567 -10682 40575 -10638
rect 40667 -10682 40675 -10638
rect 40767 -10682 40775 -10638
rect 41267 -10682 41275 -10638
rect 41367 -10682 41375 -10638
rect 41467 -10682 41475 -10638
rect 41567 -10682 41575 -10638
rect 41667 -10682 41675 -10638
rect 41767 -10682 41775 -10638
rect 41867 -10682 41875 -10638
rect 41967 -10682 41975 -10638
rect 42067 -10682 42075 -10638
rect 42167 -10682 42175 -10638
rect 42267 -10682 42275 -10638
rect 42367 -10682 42375 -10638
rect 42467 -10682 42475 -10638
rect 42567 -10682 42575 -10638
rect 42667 -10682 42675 -10638
rect 42767 -10682 42775 -10638
rect 43267 -10682 43275 -10638
rect 43367 -10682 43375 -10638
rect 43467 -10682 43475 -10638
rect 43567 -10682 43575 -10638
rect 43667 -10682 43675 -10638
rect 43767 -10682 43775 -10638
rect 43867 -10682 43875 -10638
rect 43967 -10682 43975 -10638
rect 44067 -10682 44075 -10638
rect 44167 -10682 44175 -10638
rect 44267 -10682 44275 -10638
rect 44367 -10682 44375 -10638
rect 44467 -10682 44475 -10638
rect 44567 -10682 44575 -10638
rect 44667 -10682 44675 -10638
rect 44767 -10682 44775 -10638
rect 37223 -10738 37267 -10730
rect 37323 -10738 37367 -10730
rect 37423 -10738 37467 -10730
rect 37523 -10738 37567 -10730
rect 37623 -10738 37667 -10730
rect 37723 -10738 37767 -10730
rect 37823 -10738 37867 -10730
rect 37923 -10738 37967 -10730
rect 38023 -10738 38067 -10730
rect 38123 -10738 38167 -10730
rect 38223 -10738 38267 -10730
rect 38323 -10738 38367 -10730
rect 38423 -10738 38467 -10730
rect 38523 -10738 38567 -10730
rect 38623 -10738 38667 -10730
rect 38723 -10738 38767 -10730
rect 39223 -10738 39267 -10730
rect 39323 -10738 39367 -10730
rect 39423 -10738 39467 -10730
rect 39523 -10738 39567 -10730
rect 39623 -10738 39667 -10730
rect 39723 -10738 39767 -10730
rect 39823 -10738 39867 -10730
rect 39923 -10738 39967 -10730
rect 40023 -10738 40067 -10730
rect 40123 -10738 40167 -10730
rect 40223 -10738 40267 -10730
rect 40323 -10738 40367 -10730
rect 40423 -10738 40467 -10730
rect 40523 -10738 40567 -10730
rect 40623 -10738 40667 -10730
rect 40723 -10738 40767 -10730
rect 41223 -10738 41267 -10730
rect 41323 -10738 41367 -10730
rect 41423 -10738 41467 -10730
rect 41523 -10738 41567 -10730
rect 41623 -10738 41667 -10730
rect 41723 -10738 41767 -10730
rect 41823 -10738 41867 -10730
rect 41923 -10738 41967 -10730
rect 42023 -10738 42067 -10730
rect 42123 -10738 42167 -10730
rect 42223 -10738 42267 -10730
rect 42323 -10738 42367 -10730
rect 42423 -10738 42467 -10730
rect 42523 -10738 42567 -10730
rect 42623 -10738 42667 -10730
rect 42723 -10738 42767 -10730
rect 43223 -10738 43267 -10730
rect 43323 -10738 43367 -10730
rect 43423 -10738 43467 -10730
rect 43523 -10738 43567 -10730
rect 43623 -10738 43667 -10730
rect 43723 -10738 43767 -10730
rect 43823 -10738 43867 -10730
rect 43923 -10738 43967 -10730
rect 44023 -10738 44067 -10730
rect 44123 -10738 44167 -10730
rect 44223 -10738 44267 -10730
rect 44323 -10738 44367 -10730
rect 44423 -10738 44467 -10730
rect 44523 -10738 44567 -10730
rect 44623 -10738 44667 -10730
rect 44723 -10738 44767 -10730
rect 9195 -10756 9239 -10748
rect 9295 -10756 9339 -10748
rect 9395 -10756 9439 -10748
rect 9495 -10756 9539 -10748
rect 9595 -10756 9639 -10748
rect 9695 -10756 9739 -10748
rect 9795 -10756 9839 -10748
rect 9895 -10756 9939 -10748
rect 9995 -10756 10039 -10748
rect 10095 -10756 10139 -10748
rect 10195 -10756 10239 -10748
rect 10295 -10756 10339 -10748
rect 10395 -10756 10439 -10748
rect 10495 -10756 10539 -10748
rect 10595 -10756 10639 -10748
rect 10695 -10756 10739 -10748
rect 11195 -10756 11239 -10748
rect 11295 -10756 11339 -10748
rect 11395 -10756 11439 -10748
rect 11495 -10756 11539 -10748
rect 11595 -10756 11639 -10748
rect 11695 -10756 11739 -10748
rect 11795 -10756 11839 -10748
rect 11895 -10756 11939 -10748
rect 11995 -10756 12039 -10748
rect 12095 -10756 12139 -10748
rect 12195 -10756 12239 -10748
rect 12295 -10756 12339 -10748
rect 12395 -10756 12439 -10748
rect 12495 -10756 12539 -10748
rect 12595 -10756 12639 -10748
rect 12695 -10756 12739 -10748
rect 13195 -10756 13239 -10748
rect 13295 -10756 13339 -10748
rect 13395 -10756 13439 -10748
rect 13495 -10756 13539 -10748
rect 13595 -10756 13639 -10748
rect 13695 -10756 13739 -10748
rect 13795 -10756 13839 -10748
rect 13895 -10756 13939 -10748
rect 13995 -10756 14039 -10748
rect 14095 -10756 14139 -10748
rect 14195 -10756 14239 -10748
rect 14295 -10756 14339 -10748
rect 14395 -10756 14439 -10748
rect 14495 -10756 14539 -10748
rect 14595 -10756 14639 -10748
rect 14695 -10756 14739 -10748
rect 15195 -10756 15239 -10748
rect 15295 -10756 15339 -10748
rect 15395 -10756 15439 -10748
rect 15495 -10756 15539 -10748
rect 15595 -10756 15639 -10748
rect 15695 -10756 15739 -10748
rect 15795 -10756 15839 -10748
rect 15895 -10756 15939 -10748
rect 15995 -10756 16039 -10748
rect 16095 -10756 16139 -10748
rect 16195 -10756 16239 -10748
rect 16295 -10756 16339 -10748
rect 16395 -10756 16439 -10748
rect 16495 -10756 16539 -10748
rect 16595 -10756 16639 -10748
rect 16695 -10756 16739 -10748
rect 9239 -10800 9247 -10756
rect 9339 -10800 9347 -10756
rect 9439 -10800 9447 -10756
rect 9539 -10800 9547 -10756
rect 9639 -10800 9647 -10756
rect 9739 -10800 9747 -10756
rect 9839 -10800 9847 -10756
rect 9939 -10800 9947 -10756
rect 10039 -10800 10047 -10756
rect 10139 -10800 10147 -10756
rect 10239 -10800 10247 -10756
rect 10339 -10800 10347 -10756
rect 10439 -10800 10447 -10756
rect 10539 -10800 10547 -10756
rect 10639 -10800 10647 -10756
rect 10739 -10800 10747 -10756
rect 11239 -10800 11247 -10756
rect 11339 -10800 11347 -10756
rect 11439 -10800 11447 -10756
rect 11539 -10800 11547 -10756
rect 11639 -10800 11647 -10756
rect 11739 -10800 11747 -10756
rect 11839 -10800 11847 -10756
rect 11939 -10800 11947 -10756
rect 12039 -10800 12047 -10756
rect 12139 -10800 12147 -10756
rect 12239 -10800 12247 -10756
rect 12339 -10800 12347 -10756
rect 12439 -10800 12447 -10756
rect 12539 -10800 12547 -10756
rect 12639 -10800 12647 -10756
rect 12739 -10800 12747 -10756
rect 13239 -10800 13247 -10756
rect 13339 -10800 13347 -10756
rect 13439 -10800 13447 -10756
rect 13539 -10800 13547 -10756
rect 13639 -10800 13647 -10756
rect 13739 -10800 13747 -10756
rect 13839 -10800 13847 -10756
rect 13939 -10800 13947 -10756
rect 14039 -10800 14047 -10756
rect 14139 -10800 14147 -10756
rect 14239 -10800 14247 -10756
rect 14339 -10800 14347 -10756
rect 14439 -10800 14447 -10756
rect 14539 -10800 14547 -10756
rect 14639 -10800 14647 -10756
rect 14739 -10800 14747 -10756
rect 15239 -10800 15247 -10756
rect 15339 -10800 15347 -10756
rect 15439 -10800 15447 -10756
rect 15539 -10800 15547 -10756
rect 15639 -10800 15647 -10756
rect 15739 -10800 15747 -10756
rect 15839 -10800 15847 -10756
rect 15939 -10800 15947 -10756
rect 16039 -10800 16047 -10756
rect 16139 -10800 16147 -10756
rect 16239 -10800 16247 -10756
rect 16339 -10800 16347 -10756
rect 16439 -10800 16447 -10756
rect 16539 -10800 16547 -10756
rect 16639 -10800 16647 -10756
rect 16739 -10800 16747 -10756
rect 37267 -10782 37275 -10738
rect 37367 -10782 37375 -10738
rect 37467 -10782 37475 -10738
rect 37567 -10782 37575 -10738
rect 37667 -10782 37675 -10738
rect 37767 -10782 37775 -10738
rect 37867 -10782 37875 -10738
rect 37967 -10782 37975 -10738
rect 38067 -10782 38075 -10738
rect 38167 -10782 38175 -10738
rect 38267 -10782 38275 -10738
rect 38367 -10782 38375 -10738
rect 38467 -10782 38475 -10738
rect 38567 -10782 38575 -10738
rect 38667 -10782 38675 -10738
rect 38767 -10782 38775 -10738
rect 39267 -10782 39275 -10738
rect 39367 -10782 39375 -10738
rect 39467 -10782 39475 -10738
rect 39567 -10782 39575 -10738
rect 39667 -10782 39675 -10738
rect 39767 -10782 39775 -10738
rect 39867 -10782 39875 -10738
rect 39967 -10782 39975 -10738
rect 40067 -10782 40075 -10738
rect 40167 -10782 40175 -10738
rect 40267 -10782 40275 -10738
rect 40367 -10782 40375 -10738
rect 40467 -10782 40475 -10738
rect 40567 -10782 40575 -10738
rect 40667 -10782 40675 -10738
rect 40767 -10782 40775 -10738
rect 41267 -10782 41275 -10738
rect 41367 -10782 41375 -10738
rect 41467 -10782 41475 -10738
rect 41567 -10782 41575 -10738
rect 41667 -10782 41675 -10738
rect 41767 -10782 41775 -10738
rect 41867 -10782 41875 -10738
rect 41967 -10782 41975 -10738
rect 42067 -10782 42075 -10738
rect 42167 -10782 42175 -10738
rect 42267 -10782 42275 -10738
rect 42367 -10782 42375 -10738
rect 42467 -10782 42475 -10738
rect 42567 -10782 42575 -10738
rect 42667 -10782 42675 -10738
rect 42767 -10782 42775 -10738
rect 43267 -10782 43275 -10738
rect 43367 -10782 43375 -10738
rect 43467 -10782 43475 -10738
rect 43567 -10782 43575 -10738
rect 43667 -10782 43675 -10738
rect 43767 -10782 43775 -10738
rect 43867 -10782 43875 -10738
rect 43967 -10782 43975 -10738
rect 44067 -10782 44075 -10738
rect 44167 -10782 44175 -10738
rect 44267 -10782 44275 -10738
rect 44367 -10782 44375 -10738
rect 44467 -10782 44475 -10738
rect 44567 -10782 44575 -10738
rect 44667 -10782 44675 -10738
rect 44767 -10782 44775 -10738
rect 37223 -10838 37267 -10830
rect 37323 -10838 37367 -10830
rect 37423 -10838 37467 -10830
rect 37523 -10838 37567 -10830
rect 37623 -10838 37667 -10830
rect 37723 -10838 37767 -10830
rect 37823 -10838 37867 -10830
rect 37923 -10838 37967 -10830
rect 38023 -10838 38067 -10830
rect 38123 -10838 38167 -10830
rect 38223 -10838 38267 -10830
rect 38323 -10838 38367 -10830
rect 38423 -10838 38467 -10830
rect 38523 -10838 38567 -10830
rect 38623 -10838 38667 -10830
rect 38723 -10838 38767 -10830
rect 39223 -10838 39267 -10830
rect 39323 -10838 39367 -10830
rect 39423 -10838 39467 -10830
rect 39523 -10838 39567 -10830
rect 39623 -10838 39667 -10830
rect 39723 -10838 39767 -10830
rect 39823 -10838 39867 -10830
rect 39923 -10838 39967 -10830
rect 40023 -10838 40067 -10830
rect 40123 -10838 40167 -10830
rect 40223 -10838 40267 -10830
rect 40323 -10838 40367 -10830
rect 40423 -10838 40467 -10830
rect 40523 -10838 40567 -10830
rect 40623 -10838 40667 -10830
rect 40723 -10838 40767 -10830
rect 41223 -10838 41267 -10830
rect 41323 -10838 41367 -10830
rect 41423 -10838 41467 -10830
rect 41523 -10838 41567 -10830
rect 41623 -10838 41667 -10830
rect 41723 -10838 41767 -10830
rect 41823 -10838 41867 -10830
rect 41923 -10838 41967 -10830
rect 42023 -10838 42067 -10830
rect 42123 -10838 42167 -10830
rect 42223 -10838 42267 -10830
rect 42323 -10838 42367 -10830
rect 42423 -10838 42467 -10830
rect 42523 -10838 42567 -10830
rect 42623 -10838 42667 -10830
rect 42723 -10838 42767 -10830
rect 43223 -10838 43267 -10830
rect 43323 -10838 43367 -10830
rect 43423 -10838 43467 -10830
rect 43523 -10838 43567 -10830
rect 43623 -10838 43667 -10830
rect 43723 -10838 43767 -10830
rect 43823 -10838 43867 -10830
rect 43923 -10838 43967 -10830
rect 44023 -10838 44067 -10830
rect 44123 -10838 44167 -10830
rect 44223 -10838 44267 -10830
rect 44323 -10838 44367 -10830
rect 44423 -10838 44467 -10830
rect 44523 -10838 44567 -10830
rect 44623 -10838 44667 -10830
rect 44723 -10838 44767 -10830
rect 9195 -10856 9239 -10848
rect 9295 -10856 9339 -10848
rect 9395 -10856 9439 -10848
rect 9495 -10856 9539 -10848
rect 9595 -10856 9639 -10848
rect 9695 -10856 9739 -10848
rect 9795 -10856 9839 -10848
rect 9895 -10856 9939 -10848
rect 9995 -10856 10039 -10848
rect 10095 -10856 10139 -10848
rect 10195 -10856 10239 -10848
rect 10295 -10856 10339 -10848
rect 10395 -10856 10439 -10848
rect 10495 -10856 10539 -10848
rect 10595 -10856 10639 -10848
rect 10695 -10856 10739 -10848
rect 11195 -10856 11239 -10848
rect 11295 -10856 11339 -10848
rect 11395 -10856 11439 -10848
rect 11495 -10856 11539 -10848
rect 11595 -10856 11639 -10848
rect 11695 -10856 11739 -10848
rect 11795 -10856 11839 -10848
rect 11895 -10856 11939 -10848
rect 11995 -10856 12039 -10848
rect 12095 -10856 12139 -10848
rect 12195 -10856 12239 -10848
rect 12295 -10856 12339 -10848
rect 12395 -10856 12439 -10848
rect 12495 -10856 12539 -10848
rect 12595 -10856 12639 -10848
rect 12695 -10856 12739 -10848
rect 13195 -10856 13239 -10848
rect 13295 -10856 13339 -10848
rect 13395 -10856 13439 -10848
rect 13495 -10856 13539 -10848
rect 13595 -10856 13639 -10848
rect 13695 -10856 13739 -10848
rect 13795 -10856 13839 -10848
rect 13895 -10856 13939 -10848
rect 13995 -10856 14039 -10848
rect 14095 -10856 14139 -10848
rect 14195 -10856 14239 -10848
rect 14295 -10856 14339 -10848
rect 14395 -10856 14439 -10848
rect 14495 -10856 14539 -10848
rect 14595 -10856 14639 -10848
rect 14695 -10856 14739 -10848
rect 15195 -10856 15239 -10848
rect 15295 -10856 15339 -10848
rect 15395 -10856 15439 -10848
rect 15495 -10856 15539 -10848
rect 15595 -10856 15639 -10848
rect 15695 -10856 15739 -10848
rect 15795 -10856 15839 -10848
rect 15895 -10856 15939 -10848
rect 15995 -10856 16039 -10848
rect 16095 -10856 16139 -10848
rect 16195 -10856 16239 -10848
rect 16295 -10856 16339 -10848
rect 16395 -10856 16439 -10848
rect 16495 -10856 16539 -10848
rect 16595 -10856 16639 -10848
rect 16695 -10856 16739 -10848
rect 9239 -10900 9247 -10856
rect 9339 -10900 9347 -10856
rect 9439 -10900 9447 -10856
rect 9539 -10900 9547 -10856
rect 9639 -10900 9647 -10856
rect 9739 -10900 9747 -10856
rect 9839 -10900 9847 -10856
rect 9939 -10900 9947 -10856
rect 10039 -10900 10047 -10856
rect 10139 -10900 10147 -10856
rect 10239 -10900 10247 -10856
rect 10339 -10900 10347 -10856
rect 10439 -10900 10447 -10856
rect 10539 -10900 10547 -10856
rect 10639 -10900 10647 -10856
rect 10739 -10900 10747 -10856
rect 11239 -10900 11247 -10856
rect 11339 -10900 11347 -10856
rect 11439 -10900 11447 -10856
rect 11539 -10900 11547 -10856
rect 11639 -10900 11647 -10856
rect 11739 -10900 11747 -10856
rect 11839 -10900 11847 -10856
rect 11939 -10900 11947 -10856
rect 12039 -10900 12047 -10856
rect 12139 -10900 12147 -10856
rect 12239 -10900 12247 -10856
rect 12339 -10900 12347 -10856
rect 12439 -10900 12447 -10856
rect 12539 -10900 12547 -10856
rect 12639 -10900 12647 -10856
rect 12739 -10900 12747 -10856
rect 13239 -10900 13247 -10856
rect 13339 -10900 13347 -10856
rect 13439 -10900 13447 -10856
rect 13539 -10900 13547 -10856
rect 13639 -10900 13647 -10856
rect 13739 -10900 13747 -10856
rect 13839 -10900 13847 -10856
rect 13939 -10900 13947 -10856
rect 14039 -10900 14047 -10856
rect 14139 -10900 14147 -10856
rect 14239 -10900 14247 -10856
rect 14339 -10900 14347 -10856
rect 14439 -10900 14447 -10856
rect 14539 -10900 14547 -10856
rect 14639 -10900 14647 -10856
rect 14739 -10900 14747 -10856
rect 15239 -10900 15247 -10856
rect 15339 -10900 15347 -10856
rect 15439 -10900 15447 -10856
rect 15539 -10900 15547 -10856
rect 15639 -10900 15647 -10856
rect 15739 -10900 15747 -10856
rect 15839 -10900 15847 -10856
rect 15939 -10900 15947 -10856
rect 16039 -10900 16047 -10856
rect 16139 -10900 16147 -10856
rect 16239 -10900 16247 -10856
rect 16339 -10900 16347 -10856
rect 16439 -10900 16447 -10856
rect 16539 -10900 16547 -10856
rect 16639 -10900 16647 -10856
rect 16739 -10900 16747 -10856
rect 37267 -10882 37275 -10838
rect 37367 -10882 37375 -10838
rect 37467 -10882 37475 -10838
rect 37567 -10882 37575 -10838
rect 37667 -10882 37675 -10838
rect 37767 -10882 37775 -10838
rect 37867 -10882 37875 -10838
rect 37967 -10882 37975 -10838
rect 38067 -10882 38075 -10838
rect 38167 -10882 38175 -10838
rect 38267 -10882 38275 -10838
rect 38367 -10882 38375 -10838
rect 38467 -10882 38475 -10838
rect 38567 -10882 38575 -10838
rect 38667 -10882 38675 -10838
rect 38767 -10882 38775 -10838
rect 39267 -10882 39275 -10838
rect 39367 -10882 39375 -10838
rect 39467 -10882 39475 -10838
rect 39567 -10882 39575 -10838
rect 39667 -10882 39675 -10838
rect 39767 -10882 39775 -10838
rect 39867 -10882 39875 -10838
rect 39967 -10882 39975 -10838
rect 40067 -10882 40075 -10838
rect 40167 -10882 40175 -10838
rect 40267 -10882 40275 -10838
rect 40367 -10882 40375 -10838
rect 40467 -10882 40475 -10838
rect 40567 -10882 40575 -10838
rect 40667 -10882 40675 -10838
rect 40767 -10882 40775 -10838
rect 41267 -10882 41275 -10838
rect 41367 -10882 41375 -10838
rect 41467 -10882 41475 -10838
rect 41567 -10882 41575 -10838
rect 41667 -10882 41675 -10838
rect 41767 -10882 41775 -10838
rect 41867 -10882 41875 -10838
rect 41967 -10882 41975 -10838
rect 42067 -10882 42075 -10838
rect 42167 -10882 42175 -10838
rect 42267 -10882 42275 -10838
rect 42367 -10882 42375 -10838
rect 42467 -10882 42475 -10838
rect 42567 -10882 42575 -10838
rect 42667 -10882 42675 -10838
rect 42767 -10882 42775 -10838
rect 43267 -10882 43275 -10838
rect 43367 -10882 43375 -10838
rect 43467 -10882 43475 -10838
rect 43567 -10882 43575 -10838
rect 43667 -10882 43675 -10838
rect 43767 -10882 43775 -10838
rect 43867 -10882 43875 -10838
rect 43967 -10882 43975 -10838
rect 44067 -10882 44075 -10838
rect 44167 -10882 44175 -10838
rect 44267 -10882 44275 -10838
rect 44367 -10882 44375 -10838
rect 44467 -10882 44475 -10838
rect 44567 -10882 44575 -10838
rect 44667 -10882 44675 -10838
rect 44767 -10882 44775 -10838
rect 37223 -10938 37267 -10930
rect 37323 -10938 37367 -10930
rect 37423 -10938 37467 -10930
rect 37523 -10938 37567 -10930
rect 37623 -10938 37667 -10930
rect 37723 -10938 37767 -10930
rect 37823 -10938 37867 -10930
rect 37923 -10938 37967 -10930
rect 38023 -10938 38067 -10930
rect 38123 -10938 38167 -10930
rect 38223 -10938 38267 -10930
rect 38323 -10938 38367 -10930
rect 38423 -10938 38467 -10930
rect 38523 -10938 38567 -10930
rect 38623 -10938 38667 -10930
rect 38723 -10938 38767 -10930
rect 39223 -10938 39267 -10930
rect 39323 -10938 39367 -10930
rect 39423 -10938 39467 -10930
rect 39523 -10938 39567 -10930
rect 39623 -10938 39667 -10930
rect 39723 -10938 39767 -10930
rect 39823 -10938 39867 -10930
rect 39923 -10938 39967 -10930
rect 40023 -10938 40067 -10930
rect 40123 -10938 40167 -10930
rect 40223 -10938 40267 -10930
rect 40323 -10938 40367 -10930
rect 40423 -10938 40467 -10930
rect 40523 -10938 40567 -10930
rect 40623 -10938 40667 -10930
rect 40723 -10938 40767 -10930
rect 41223 -10938 41267 -10930
rect 41323 -10938 41367 -10930
rect 41423 -10938 41467 -10930
rect 41523 -10938 41567 -10930
rect 41623 -10938 41667 -10930
rect 41723 -10938 41767 -10930
rect 41823 -10938 41867 -10930
rect 41923 -10938 41967 -10930
rect 42023 -10938 42067 -10930
rect 42123 -10938 42167 -10930
rect 42223 -10938 42267 -10930
rect 42323 -10938 42367 -10930
rect 42423 -10938 42467 -10930
rect 42523 -10938 42567 -10930
rect 42623 -10938 42667 -10930
rect 42723 -10938 42767 -10930
rect 43223 -10938 43267 -10930
rect 43323 -10938 43367 -10930
rect 43423 -10938 43467 -10930
rect 43523 -10938 43567 -10930
rect 43623 -10938 43667 -10930
rect 43723 -10938 43767 -10930
rect 43823 -10938 43867 -10930
rect 43923 -10938 43967 -10930
rect 44023 -10938 44067 -10930
rect 44123 -10938 44167 -10930
rect 44223 -10938 44267 -10930
rect 44323 -10938 44367 -10930
rect 44423 -10938 44467 -10930
rect 44523 -10938 44567 -10930
rect 44623 -10938 44667 -10930
rect 44723 -10938 44767 -10930
rect 9195 -10956 9239 -10948
rect 9295 -10956 9339 -10948
rect 9395 -10956 9439 -10948
rect 9495 -10956 9539 -10948
rect 9595 -10956 9639 -10948
rect 9695 -10956 9739 -10948
rect 9795 -10956 9839 -10948
rect 9895 -10956 9939 -10948
rect 9995 -10956 10039 -10948
rect 10095 -10956 10139 -10948
rect 10195 -10956 10239 -10948
rect 10295 -10956 10339 -10948
rect 10395 -10956 10439 -10948
rect 10495 -10956 10539 -10948
rect 10595 -10956 10639 -10948
rect 10695 -10956 10739 -10948
rect 11195 -10956 11239 -10948
rect 11295 -10956 11339 -10948
rect 11395 -10956 11439 -10948
rect 11495 -10956 11539 -10948
rect 11595 -10956 11639 -10948
rect 11695 -10956 11739 -10948
rect 11795 -10956 11839 -10948
rect 11895 -10956 11939 -10948
rect 11995 -10956 12039 -10948
rect 12095 -10956 12139 -10948
rect 12195 -10956 12239 -10948
rect 12295 -10956 12339 -10948
rect 12395 -10956 12439 -10948
rect 12495 -10956 12539 -10948
rect 12595 -10956 12639 -10948
rect 12695 -10956 12739 -10948
rect 13195 -10956 13239 -10948
rect 13295 -10956 13339 -10948
rect 13395 -10956 13439 -10948
rect 13495 -10956 13539 -10948
rect 13595 -10956 13639 -10948
rect 13695 -10956 13739 -10948
rect 13795 -10956 13839 -10948
rect 13895 -10956 13939 -10948
rect 13995 -10956 14039 -10948
rect 14095 -10956 14139 -10948
rect 14195 -10956 14239 -10948
rect 14295 -10956 14339 -10948
rect 14395 -10956 14439 -10948
rect 14495 -10956 14539 -10948
rect 14595 -10956 14639 -10948
rect 14695 -10956 14739 -10948
rect 15195 -10956 15239 -10948
rect 15295 -10956 15339 -10948
rect 15395 -10956 15439 -10948
rect 15495 -10956 15539 -10948
rect 15595 -10956 15639 -10948
rect 15695 -10956 15739 -10948
rect 15795 -10956 15839 -10948
rect 15895 -10956 15939 -10948
rect 15995 -10956 16039 -10948
rect 16095 -10956 16139 -10948
rect 16195 -10956 16239 -10948
rect 16295 -10956 16339 -10948
rect 16395 -10956 16439 -10948
rect 16495 -10956 16539 -10948
rect 16595 -10956 16639 -10948
rect 16695 -10956 16739 -10948
rect 9239 -11000 9247 -10956
rect 9339 -11000 9347 -10956
rect 9439 -11000 9447 -10956
rect 9539 -11000 9547 -10956
rect 9639 -11000 9647 -10956
rect 9739 -11000 9747 -10956
rect 9839 -11000 9847 -10956
rect 9939 -11000 9947 -10956
rect 10039 -11000 10047 -10956
rect 10139 -11000 10147 -10956
rect 10239 -11000 10247 -10956
rect 10339 -11000 10347 -10956
rect 10439 -11000 10447 -10956
rect 10539 -11000 10547 -10956
rect 10639 -11000 10647 -10956
rect 10739 -11000 10747 -10956
rect 11239 -11000 11247 -10956
rect 11339 -11000 11347 -10956
rect 11439 -11000 11447 -10956
rect 11539 -11000 11547 -10956
rect 11639 -11000 11647 -10956
rect 11739 -11000 11747 -10956
rect 11839 -11000 11847 -10956
rect 11939 -11000 11947 -10956
rect 12039 -11000 12047 -10956
rect 12139 -11000 12147 -10956
rect 12239 -11000 12247 -10956
rect 12339 -11000 12347 -10956
rect 12439 -11000 12447 -10956
rect 12539 -11000 12547 -10956
rect 12639 -11000 12647 -10956
rect 12739 -11000 12747 -10956
rect 13239 -11000 13247 -10956
rect 13339 -11000 13347 -10956
rect 13439 -11000 13447 -10956
rect 13539 -11000 13547 -10956
rect 13639 -11000 13647 -10956
rect 13739 -11000 13747 -10956
rect 13839 -11000 13847 -10956
rect 13939 -11000 13947 -10956
rect 14039 -11000 14047 -10956
rect 14139 -11000 14147 -10956
rect 14239 -11000 14247 -10956
rect 14339 -11000 14347 -10956
rect 14439 -11000 14447 -10956
rect 14539 -11000 14547 -10956
rect 14639 -11000 14647 -10956
rect 14739 -11000 14747 -10956
rect 15239 -11000 15247 -10956
rect 15339 -11000 15347 -10956
rect 15439 -11000 15447 -10956
rect 15539 -11000 15547 -10956
rect 15639 -11000 15647 -10956
rect 15739 -11000 15747 -10956
rect 15839 -11000 15847 -10956
rect 15939 -11000 15947 -10956
rect 16039 -11000 16047 -10956
rect 16139 -11000 16147 -10956
rect 16239 -11000 16247 -10956
rect 16339 -11000 16347 -10956
rect 16439 -11000 16447 -10956
rect 16539 -11000 16547 -10956
rect 16639 -11000 16647 -10956
rect 16739 -11000 16747 -10956
rect 37267 -10982 37275 -10938
rect 37367 -10982 37375 -10938
rect 37467 -10982 37475 -10938
rect 37567 -10982 37575 -10938
rect 37667 -10982 37675 -10938
rect 37767 -10982 37775 -10938
rect 37867 -10982 37875 -10938
rect 37967 -10982 37975 -10938
rect 38067 -10982 38075 -10938
rect 38167 -10982 38175 -10938
rect 38267 -10982 38275 -10938
rect 38367 -10982 38375 -10938
rect 38467 -10982 38475 -10938
rect 38567 -10982 38575 -10938
rect 38667 -10982 38675 -10938
rect 38767 -10982 38775 -10938
rect 39267 -10982 39275 -10938
rect 39367 -10982 39375 -10938
rect 39467 -10982 39475 -10938
rect 39567 -10982 39575 -10938
rect 39667 -10982 39675 -10938
rect 39767 -10982 39775 -10938
rect 39867 -10982 39875 -10938
rect 39967 -10982 39975 -10938
rect 40067 -10982 40075 -10938
rect 40167 -10982 40175 -10938
rect 40267 -10982 40275 -10938
rect 40367 -10982 40375 -10938
rect 40467 -10982 40475 -10938
rect 40567 -10982 40575 -10938
rect 40667 -10982 40675 -10938
rect 40767 -10982 40775 -10938
rect 41267 -10982 41275 -10938
rect 41367 -10982 41375 -10938
rect 41467 -10982 41475 -10938
rect 41567 -10982 41575 -10938
rect 41667 -10982 41675 -10938
rect 41767 -10982 41775 -10938
rect 41867 -10982 41875 -10938
rect 41967 -10982 41975 -10938
rect 42067 -10982 42075 -10938
rect 42167 -10982 42175 -10938
rect 42267 -10982 42275 -10938
rect 42367 -10982 42375 -10938
rect 42467 -10982 42475 -10938
rect 42567 -10982 42575 -10938
rect 42667 -10982 42675 -10938
rect 42767 -10982 42775 -10938
rect 43267 -10982 43275 -10938
rect 43367 -10982 43375 -10938
rect 43467 -10982 43475 -10938
rect 43567 -10982 43575 -10938
rect 43667 -10982 43675 -10938
rect 43767 -10982 43775 -10938
rect 43867 -10982 43875 -10938
rect 43967 -10982 43975 -10938
rect 44067 -10982 44075 -10938
rect 44167 -10982 44175 -10938
rect 44267 -10982 44275 -10938
rect 44367 -10982 44375 -10938
rect 44467 -10982 44475 -10938
rect 44567 -10982 44575 -10938
rect 44667 -10982 44675 -10938
rect 44767 -10982 44775 -10938
rect 37223 -11038 37267 -11030
rect 37323 -11038 37367 -11030
rect 37423 -11038 37467 -11030
rect 37523 -11038 37567 -11030
rect 37623 -11038 37667 -11030
rect 37723 -11038 37767 -11030
rect 37823 -11038 37867 -11030
rect 37923 -11038 37967 -11030
rect 38023 -11038 38067 -11030
rect 38123 -11038 38167 -11030
rect 38223 -11038 38267 -11030
rect 38323 -11038 38367 -11030
rect 38423 -11038 38467 -11030
rect 38523 -11038 38567 -11030
rect 38623 -11038 38667 -11030
rect 38723 -11038 38767 -11030
rect 39223 -11038 39267 -11030
rect 39323 -11038 39367 -11030
rect 39423 -11038 39467 -11030
rect 39523 -11038 39567 -11030
rect 39623 -11038 39667 -11030
rect 39723 -11038 39767 -11030
rect 39823 -11038 39867 -11030
rect 39923 -11038 39967 -11030
rect 40023 -11038 40067 -11030
rect 40123 -11038 40167 -11030
rect 40223 -11038 40267 -11030
rect 40323 -11038 40367 -11030
rect 40423 -11038 40467 -11030
rect 40523 -11038 40567 -11030
rect 40623 -11038 40667 -11030
rect 40723 -11038 40767 -11030
rect 41223 -11038 41267 -11030
rect 41323 -11038 41367 -11030
rect 41423 -11038 41467 -11030
rect 41523 -11038 41567 -11030
rect 41623 -11038 41667 -11030
rect 41723 -11038 41767 -11030
rect 41823 -11038 41867 -11030
rect 41923 -11038 41967 -11030
rect 42023 -11038 42067 -11030
rect 42123 -11038 42167 -11030
rect 42223 -11038 42267 -11030
rect 42323 -11038 42367 -11030
rect 42423 -11038 42467 -11030
rect 42523 -11038 42567 -11030
rect 42623 -11038 42667 -11030
rect 42723 -11038 42767 -11030
rect 43223 -11038 43267 -11030
rect 43323 -11038 43367 -11030
rect 43423 -11038 43467 -11030
rect 43523 -11038 43567 -11030
rect 43623 -11038 43667 -11030
rect 43723 -11038 43767 -11030
rect 43823 -11038 43867 -11030
rect 43923 -11038 43967 -11030
rect 44023 -11038 44067 -11030
rect 44123 -11038 44167 -11030
rect 44223 -11038 44267 -11030
rect 44323 -11038 44367 -11030
rect 44423 -11038 44467 -11030
rect 44523 -11038 44567 -11030
rect 44623 -11038 44667 -11030
rect 44723 -11038 44767 -11030
rect 9195 -11056 9239 -11048
rect 9295 -11056 9339 -11048
rect 9395 -11056 9439 -11048
rect 9495 -11056 9539 -11048
rect 9595 -11056 9639 -11048
rect 9695 -11056 9739 -11048
rect 9795 -11056 9839 -11048
rect 9895 -11056 9939 -11048
rect 9995 -11056 10039 -11048
rect 10095 -11056 10139 -11048
rect 10195 -11056 10239 -11048
rect 10295 -11056 10339 -11048
rect 10395 -11056 10439 -11048
rect 10495 -11056 10539 -11048
rect 10595 -11056 10639 -11048
rect 10695 -11056 10739 -11048
rect 11195 -11056 11239 -11048
rect 11295 -11056 11339 -11048
rect 11395 -11056 11439 -11048
rect 11495 -11056 11539 -11048
rect 11595 -11056 11639 -11048
rect 11695 -11056 11739 -11048
rect 11795 -11056 11839 -11048
rect 11895 -11056 11939 -11048
rect 11995 -11056 12039 -11048
rect 12095 -11056 12139 -11048
rect 12195 -11056 12239 -11048
rect 12295 -11056 12339 -11048
rect 12395 -11056 12439 -11048
rect 12495 -11056 12539 -11048
rect 12595 -11056 12639 -11048
rect 12695 -11056 12739 -11048
rect 13195 -11056 13239 -11048
rect 13295 -11056 13339 -11048
rect 13395 -11056 13439 -11048
rect 13495 -11056 13539 -11048
rect 13595 -11056 13639 -11048
rect 13695 -11056 13739 -11048
rect 13795 -11056 13839 -11048
rect 13895 -11056 13939 -11048
rect 13995 -11056 14039 -11048
rect 14095 -11056 14139 -11048
rect 14195 -11056 14239 -11048
rect 14295 -11056 14339 -11048
rect 14395 -11056 14439 -11048
rect 14495 -11056 14539 -11048
rect 14595 -11056 14639 -11048
rect 14695 -11056 14739 -11048
rect 15195 -11056 15239 -11048
rect 15295 -11056 15339 -11048
rect 15395 -11056 15439 -11048
rect 15495 -11056 15539 -11048
rect 15595 -11056 15639 -11048
rect 15695 -11056 15739 -11048
rect 15795 -11056 15839 -11048
rect 15895 -11056 15939 -11048
rect 15995 -11056 16039 -11048
rect 16095 -11056 16139 -11048
rect 16195 -11056 16239 -11048
rect 16295 -11056 16339 -11048
rect 16395 -11056 16439 -11048
rect 16495 -11056 16539 -11048
rect 16595 -11056 16639 -11048
rect 16695 -11056 16739 -11048
rect 9239 -11100 9247 -11056
rect 9339 -11100 9347 -11056
rect 9439 -11100 9447 -11056
rect 9539 -11100 9547 -11056
rect 9639 -11100 9647 -11056
rect 9739 -11100 9747 -11056
rect 9839 -11100 9847 -11056
rect 9939 -11100 9947 -11056
rect 10039 -11100 10047 -11056
rect 10139 -11100 10147 -11056
rect 10239 -11100 10247 -11056
rect 10339 -11100 10347 -11056
rect 10439 -11100 10447 -11056
rect 10539 -11100 10547 -11056
rect 10639 -11100 10647 -11056
rect 10739 -11100 10747 -11056
rect 11239 -11100 11247 -11056
rect 11339 -11100 11347 -11056
rect 11439 -11100 11447 -11056
rect 11539 -11100 11547 -11056
rect 11639 -11100 11647 -11056
rect 11739 -11100 11747 -11056
rect 11839 -11100 11847 -11056
rect 11939 -11100 11947 -11056
rect 12039 -11100 12047 -11056
rect 12139 -11100 12147 -11056
rect 12239 -11100 12247 -11056
rect 12339 -11100 12347 -11056
rect 12439 -11100 12447 -11056
rect 12539 -11100 12547 -11056
rect 12639 -11100 12647 -11056
rect 12739 -11100 12747 -11056
rect 13239 -11100 13247 -11056
rect 13339 -11100 13347 -11056
rect 13439 -11100 13447 -11056
rect 13539 -11100 13547 -11056
rect 13639 -11100 13647 -11056
rect 13739 -11100 13747 -11056
rect 13839 -11100 13847 -11056
rect 13939 -11100 13947 -11056
rect 14039 -11100 14047 -11056
rect 14139 -11100 14147 -11056
rect 14239 -11100 14247 -11056
rect 14339 -11100 14347 -11056
rect 14439 -11100 14447 -11056
rect 14539 -11100 14547 -11056
rect 14639 -11100 14647 -11056
rect 14739 -11100 14747 -11056
rect 15239 -11100 15247 -11056
rect 15339 -11100 15347 -11056
rect 15439 -11100 15447 -11056
rect 15539 -11100 15547 -11056
rect 15639 -11100 15647 -11056
rect 15739 -11100 15747 -11056
rect 15839 -11100 15847 -11056
rect 15939 -11100 15947 -11056
rect 16039 -11100 16047 -11056
rect 16139 -11100 16147 -11056
rect 16239 -11100 16247 -11056
rect 16339 -11100 16347 -11056
rect 16439 -11100 16447 -11056
rect 16539 -11100 16547 -11056
rect 16639 -11100 16647 -11056
rect 16739 -11100 16747 -11056
rect 37267 -11082 37275 -11038
rect 37367 -11082 37375 -11038
rect 37467 -11082 37475 -11038
rect 37567 -11082 37575 -11038
rect 37667 -11082 37675 -11038
rect 37767 -11082 37775 -11038
rect 37867 -11082 37875 -11038
rect 37967 -11082 37975 -11038
rect 38067 -11082 38075 -11038
rect 38167 -11082 38175 -11038
rect 38267 -11082 38275 -11038
rect 38367 -11082 38375 -11038
rect 38467 -11082 38475 -11038
rect 38567 -11082 38575 -11038
rect 38667 -11082 38675 -11038
rect 38767 -11082 38775 -11038
rect 39267 -11082 39275 -11038
rect 39367 -11082 39375 -11038
rect 39467 -11082 39475 -11038
rect 39567 -11082 39575 -11038
rect 39667 -11082 39675 -11038
rect 39767 -11082 39775 -11038
rect 39867 -11082 39875 -11038
rect 39967 -11082 39975 -11038
rect 40067 -11082 40075 -11038
rect 40167 -11082 40175 -11038
rect 40267 -11082 40275 -11038
rect 40367 -11082 40375 -11038
rect 40467 -11082 40475 -11038
rect 40567 -11082 40575 -11038
rect 40667 -11082 40675 -11038
rect 40767 -11082 40775 -11038
rect 41267 -11082 41275 -11038
rect 41367 -11082 41375 -11038
rect 41467 -11082 41475 -11038
rect 41567 -11082 41575 -11038
rect 41667 -11082 41675 -11038
rect 41767 -11082 41775 -11038
rect 41867 -11082 41875 -11038
rect 41967 -11082 41975 -11038
rect 42067 -11082 42075 -11038
rect 42167 -11082 42175 -11038
rect 42267 -11082 42275 -11038
rect 42367 -11082 42375 -11038
rect 42467 -11082 42475 -11038
rect 42567 -11082 42575 -11038
rect 42667 -11082 42675 -11038
rect 42767 -11082 42775 -11038
rect 43267 -11082 43275 -11038
rect 43367 -11082 43375 -11038
rect 43467 -11082 43475 -11038
rect 43567 -11082 43575 -11038
rect 43667 -11082 43675 -11038
rect 43767 -11082 43775 -11038
rect 43867 -11082 43875 -11038
rect 43967 -11082 43975 -11038
rect 44067 -11082 44075 -11038
rect 44167 -11082 44175 -11038
rect 44267 -11082 44275 -11038
rect 44367 -11082 44375 -11038
rect 44467 -11082 44475 -11038
rect 44567 -11082 44575 -11038
rect 44667 -11082 44675 -11038
rect 44767 -11082 44775 -11038
rect 37223 -11138 37267 -11130
rect 37323 -11138 37367 -11130
rect 37423 -11138 37467 -11130
rect 37523 -11138 37567 -11130
rect 37623 -11138 37667 -11130
rect 37723 -11138 37767 -11130
rect 37823 -11138 37867 -11130
rect 37923 -11138 37967 -11130
rect 38023 -11138 38067 -11130
rect 38123 -11138 38167 -11130
rect 38223 -11138 38267 -11130
rect 38323 -11138 38367 -11130
rect 38423 -11138 38467 -11130
rect 38523 -11138 38567 -11130
rect 38623 -11138 38667 -11130
rect 38723 -11138 38767 -11130
rect 39223 -11138 39267 -11130
rect 39323 -11138 39367 -11130
rect 39423 -11138 39467 -11130
rect 39523 -11138 39567 -11130
rect 39623 -11138 39667 -11130
rect 39723 -11138 39767 -11130
rect 39823 -11138 39867 -11130
rect 39923 -11138 39967 -11130
rect 40023 -11138 40067 -11130
rect 40123 -11138 40167 -11130
rect 40223 -11138 40267 -11130
rect 40323 -11138 40367 -11130
rect 40423 -11138 40467 -11130
rect 40523 -11138 40567 -11130
rect 40623 -11138 40667 -11130
rect 40723 -11138 40767 -11130
rect 41223 -11138 41267 -11130
rect 41323 -11138 41367 -11130
rect 41423 -11138 41467 -11130
rect 41523 -11138 41567 -11130
rect 41623 -11138 41667 -11130
rect 41723 -11138 41767 -11130
rect 41823 -11138 41867 -11130
rect 41923 -11138 41967 -11130
rect 42023 -11138 42067 -11130
rect 42123 -11138 42167 -11130
rect 42223 -11138 42267 -11130
rect 42323 -11138 42367 -11130
rect 42423 -11138 42467 -11130
rect 42523 -11138 42567 -11130
rect 42623 -11138 42667 -11130
rect 42723 -11138 42767 -11130
rect 43223 -11138 43267 -11130
rect 43323 -11138 43367 -11130
rect 43423 -11138 43467 -11130
rect 43523 -11138 43567 -11130
rect 43623 -11138 43667 -11130
rect 43723 -11138 43767 -11130
rect 43823 -11138 43867 -11130
rect 43923 -11138 43967 -11130
rect 44023 -11138 44067 -11130
rect 44123 -11138 44167 -11130
rect 44223 -11138 44267 -11130
rect 44323 -11138 44367 -11130
rect 44423 -11138 44467 -11130
rect 44523 -11138 44567 -11130
rect 44623 -11138 44667 -11130
rect 44723 -11138 44767 -11130
rect 9195 -11156 9239 -11148
rect 9295 -11156 9339 -11148
rect 9395 -11156 9439 -11148
rect 9495 -11156 9539 -11148
rect 9595 -11156 9639 -11148
rect 9695 -11156 9739 -11148
rect 9795 -11156 9839 -11148
rect 9895 -11156 9939 -11148
rect 9995 -11156 10039 -11148
rect 10095 -11156 10139 -11148
rect 10195 -11156 10239 -11148
rect 10295 -11156 10339 -11148
rect 10395 -11156 10439 -11148
rect 10495 -11156 10539 -11148
rect 10595 -11156 10639 -11148
rect 10695 -11156 10739 -11148
rect 11195 -11156 11239 -11148
rect 11295 -11156 11339 -11148
rect 11395 -11156 11439 -11148
rect 11495 -11156 11539 -11148
rect 11595 -11156 11639 -11148
rect 11695 -11156 11739 -11148
rect 11795 -11156 11839 -11148
rect 11895 -11156 11939 -11148
rect 11995 -11156 12039 -11148
rect 12095 -11156 12139 -11148
rect 12195 -11156 12239 -11148
rect 12295 -11156 12339 -11148
rect 12395 -11156 12439 -11148
rect 12495 -11156 12539 -11148
rect 12595 -11156 12639 -11148
rect 12695 -11156 12739 -11148
rect 13195 -11156 13239 -11148
rect 13295 -11156 13339 -11148
rect 13395 -11156 13439 -11148
rect 13495 -11156 13539 -11148
rect 13595 -11156 13639 -11148
rect 13695 -11156 13739 -11148
rect 13795 -11156 13839 -11148
rect 13895 -11156 13939 -11148
rect 13995 -11156 14039 -11148
rect 14095 -11156 14139 -11148
rect 14195 -11156 14239 -11148
rect 14295 -11156 14339 -11148
rect 14395 -11156 14439 -11148
rect 14495 -11156 14539 -11148
rect 14595 -11156 14639 -11148
rect 14695 -11156 14739 -11148
rect 15195 -11156 15239 -11148
rect 15295 -11156 15339 -11148
rect 15395 -11156 15439 -11148
rect 15495 -11156 15539 -11148
rect 15595 -11156 15639 -11148
rect 15695 -11156 15739 -11148
rect 15795 -11156 15839 -11148
rect 15895 -11156 15939 -11148
rect 15995 -11156 16039 -11148
rect 16095 -11156 16139 -11148
rect 16195 -11156 16239 -11148
rect 16295 -11156 16339 -11148
rect 16395 -11156 16439 -11148
rect 16495 -11156 16539 -11148
rect 16595 -11156 16639 -11148
rect 16695 -11156 16739 -11148
rect 9239 -11200 9247 -11156
rect 9339 -11200 9347 -11156
rect 9439 -11200 9447 -11156
rect 9539 -11200 9547 -11156
rect 9639 -11200 9647 -11156
rect 9739 -11200 9747 -11156
rect 9839 -11200 9847 -11156
rect 9939 -11200 9947 -11156
rect 10039 -11200 10047 -11156
rect 10139 -11200 10147 -11156
rect 10239 -11200 10247 -11156
rect 10339 -11200 10347 -11156
rect 10439 -11200 10447 -11156
rect 10539 -11200 10547 -11156
rect 10639 -11200 10647 -11156
rect 10739 -11200 10747 -11156
rect 11239 -11200 11247 -11156
rect 11339 -11200 11347 -11156
rect 11439 -11200 11447 -11156
rect 11539 -11200 11547 -11156
rect 11639 -11200 11647 -11156
rect 11739 -11200 11747 -11156
rect 11839 -11200 11847 -11156
rect 11939 -11200 11947 -11156
rect 12039 -11200 12047 -11156
rect 12139 -11200 12147 -11156
rect 12239 -11200 12247 -11156
rect 12339 -11200 12347 -11156
rect 12439 -11200 12447 -11156
rect 12539 -11200 12547 -11156
rect 12639 -11200 12647 -11156
rect 12739 -11200 12747 -11156
rect 13239 -11200 13247 -11156
rect 13339 -11200 13347 -11156
rect 13439 -11200 13447 -11156
rect 13539 -11200 13547 -11156
rect 13639 -11200 13647 -11156
rect 13739 -11200 13747 -11156
rect 13839 -11200 13847 -11156
rect 13939 -11200 13947 -11156
rect 14039 -11200 14047 -11156
rect 14139 -11200 14147 -11156
rect 14239 -11200 14247 -11156
rect 14339 -11200 14347 -11156
rect 14439 -11200 14447 -11156
rect 14539 -11200 14547 -11156
rect 14639 -11200 14647 -11156
rect 14739 -11200 14747 -11156
rect 15239 -11200 15247 -11156
rect 15339 -11200 15347 -11156
rect 15439 -11200 15447 -11156
rect 15539 -11200 15547 -11156
rect 15639 -11200 15647 -11156
rect 15739 -11200 15747 -11156
rect 15839 -11200 15847 -11156
rect 15939 -11200 15947 -11156
rect 16039 -11200 16047 -11156
rect 16139 -11200 16147 -11156
rect 16239 -11200 16247 -11156
rect 16339 -11200 16347 -11156
rect 16439 -11200 16447 -11156
rect 16539 -11200 16547 -11156
rect 16639 -11200 16647 -11156
rect 16739 -11200 16747 -11156
rect 37267 -11182 37275 -11138
rect 37367 -11182 37375 -11138
rect 37467 -11182 37475 -11138
rect 37567 -11182 37575 -11138
rect 37667 -11182 37675 -11138
rect 37767 -11182 37775 -11138
rect 37867 -11182 37875 -11138
rect 37967 -11182 37975 -11138
rect 38067 -11182 38075 -11138
rect 38167 -11182 38175 -11138
rect 38267 -11182 38275 -11138
rect 38367 -11182 38375 -11138
rect 38467 -11182 38475 -11138
rect 38567 -11182 38575 -11138
rect 38667 -11182 38675 -11138
rect 38767 -11182 38775 -11138
rect 39267 -11182 39275 -11138
rect 39367 -11182 39375 -11138
rect 39467 -11182 39475 -11138
rect 39567 -11182 39575 -11138
rect 39667 -11182 39675 -11138
rect 39767 -11182 39775 -11138
rect 39867 -11182 39875 -11138
rect 39967 -11182 39975 -11138
rect 40067 -11182 40075 -11138
rect 40167 -11182 40175 -11138
rect 40267 -11182 40275 -11138
rect 40367 -11182 40375 -11138
rect 40467 -11182 40475 -11138
rect 40567 -11182 40575 -11138
rect 40667 -11182 40675 -11138
rect 40767 -11182 40775 -11138
rect 41267 -11182 41275 -11138
rect 41367 -11182 41375 -11138
rect 41467 -11182 41475 -11138
rect 41567 -11182 41575 -11138
rect 41667 -11182 41675 -11138
rect 41767 -11182 41775 -11138
rect 41867 -11182 41875 -11138
rect 41967 -11182 41975 -11138
rect 42067 -11182 42075 -11138
rect 42167 -11182 42175 -11138
rect 42267 -11182 42275 -11138
rect 42367 -11182 42375 -11138
rect 42467 -11182 42475 -11138
rect 42567 -11182 42575 -11138
rect 42667 -11182 42675 -11138
rect 42767 -11182 42775 -11138
rect 43267 -11182 43275 -11138
rect 43367 -11182 43375 -11138
rect 43467 -11182 43475 -11138
rect 43567 -11182 43575 -11138
rect 43667 -11182 43675 -11138
rect 43767 -11182 43775 -11138
rect 43867 -11182 43875 -11138
rect 43967 -11182 43975 -11138
rect 44067 -11182 44075 -11138
rect 44167 -11182 44175 -11138
rect 44267 -11182 44275 -11138
rect 44367 -11182 44375 -11138
rect 44467 -11182 44475 -11138
rect 44567 -11182 44575 -11138
rect 44667 -11182 44675 -11138
rect 44767 -11182 44775 -11138
rect 9195 -11256 9239 -11248
rect 9295 -11256 9339 -11248
rect 9395 -11256 9439 -11248
rect 9495 -11256 9539 -11248
rect 9595 -11256 9639 -11248
rect 9695 -11256 9739 -11248
rect 9795 -11256 9839 -11248
rect 9895 -11256 9939 -11248
rect 9995 -11256 10039 -11248
rect 10095 -11256 10139 -11248
rect 10195 -11256 10239 -11248
rect 10295 -11256 10339 -11248
rect 10395 -11256 10439 -11248
rect 10495 -11256 10539 -11248
rect 10595 -11256 10639 -11248
rect 10695 -11256 10739 -11248
rect 11195 -11256 11239 -11248
rect 11295 -11256 11339 -11248
rect 11395 -11256 11439 -11248
rect 11495 -11256 11539 -11248
rect 11595 -11256 11639 -11248
rect 11695 -11256 11739 -11248
rect 11795 -11256 11839 -11248
rect 11895 -11256 11939 -11248
rect 11995 -11256 12039 -11248
rect 12095 -11256 12139 -11248
rect 12195 -11256 12239 -11248
rect 12295 -11256 12339 -11248
rect 12395 -11256 12439 -11248
rect 12495 -11256 12539 -11248
rect 12595 -11256 12639 -11248
rect 12695 -11256 12739 -11248
rect 13195 -11256 13239 -11248
rect 13295 -11256 13339 -11248
rect 13395 -11256 13439 -11248
rect 13495 -11256 13539 -11248
rect 13595 -11256 13639 -11248
rect 13695 -11256 13739 -11248
rect 13795 -11256 13839 -11248
rect 13895 -11256 13939 -11248
rect 13995 -11256 14039 -11248
rect 14095 -11256 14139 -11248
rect 14195 -11256 14239 -11248
rect 14295 -11256 14339 -11248
rect 14395 -11256 14439 -11248
rect 14495 -11256 14539 -11248
rect 14595 -11256 14639 -11248
rect 14695 -11256 14739 -11248
rect 15195 -11256 15239 -11248
rect 15295 -11256 15339 -11248
rect 15395 -11256 15439 -11248
rect 15495 -11256 15539 -11248
rect 15595 -11256 15639 -11248
rect 15695 -11256 15739 -11248
rect 15795 -11256 15839 -11248
rect 15895 -11256 15939 -11248
rect 15995 -11256 16039 -11248
rect 16095 -11256 16139 -11248
rect 16195 -11256 16239 -11248
rect 16295 -11256 16339 -11248
rect 16395 -11256 16439 -11248
rect 16495 -11256 16539 -11248
rect 16595 -11256 16639 -11248
rect 16695 -11256 16739 -11248
rect 9239 -11300 9247 -11256
rect 9339 -11300 9347 -11256
rect 9439 -11300 9447 -11256
rect 9539 -11300 9547 -11256
rect 9639 -11300 9647 -11256
rect 9739 -11300 9747 -11256
rect 9839 -11300 9847 -11256
rect 9939 -11300 9947 -11256
rect 10039 -11300 10047 -11256
rect 10139 -11300 10147 -11256
rect 10239 -11300 10247 -11256
rect 10339 -11300 10347 -11256
rect 10439 -11300 10447 -11256
rect 10539 -11300 10547 -11256
rect 10639 -11300 10647 -11256
rect 10739 -11300 10747 -11256
rect 11239 -11300 11247 -11256
rect 11339 -11300 11347 -11256
rect 11439 -11300 11447 -11256
rect 11539 -11300 11547 -11256
rect 11639 -11300 11647 -11256
rect 11739 -11300 11747 -11256
rect 11839 -11300 11847 -11256
rect 11939 -11300 11947 -11256
rect 12039 -11300 12047 -11256
rect 12139 -11300 12147 -11256
rect 12239 -11300 12247 -11256
rect 12339 -11300 12347 -11256
rect 12439 -11300 12447 -11256
rect 12539 -11300 12547 -11256
rect 12639 -11300 12647 -11256
rect 12739 -11300 12747 -11256
rect 13239 -11300 13247 -11256
rect 13339 -11300 13347 -11256
rect 13439 -11300 13447 -11256
rect 13539 -11300 13547 -11256
rect 13639 -11300 13647 -11256
rect 13739 -11300 13747 -11256
rect 13839 -11300 13847 -11256
rect 13939 -11300 13947 -11256
rect 14039 -11300 14047 -11256
rect 14139 -11300 14147 -11256
rect 14239 -11300 14247 -11256
rect 14339 -11300 14347 -11256
rect 14439 -11300 14447 -11256
rect 14539 -11300 14547 -11256
rect 14639 -11300 14647 -11256
rect 14739 -11300 14747 -11256
rect 15239 -11300 15247 -11256
rect 15339 -11300 15347 -11256
rect 15439 -11300 15447 -11256
rect 15539 -11300 15547 -11256
rect 15639 -11300 15647 -11256
rect 15739 -11300 15747 -11256
rect 15839 -11300 15847 -11256
rect 15939 -11300 15947 -11256
rect 16039 -11300 16047 -11256
rect 16139 -11300 16147 -11256
rect 16239 -11300 16247 -11256
rect 16339 -11300 16347 -11256
rect 16439 -11300 16447 -11256
rect 16539 -11300 16547 -11256
rect 16639 -11300 16647 -11256
rect 16739 -11300 16747 -11256
rect 57950 -19693 57952 307
rect 58016 -19693 58018 307
rect 84950 -19693 84952 307
rect 85016 -19693 85018 307
rect 80849 -24026 80893 -24018
rect 80949 -24026 80993 -24018
rect 81049 -24026 81093 -24018
rect 81149 -24026 81193 -24018
rect 81249 -24026 81293 -24018
rect 81349 -24026 81393 -24018
rect 81449 -24026 81493 -24018
rect 81549 -24026 81593 -24018
rect 81649 -24026 81693 -24018
rect 81749 -24026 81793 -24018
rect 81849 -24026 81893 -24018
rect 81949 -24026 81993 -24018
rect 82049 -24026 82093 -24018
rect 82149 -24026 82193 -24018
rect 82249 -24026 82293 -24018
rect 82349 -24026 82393 -24018
rect 82849 -24026 82893 -24018
rect 82949 -24026 82993 -24018
rect 83049 -24026 83093 -24018
rect 83149 -24026 83193 -24018
rect 83249 -24026 83293 -24018
rect 83349 -24026 83393 -24018
rect 83449 -24026 83493 -24018
rect 83549 -24026 83593 -24018
rect 83649 -24026 83693 -24018
rect 83749 -24026 83793 -24018
rect 83849 -24026 83893 -24018
rect 83949 -24026 83993 -24018
rect 84049 -24026 84093 -24018
rect 84149 -24026 84193 -24018
rect 84249 -24026 84293 -24018
rect 84349 -24026 84393 -24018
rect 84849 -24026 84893 -24018
rect 84949 -24026 84993 -24018
rect 85049 -24026 85093 -24018
rect 85149 -24026 85193 -24018
rect 85249 -24026 85293 -24018
rect 85349 -24026 85393 -24018
rect 85449 -24026 85493 -24018
rect 85549 -24026 85593 -24018
rect 85649 -24026 85693 -24018
rect 85749 -24026 85793 -24018
rect 85849 -24026 85893 -24018
rect 85949 -24026 85993 -24018
rect 86049 -24026 86093 -24018
rect 86149 -24026 86193 -24018
rect 86249 -24026 86293 -24018
rect 86349 -24026 86393 -24018
rect 86849 -24026 86893 -24018
rect 86949 -24026 86993 -24018
rect 87049 -24026 87093 -24018
rect 87149 -24026 87193 -24018
rect 87249 -24026 87293 -24018
rect 87349 -24026 87393 -24018
rect 87449 -24026 87493 -24018
rect 87549 -24026 87593 -24018
rect 87649 -24026 87693 -24018
rect 87749 -24026 87793 -24018
rect 87849 -24026 87893 -24018
rect 87949 -24026 87993 -24018
rect 88049 -24026 88093 -24018
rect 88149 -24026 88193 -24018
rect 88249 -24026 88293 -24018
rect 88349 -24026 88393 -24018
rect 80893 -24070 80901 -24026
rect 80993 -24070 81001 -24026
rect 81093 -24070 81101 -24026
rect 81193 -24070 81201 -24026
rect 81293 -24070 81301 -24026
rect 81393 -24070 81401 -24026
rect 81493 -24070 81501 -24026
rect 81593 -24070 81601 -24026
rect 81693 -24070 81701 -24026
rect 81793 -24070 81801 -24026
rect 81893 -24070 81901 -24026
rect 81993 -24070 82001 -24026
rect 82093 -24070 82101 -24026
rect 82193 -24070 82201 -24026
rect 82293 -24070 82301 -24026
rect 82393 -24070 82401 -24026
rect 82893 -24070 82901 -24026
rect 82993 -24070 83001 -24026
rect 83093 -24070 83101 -24026
rect 83193 -24070 83201 -24026
rect 83293 -24070 83301 -24026
rect 83393 -24070 83401 -24026
rect 83493 -24070 83501 -24026
rect 83593 -24070 83601 -24026
rect 83693 -24070 83701 -24026
rect 83793 -24070 83801 -24026
rect 83893 -24070 83901 -24026
rect 83993 -24070 84001 -24026
rect 84093 -24070 84101 -24026
rect 84193 -24070 84201 -24026
rect 84293 -24070 84301 -24026
rect 84393 -24070 84401 -24026
rect 84893 -24070 84901 -24026
rect 84993 -24070 85001 -24026
rect 85093 -24070 85101 -24026
rect 85193 -24070 85201 -24026
rect 85293 -24070 85301 -24026
rect 85393 -24070 85401 -24026
rect 85493 -24070 85501 -24026
rect 85593 -24070 85601 -24026
rect 85693 -24070 85701 -24026
rect 85793 -24070 85801 -24026
rect 85893 -24070 85901 -24026
rect 85993 -24070 86001 -24026
rect 86093 -24070 86101 -24026
rect 86193 -24070 86201 -24026
rect 86293 -24070 86301 -24026
rect 86393 -24070 86401 -24026
rect 86893 -24070 86901 -24026
rect 86993 -24070 87001 -24026
rect 87093 -24070 87101 -24026
rect 87193 -24070 87201 -24026
rect 87293 -24070 87301 -24026
rect 87393 -24070 87401 -24026
rect 87493 -24070 87501 -24026
rect 87593 -24070 87601 -24026
rect 87693 -24070 87701 -24026
rect 87793 -24070 87801 -24026
rect 87893 -24070 87901 -24026
rect 87993 -24070 88001 -24026
rect 88093 -24070 88101 -24026
rect 88193 -24070 88201 -24026
rect 88293 -24070 88301 -24026
rect 88393 -24070 88401 -24026
rect 80849 -24126 80893 -24118
rect 80949 -24126 80993 -24118
rect 81049 -24126 81093 -24118
rect 81149 -24126 81193 -24118
rect 81249 -24126 81293 -24118
rect 81349 -24126 81393 -24118
rect 81449 -24126 81493 -24118
rect 81549 -24126 81593 -24118
rect 81649 -24126 81693 -24118
rect 81749 -24126 81793 -24118
rect 81849 -24126 81893 -24118
rect 81949 -24126 81993 -24118
rect 82049 -24126 82093 -24118
rect 82149 -24126 82193 -24118
rect 82249 -24126 82293 -24118
rect 82349 -24126 82393 -24118
rect 82849 -24126 82893 -24118
rect 82949 -24126 82993 -24118
rect 83049 -24126 83093 -24118
rect 83149 -24126 83193 -24118
rect 83249 -24126 83293 -24118
rect 83349 -24126 83393 -24118
rect 83449 -24126 83493 -24118
rect 83549 -24126 83593 -24118
rect 83649 -24126 83693 -24118
rect 83749 -24126 83793 -24118
rect 83849 -24126 83893 -24118
rect 83949 -24126 83993 -24118
rect 84049 -24126 84093 -24118
rect 84149 -24126 84193 -24118
rect 84249 -24126 84293 -24118
rect 84349 -24126 84393 -24118
rect 84849 -24126 84893 -24118
rect 84949 -24126 84993 -24118
rect 85049 -24126 85093 -24118
rect 85149 -24126 85193 -24118
rect 85249 -24126 85293 -24118
rect 85349 -24126 85393 -24118
rect 85449 -24126 85493 -24118
rect 85549 -24126 85593 -24118
rect 85649 -24126 85693 -24118
rect 85749 -24126 85793 -24118
rect 85849 -24126 85893 -24118
rect 85949 -24126 85993 -24118
rect 86049 -24126 86093 -24118
rect 86149 -24126 86193 -24118
rect 86249 -24126 86293 -24118
rect 86349 -24126 86393 -24118
rect 86849 -24126 86893 -24118
rect 86949 -24126 86993 -24118
rect 87049 -24126 87093 -24118
rect 87149 -24126 87193 -24118
rect 87249 -24126 87293 -24118
rect 87349 -24126 87393 -24118
rect 87449 -24126 87493 -24118
rect 87549 -24126 87593 -24118
rect 87649 -24126 87693 -24118
rect 87749 -24126 87793 -24118
rect 87849 -24126 87893 -24118
rect 87949 -24126 87993 -24118
rect 88049 -24126 88093 -24118
rect 88149 -24126 88193 -24118
rect 88249 -24126 88293 -24118
rect 88349 -24126 88393 -24118
rect 80893 -24170 80901 -24126
rect 80993 -24170 81001 -24126
rect 81093 -24170 81101 -24126
rect 81193 -24170 81201 -24126
rect 81293 -24170 81301 -24126
rect 81393 -24170 81401 -24126
rect 81493 -24170 81501 -24126
rect 81593 -24170 81601 -24126
rect 81693 -24170 81701 -24126
rect 81793 -24170 81801 -24126
rect 81893 -24170 81901 -24126
rect 81993 -24170 82001 -24126
rect 82093 -24170 82101 -24126
rect 82193 -24170 82201 -24126
rect 82293 -24170 82301 -24126
rect 82393 -24170 82401 -24126
rect 82893 -24170 82901 -24126
rect 82993 -24170 83001 -24126
rect 83093 -24170 83101 -24126
rect 83193 -24170 83201 -24126
rect 83293 -24170 83301 -24126
rect 83393 -24170 83401 -24126
rect 83493 -24170 83501 -24126
rect 83593 -24170 83601 -24126
rect 83693 -24170 83701 -24126
rect 83793 -24170 83801 -24126
rect 83893 -24170 83901 -24126
rect 83993 -24170 84001 -24126
rect 84093 -24170 84101 -24126
rect 84193 -24170 84201 -24126
rect 84293 -24170 84301 -24126
rect 84393 -24170 84401 -24126
rect 84893 -24170 84901 -24126
rect 84993 -24170 85001 -24126
rect 85093 -24170 85101 -24126
rect 85193 -24170 85201 -24126
rect 85293 -24170 85301 -24126
rect 85393 -24170 85401 -24126
rect 85493 -24170 85501 -24126
rect 85593 -24170 85601 -24126
rect 85693 -24170 85701 -24126
rect 85793 -24170 85801 -24126
rect 85893 -24170 85901 -24126
rect 85993 -24170 86001 -24126
rect 86093 -24170 86101 -24126
rect 86193 -24170 86201 -24126
rect 86293 -24170 86301 -24126
rect 86393 -24170 86401 -24126
rect 86893 -24170 86901 -24126
rect 86993 -24170 87001 -24126
rect 87093 -24170 87101 -24126
rect 87193 -24170 87201 -24126
rect 87293 -24170 87301 -24126
rect 87393 -24170 87401 -24126
rect 87493 -24170 87501 -24126
rect 87593 -24170 87601 -24126
rect 87693 -24170 87701 -24126
rect 87793 -24170 87801 -24126
rect 87893 -24170 87901 -24126
rect 87993 -24170 88001 -24126
rect 88093 -24170 88101 -24126
rect 88193 -24170 88201 -24126
rect 88293 -24170 88301 -24126
rect 88393 -24170 88401 -24126
rect 109104 -24195 109148 -24187
rect 109204 -24195 109248 -24187
rect 109304 -24195 109348 -24187
rect 109404 -24195 109448 -24187
rect 109504 -24195 109548 -24187
rect 109604 -24195 109648 -24187
rect 109704 -24195 109748 -24187
rect 109804 -24195 109848 -24187
rect 109904 -24195 109948 -24187
rect 110004 -24195 110048 -24187
rect 110104 -24195 110148 -24187
rect 110204 -24195 110248 -24187
rect 110304 -24195 110348 -24187
rect 110404 -24195 110448 -24187
rect 110504 -24195 110548 -24187
rect 110604 -24195 110648 -24187
rect 111104 -24195 111148 -24187
rect 111204 -24195 111248 -24187
rect 111304 -24195 111348 -24187
rect 111404 -24195 111448 -24187
rect 111504 -24195 111548 -24187
rect 111604 -24195 111648 -24187
rect 111704 -24195 111748 -24187
rect 111804 -24195 111848 -24187
rect 111904 -24195 111948 -24187
rect 112004 -24195 112048 -24187
rect 112104 -24195 112148 -24187
rect 112204 -24195 112248 -24187
rect 112304 -24195 112348 -24187
rect 112404 -24195 112448 -24187
rect 112504 -24195 112548 -24187
rect 112604 -24195 112648 -24187
rect 113104 -24195 113148 -24187
rect 113204 -24195 113248 -24187
rect 113304 -24195 113348 -24187
rect 113404 -24195 113448 -24187
rect 113504 -24195 113548 -24187
rect 113604 -24195 113648 -24187
rect 113704 -24195 113748 -24187
rect 113804 -24195 113848 -24187
rect 113904 -24195 113948 -24187
rect 114004 -24195 114048 -24187
rect 114104 -24195 114148 -24187
rect 114204 -24195 114248 -24187
rect 114304 -24195 114348 -24187
rect 114404 -24195 114448 -24187
rect 114504 -24195 114548 -24187
rect 114604 -24195 114648 -24187
rect 115104 -24195 115148 -24187
rect 115204 -24195 115248 -24187
rect 115304 -24195 115348 -24187
rect 115404 -24195 115448 -24187
rect 115504 -24195 115548 -24187
rect 115604 -24195 115648 -24187
rect 115704 -24195 115748 -24187
rect 115804 -24195 115848 -24187
rect 115904 -24195 115948 -24187
rect 116004 -24195 116048 -24187
rect 116104 -24195 116148 -24187
rect 116204 -24195 116248 -24187
rect 116304 -24195 116348 -24187
rect 116404 -24195 116448 -24187
rect 116504 -24195 116548 -24187
rect 116604 -24195 116648 -24187
rect 80849 -24226 80893 -24218
rect 80949 -24226 80993 -24218
rect 81049 -24226 81093 -24218
rect 81149 -24226 81193 -24218
rect 81249 -24226 81293 -24218
rect 81349 -24226 81393 -24218
rect 81449 -24226 81493 -24218
rect 81549 -24226 81593 -24218
rect 81649 -24226 81693 -24218
rect 81749 -24226 81793 -24218
rect 81849 -24226 81893 -24218
rect 81949 -24226 81993 -24218
rect 82049 -24226 82093 -24218
rect 82149 -24226 82193 -24218
rect 82249 -24226 82293 -24218
rect 82349 -24226 82393 -24218
rect 82849 -24226 82893 -24218
rect 82949 -24226 82993 -24218
rect 83049 -24226 83093 -24218
rect 83149 -24226 83193 -24218
rect 83249 -24226 83293 -24218
rect 83349 -24226 83393 -24218
rect 83449 -24226 83493 -24218
rect 83549 -24226 83593 -24218
rect 83649 -24226 83693 -24218
rect 83749 -24226 83793 -24218
rect 83849 -24226 83893 -24218
rect 83949 -24226 83993 -24218
rect 84049 -24226 84093 -24218
rect 84149 -24226 84193 -24218
rect 84249 -24226 84293 -24218
rect 84349 -24226 84393 -24218
rect 84849 -24226 84893 -24218
rect 84949 -24226 84993 -24218
rect 85049 -24226 85093 -24218
rect 85149 -24226 85193 -24218
rect 85249 -24226 85293 -24218
rect 85349 -24226 85393 -24218
rect 85449 -24226 85493 -24218
rect 85549 -24226 85593 -24218
rect 85649 -24226 85693 -24218
rect 85749 -24226 85793 -24218
rect 85849 -24226 85893 -24218
rect 85949 -24226 85993 -24218
rect 86049 -24226 86093 -24218
rect 86149 -24226 86193 -24218
rect 86249 -24226 86293 -24218
rect 86349 -24226 86393 -24218
rect 86849 -24226 86893 -24218
rect 86949 -24226 86993 -24218
rect 87049 -24226 87093 -24218
rect 87149 -24226 87193 -24218
rect 87249 -24226 87293 -24218
rect 87349 -24226 87393 -24218
rect 87449 -24226 87493 -24218
rect 87549 -24226 87593 -24218
rect 87649 -24226 87693 -24218
rect 87749 -24226 87793 -24218
rect 87849 -24226 87893 -24218
rect 87949 -24226 87993 -24218
rect 88049 -24226 88093 -24218
rect 88149 -24226 88193 -24218
rect 88249 -24226 88293 -24218
rect 88349 -24226 88393 -24218
rect 80893 -24270 80901 -24226
rect 80993 -24270 81001 -24226
rect 81093 -24270 81101 -24226
rect 81193 -24270 81201 -24226
rect 81293 -24270 81301 -24226
rect 81393 -24270 81401 -24226
rect 81493 -24270 81501 -24226
rect 81593 -24270 81601 -24226
rect 81693 -24270 81701 -24226
rect 81793 -24270 81801 -24226
rect 81893 -24270 81901 -24226
rect 81993 -24270 82001 -24226
rect 82093 -24270 82101 -24226
rect 82193 -24270 82201 -24226
rect 82293 -24270 82301 -24226
rect 82393 -24270 82401 -24226
rect 82893 -24270 82901 -24226
rect 82993 -24270 83001 -24226
rect 83093 -24270 83101 -24226
rect 83193 -24270 83201 -24226
rect 83293 -24270 83301 -24226
rect 83393 -24270 83401 -24226
rect 83493 -24270 83501 -24226
rect 83593 -24270 83601 -24226
rect 83693 -24270 83701 -24226
rect 83793 -24270 83801 -24226
rect 83893 -24270 83901 -24226
rect 83993 -24270 84001 -24226
rect 84093 -24270 84101 -24226
rect 84193 -24270 84201 -24226
rect 84293 -24270 84301 -24226
rect 84393 -24270 84401 -24226
rect 84893 -24270 84901 -24226
rect 84993 -24270 85001 -24226
rect 85093 -24270 85101 -24226
rect 85193 -24270 85201 -24226
rect 85293 -24270 85301 -24226
rect 85393 -24270 85401 -24226
rect 85493 -24270 85501 -24226
rect 85593 -24270 85601 -24226
rect 85693 -24270 85701 -24226
rect 85793 -24270 85801 -24226
rect 85893 -24270 85901 -24226
rect 85993 -24270 86001 -24226
rect 86093 -24270 86101 -24226
rect 86193 -24270 86201 -24226
rect 86293 -24270 86301 -24226
rect 86393 -24270 86401 -24226
rect 86893 -24270 86901 -24226
rect 86993 -24270 87001 -24226
rect 87093 -24270 87101 -24226
rect 87193 -24270 87201 -24226
rect 87293 -24270 87301 -24226
rect 87393 -24270 87401 -24226
rect 87493 -24270 87501 -24226
rect 87593 -24270 87601 -24226
rect 87693 -24270 87701 -24226
rect 87793 -24270 87801 -24226
rect 87893 -24270 87901 -24226
rect 87993 -24270 88001 -24226
rect 88093 -24270 88101 -24226
rect 88193 -24270 88201 -24226
rect 88293 -24270 88301 -24226
rect 88393 -24270 88401 -24226
rect 109148 -24239 109156 -24195
rect 109248 -24239 109256 -24195
rect 109348 -24239 109356 -24195
rect 109448 -24239 109456 -24195
rect 109548 -24239 109556 -24195
rect 109648 -24239 109656 -24195
rect 109748 -24239 109756 -24195
rect 109848 -24239 109856 -24195
rect 109948 -24239 109956 -24195
rect 110048 -24239 110056 -24195
rect 110148 -24239 110156 -24195
rect 110248 -24239 110256 -24195
rect 110348 -24239 110356 -24195
rect 110448 -24239 110456 -24195
rect 110548 -24239 110556 -24195
rect 110648 -24239 110656 -24195
rect 111148 -24239 111156 -24195
rect 111248 -24239 111256 -24195
rect 111348 -24239 111356 -24195
rect 111448 -24239 111456 -24195
rect 111548 -24239 111556 -24195
rect 111648 -24239 111656 -24195
rect 111748 -24239 111756 -24195
rect 111848 -24239 111856 -24195
rect 111948 -24239 111956 -24195
rect 112048 -24239 112056 -24195
rect 112148 -24239 112156 -24195
rect 112248 -24239 112256 -24195
rect 112348 -24239 112356 -24195
rect 112448 -24239 112456 -24195
rect 112548 -24239 112556 -24195
rect 112648 -24239 112656 -24195
rect 113148 -24239 113156 -24195
rect 113248 -24239 113256 -24195
rect 113348 -24239 113356 -24195
rect 113448 -24239 113456 -24195
rect 113548 -24239 113556 -24195
rect 113648 -24239 113656 -24195
rect 113748 -24239 113756 -24195
rect 113848 -24239 113856 -24195
rect 113948 -24239 113956 -24195
rect 114048 -24239 114056 -24195
rect 114148 -24239 114156 -24195
rect 114248 -24239 114256 -24195
rect 114348 -24239 114356 -24195
rect 114448 -24239 114456 -24195
rect 114548 -24239 114556 -24195
rect 114648 -24239 114656 -24195
rect 115148 -24239 115156 -24195
rect 115248 -24239 115256 -24195
rect 115348 -24239 115356 -24195
rect 115448 -24239 115456 -24195
rect 115548 -24239 115556 -24195
rect 115648 -24239 115656 -24195
rect 115748 -24239 115756 -24195
rect 115848 -24239 115856 -24195
rect 115948 -24239 115956 -24195
rect 116048 -24239 116056 -24195
rect 116148 -24239 116156 -24195
rect 116248 -24239 116256 -24195
rect 116348 -24239 116356 -24195
rect 116448 -24239 116456 -24195
rect 116548 -24239 116556 -24195
rect 116648 -24239 116656 -24195
rect 109104 -24295 109148 -24287
rect 109204 -24295 109248 -24287
rect 109304 -24295 109348 -24287
rect 109404 -24295 109448 -24287
rect 109504 -24295 109548 -24287
rect 109604 -24295 109648 -24287
rect 109704 -24295 109748 -24287
rect 109804 -24295 109848 -24287
rect 109904 -24295 109948 -24287
rect 110004 -24295 110048 -24287
rect 110104 -24295 110148 -24287
rect 110204 -24295 110248 -24287
rect 110304 -24295 110348 -24287
rect 110404 -24295 110448 -24287
rect 110504 -24295 110548 -24287
rect 110604 -24295 110648 -24287
rect 111104 -24295 111148 -24287
rect 111204 -24295 111248 -24287
rect 111304 -24295 111348 -24287
rect 111404 -24295 111448 -24287
rect 111504 -24295 111548 -24287
rect 111604 -24295 111648 -24287
rect 111704 -24295 111748 -24287
rect 111804 -24295 111848 -24287
rect 111904 -24295 111948 -24287
rect 112004 -24295 112048 -24287
rect 112104 -24295 112148 -24287
rect 112204 -24295 112248 -24287
rect 112304 -24295 112348 -24287
rect 112404 -24295 112448 -24287
rect 112504 -24295 112548 -24287
rect 112604 -24295 112648 -24287
rect 113104 -24295 113148 -24287
rect 113204 -24295 113248 -24287
rect 113304 -24295 113348 -24287
rect 113404 -24295 113448 -24287
rect 113504 -24295 113548 -24287
rect 113604 -24295 113648 -24287
rect 113704 -24295 113748 -24287
rect 113804 -24295 113848 -24287
rect 113904 -24295 113948 -24287
rect 114004 -24295 114048 -24287
rect 114104 -24295 114148 -24287
rect 114204 -24295 114248 -24287
rect 114304 -24295 114348 -24287
rect 114404 -24295 114448 -24287
rect 114504 -24295 114548 -24287
rect 114604 -24295 114648 -24287
rect 115104 -24295 115148 -24287
rect 115204 -24295 115248 -24287
rect 115304 -24295 115348 -24287
rect 115404 -24295 115448 -24287
rect 115504 -24295 115548 -24287
rect 115604 -24295 115648 -24287
rect 115704 -24295 115748 -24287
rect 115804 -24295 115848 -24287
rect 115904 -24295 115948 -24287
rect 116004 -24295 116048 -24287
rect 116104 -24295 116148 -24287
rect 116204 -24295 116248 -24287
rect 116304 -24295 116348 -24287
rect 116404 -24295 116448 -24287
rect 116504 -24295 116548 -24287
rect 116604 -24295 116648 -24287
rect 80849 -24326 80893 -24318
rect 80949 -24326 80993 -24318
rect 81049 -24326 81093 -24318
rect 81149 -24326 81193 -24318
rect 81249 -24326 81293 -24318
rect 81349 -24326 81393 -24318
rect 81449 -24326 81493 -24318
rect 81549 -24326 81593 -24318
rect 81649 -24326 81693 -24318
rect 81749 -24326 81793 -24318
rect 81849 -24326 81893 -24318
rect 81949 -24326 81993 -24318
rect 82049 -24326 82093 -24318
rect 82149 -24326 82193 -24318
rect 82249 -24326 82293 -24318
rect 82349 -24326 82393 -24318
rect 82849 -24326 82893 -24318
rect 82949 -24326 82993 -24318
rect 83049 -24326 83093 -24318
rect 83149 -24326 83193 -24318
rect 83249 -24326 83293 -24318
rect 83349 -24326 83393 -24318
rect 83449 -24326 83493 -24318
rect 83549 -24326 83593 -24318
rect 83649 -24326 83693 -24318
rect 83749 -24326 83793 -24318
rect 83849 -24326 83893 -24318
rect 83949 -24326 83993 -24318
rect 84049 -24326 84093 -24318
rect 84149 -24326 84193 -24318
rect 84249 -24326 84293 -24318
rect 84349 -24326 84393 -24318
rect 84849 -24326 84893 -24318
rect 84949 -24326 84993 -24318
rect 85049 -24326 85093 -24318
rect 85149 -24326 85193 -24318
rect 85249 -24326 85293 -24318
rect 85349 -24326 85393 -24318
rect 85449 -24326 85493 -24318
rect 85549 -24326 85593 -24318
rect 85649 -24326 85693 -24318
rect 85749 -24326 85793 -24318
rect 85849 -24326 85893 -24318
rect 85949 -24326 85993 -24318
rect 86049 -24326 86093 -24318
rect 86149 -24326 86193 -24318
rect 86249 -24326 86293 -24318
rect 86349 -24326 86393 -24318
rect 86849 -24326 86893 -24318
rect 86949 -24326 86993 -24318
rect 87049 -24326 87093 -24318
rect 87149 -24326 87193 -24318
rect 87249 -24326 87293 -24318
rect 87349 -24326 87393 -24318
rect 87449 -24326 87493 -24318
rect 87549 -24326 87593 -24318
rect 87649 -24326 87693 -24318
rect 87749 -24326 87793 -24318
rect 87849 -24326 87893 -24318
rect 87949 -24326 87993 -24318
rect 88049 -24326 88093 -24318
rect 88149 -24326 88193 -24318
rect 88249 -24326 88293 -24318
rect 88349 -24326 88393 -24318
rect 80893 -24370 80901 -24326
rect 80993 -24370 81001 -24326
rect 81093 -24370 81101 -24326
rect 81193 -24370 81201 -24326
rect 81293 -24370 81301 -24326
rect 81393 -24370 81401 -24326
rect 81493 -24370 81501 -24326
rect 81593 -24370 81601 -24326
rect 81693 -24370 81701 -24326
rect 81793 -24370 81801 -24326
rect 81893 -24370 81901 -24326
rect 81993 -24370 82001 -24326
rect 82093 -24370 82101 -24326
rect 82193 -24370 82201 -24326
rect 82293 -24370 82301 -24326
rect 82393 -24370 82401 -24326
rect 82893 -24370 82901 -24326
rect 82993 -24370 83001 -24326
rect 83093 -24370 83101 -24326
rect 83193 -24370 83201 -24326
rect 83293 -24370 83301 -24326
rect 83393 -24370 83401 -24326
rect 83493 -24370 83501 -24326
rect 83593 -24370 83601 -24326
rect 83693 -24370 83701 -24326
rect 83793 -24370 83801 -24326
rect 83893 -24370 83901 -24326
rect 83993 -24370 84001 -24326
rect 84093 -24370 84101 -24326
rect 84193 -24370 84201 -24326
rect 84293 -24370 84301 -24326
rect 84393 -24370 84401 -24326
rect 84893 -24370 84901 -24326
rect 84993 -24370 85001 -24326
rect 85093 -24370 85101 -24326
rect 85193 -24370 85201 -24326
rect 85293 -24370 85301 -24326
rect 85393 -24370 85401 -24326
rect 85493 -24370 85501 -24326
rect 85593 -24370 85601 -24326
rect 85693 -24370 85701 -24326
rect 85793 -24370 85801 -24326
rect 85893 -24370 85901 -24326
rect 85993 -24370 86001 -24326
rect 86093 -24370 86101 -24326
rect 86193 -24370 86201 -24326
rect 86293 -24370 86301 -24326
rect 86393 -24370 86401 -24326
rect 86893 -24370 86901 -24326
rect 86993 -24370 87001 -24326
rect 87093 -24370 87101 -24326
rect 87193 -24370 87201 -24326
rect 87293 -24370 87301 -24326
rect 87393 -24370 87401 -24326
rect 87493 -24370 87501 -24326
rect 87593 -24370 87601 -24326
rect 87693 -24370 87701 -24326
rect 87793 -24370 87801 -24326
rect 87893 -24370 87901 -24326
rect 87993 -24370 88001 -24326
rect 88093 -24370 88101 -24326
rect 88193 -24370 88201 -24326
rect 88293 -24370 88301 -24326
rect 88393 -24370 88401 -24326
rect 109148 -24339 109156 -24295
rect 109248 -24339 109256 -24295
rect 109348 -24339 109356 -24295
rect 109448 -24339 109456 -24295
rect 109548 -24339 109556 -24295
rect 109648 -24339 109656 -24295
rect 109748 -24339 109756 -24295
rect 109848 -24339 109856 -24295
rect 109948 -24339 109956 -24295
rect 110048 -24339 110056 -24295
rect 110148 -24339 110156 -24295
rect 110248 -24339 110256 -24295
rect 110348 -24339 110356 -24295
rect 110448 -24339 110456 -24295
rect 110548 -24339 110556 -24295
rect 110648 -24339 110656 -24295
rect 111148 -24339 111156 -24295
rect 111248 -24339 111256 -24295
rect 111348 -24339 111356 -24295
rect 111448 -24339 111456 -24295
rect 111548 -24339 111556 -24295
rect 111648 -24339 111656 -24295
rect 111748 -24339 111756 -24295
rect 111848 -24339 111856 -24295
rect 111948 -24339 111956 -24295
rect 112048 -24339 112056 -24295
rect 112148 -24339 112156 -24295
rect 112248 -24339 112256 -24295
rect 112348 -24339 112356 -24295
rect 112448 -24339 112456 -24295
rect 112548 -24339 112556 -24295
rect 112648 -24339 112656 -24295
rect 113148 -24339 113156 -24295
rect 113248 -24339 113256 -24295
rect 113348 -24339 113356 -24295
rect 113448 -24339 113456 -24295
rect 113548 -24339 113556 -24295
rect 113648 -24339 113656 -24295
rect 113748 -24339 113756 -24295
rect 113848 -24339 113856 -24295
rect 113948 -24339 113956 -24295
rect 114048 -24339 114056 -24295
rect 114148 -24339 114156 -24295
rect 114248 -24339 114256 -24295
rect 114348 -24339 114356 -24295
rect 114448 -24339 114456 -24295
rect 114548 -24339 114556 -24295
rect 114648 -24339 114656 -24295
rect 115148 -24339 115156 -24295
rect 115248 -24339 115256 -24295
rect 115348 -24339 115356 -24295
rect 115448 -24339 115456 -24295
rect 115548 -24339 115556 -24295
rect 115648 -24339 115656 -24295
rect 115748 -24339 115756 -24295
rect 115848 -24339 115856 -24295
rect 115948 -24339 115956 -24295
rect 116048 -24339 116056 -24295
rect 116148 -24339 116156 -24295
rect 116248 -24339 116256 -24295
rect 116348 -24339 116356 -24295
rect 116448 -24339 116456 -24295
rect 116548 -24339 116556 -24295
rect 116648 -24339 116656 -24295
rect 109104 -24395 109148 -24387
rect 109204 -24395 109248 -24387
rect 109304 -24395 109348 -24387
rect 109404 -24395 109448 -24387
rect 109504 -24395 109548 -24387
rect 109604 -24395 109648 -24387
rect 109704 -24395 109748 -24387
rect 109804 -24395 109848 -24387
rect 109904 -24395 109948 -24387
rect 110004 -24395 110048 -24387
rect 110104 -24395 110148 -24387
rect 110204 -24395 110248 -24387
rect 110304 -24395 110348 -24387
rect 110404 -24395 110448 -24387
rect 110504 -24395 110548 -24387
rect 110604 -24395 110648 -24387
rect 111104 -24395 111148 -24387
rect 111204 -24395 111248 -24387
rect 111304 -24395 111348 -24387
rect 111404 -24395 111448 -24387
rect 111504 -24395 111548 -24387
rect 111604 -24395 111648 -24387
rect 111704 -24395 111748 -24387
rect 111804 -24395 111848 -24387
rect 111904 -24395 111948 -24387
rect 112004 -24395 112048 -24387
rect 112104 -24395 112148 -24387
rect 112204 -24395 112248 -24387
rect 112304 -24395 112348 -24387
rect 112404 -24395 112448 -24387
rect 112504 -24395 112548 -24387
rect 112604 -24395 112648 -24387
rect 113104 -24395 113148 -24387
rect 113204 -24395 113248 -24387
rect 113304 -24395 113348 -24387
rect 113404 -24395 113448 -24387
rect 113504 -24395 113548 -24387
rect 113604 -24395 113648 -24387
rect 113704 -24395 113748 -24387
rect 113804 -24395 113848 -24387
rect 113904 -24395 113948 -24387
rect 114004 -24395 114048 -24387
rect 114104 -24395 114148 -24387
rect 114204 -24395 114248 -24387
rect 114304 -24395 114348 -24387
rect 114404 -24395 114448 -24387
rect 114504 -24395 114548 -24387
rect 114604 -24395 114648 -24387
rect 115104 -24395 115148 -24387
rect 115204 -24395 115248 -24387
rect 115304 -24395 115348 -24387
rect 115404 -24395 115448 -24387
rect 115504 -24395 115548 -24387
rect 115604 -24395 115648 -24387
rect 115704 -24395 115748 -24387
rect 115804 -24395 115848 -24387
rect 115904 -24395 115948 -24387
rect 116004 -24395 116048 -24387
rect 116104 -24395 116148 -24387
rect 116204 -24395 116248 -24387
rect 116304 -24395 116348 -24387
rect 116404 -24395 116448 -24387
rect 116504 -24395 116548 -24387
rect 116604 -24395 116648 -24387
rect 80849 -24426 80893 -24418
rect 80949 -24426 80993 -24418
rect 81049 -24426 81093 -24418
rect 81149 -24426 81193 -24418
rect 81249 -24426 81293 -24418
rect 81349 -24426 81393 -24418
rect 81449 -24426 81493 -24418
rect 81549 -24426 81593 -24418
rect 81649 -24426 81693 -24418
rect 81749 -24426 81793 -24418
rect 81849 -24426 81893 -24418
rect 81949 -24426 81993 -24418
rect 82049 -24426 82093 -24418
rect 82149 -24426 82193 -24418
rect 82249 -24426 82293 -24418
rect 82349 -24426 82393 -24418
rect 82849 -24426 82893 -24418
rect 82949 -24426 82993 -24418
rect 83049 -24426 83093 -24418
rect 83149 -24426 83193 -24418
rect 83249 -24426 83293 -24418
rect 83349 -24426 83393 -24418
rect 83449 -24426 83493 -24418
rect 83549 -24426 83593 -24418
rect 83649 -24426 83693 -24418
rect 83749 -24426 83793 -24418
rect 83849 -24426 83893 -24418
rect 83949 -24426 83993 -24418
rect 84049 -24426 84093 -24418
rect 84149 -24426 84193 -24418
rect 84249 -24426 84293 -24418
rect 84349 -24426 84393 -24418
rect 84849 -24426 84893 -24418
rect 84949 -24426 84993 -24418
rect 85049 -24426 85093 -24418
rect 85149 -24426 85193 -24418
rect 85249 -24426 85293 -24418
rect 85349 -24426 85393 -24418
rect 85449 -24426 85493 -24418
rect 85549 -24426 85593 -24418
rect 85649 -24426 85693 -24418
rect 85749 -24426 85793 -24418
rect 85849 -24426 85893 -24418
rect 85949 -24426 85993 -24418
rect 86049 -24426 86093 -24418
rect 86149 -24426 86193 -24418
rect 86249 -24426 86293 -24418
rect 86349 -24426 86393 -24418
rect 86849 -24426 86893 -24418
rect 86949 -24426 86993 -24418
rect 87049 -24426 87093 -24418
rect 87149 -24426 87193 -24418
rect 87249 -24426 87293 -24418
rect 87349 -24426 87393 -24418
rect 87449 -24426 87493 -24418
rect 87549 -24426 87593 -24418
rect 87649 -24426 87693 -24418
rect 87749 -24426 87793 -24418
rect 87849 -24426 87893 -24418
rect 87949 -24426 87993 -24418
rect 88049 -24426 88093 -24418
rect 88149 -24426 88193 -24418
rect 88249 -24426 88293 -24418
rect 88349 -24426 88393 -24418
rect 80893 -24470 80901 -24426
rect 80993 -24470 81001 -24426
rect 81093 -24470 81101 -24426
rect 81193 -24470 81201 -24426
rect 81293 -24470 81301 -24426
rect 81393 -24470 81401 -24426
rect 81493 -24470 81501 -24426
rect 81593 -24470 81601 -24426
rect 81693 -24470 81701 -24426
rect 81793 -24470 81801 -24426
rect 81893 -24470 81901 -24426
rect 81993 -24470 82001 -24426
rect 82093 -24470 82101 -24426
rect 82193 -24470 82201 -24426
rect 82293 -24470 82301 -24426
rect 82393 -24470 82401 -24426
rect 82893 -24470 82901 -24426
rect 82993 -24470 83001 -24426
rect 83093 -24470 83101 -24426
rect 83193 -24470 83201 -24426
rect 83293 -24470 83301 -24426
rect 83393 -24470 83401 -24426
rect 83493 -24470 83501 -24426
rect 83593 -24470 83601 -24426
rect 83693 -24470 83701 -24426
rect 83793 -24470 83801 -24426
rect 83893 -24470 83901 -24426
rect 83993 -24470 84001 -24426
rect 84093 -24470 84101 -24426
rect 84193 -24470 84201 -24426
rect 84293 -24470 84301 -24426
rect 84393 -24470 84401 -24426
rect 84893 -24470 84901 -24426
rect 84993 -24470 85001 -24426
rect 85093 -24470 85101 -24426
rect 85193 -24470 85201 -24426
rect 85293 -24470 85301 -24426
rect 85393 -24470 85401 -24426
rect 85493 -24470 85501 -24426
rect 85593 -24470 85601 -24426
rect 85693 -24470 85701 -24426
rect 85793 -24470 85801 -24426
rect 85893 -24470 85901 -24426
rect 85993 -24470 86001 -24426
rect 86093 -24470 86101 -24426
rect 86193 -24470 86201 -24426
rect 86293 -24470 86301 -24426
rect 86393 -24470 86401 -24426
rect 86893 -24470 86901 -24426
rect 86993 -24470 87001 -24426
rect 87093 -24470 87101 -24426
rect 87193 -24470 87201 -24426
rect 87293 -24470 87301 -24426
rect 87393 -24470 87401 -24426
rect 87493 -24470 87501 -24426
rect 87593 -24470 87601 -24426
rect 87693 -24470 87701 -24426
rect 87793 -24470 87801 -24426
rect 87893 -24470 87901 -24426
rect 87993 -24470 88001 -24426
rect 88093 -24470 88101 -24426
rect 88193 -24470 88201 -24426
rect 88293 -24470 88301 -24426
rect 88393 -24470 88401 -24426
rect 109148 -24439 109156 -24395
rect 109248 -24439 109256 -24395
rect 109348 -24439 109356 -24395
rect 109448 -24439 109456 -24395
rect 109548 -24439 109556 -24395
rect 109648 -24439 109656 -24395
rect 109748 -24439 109756 -24395
rect 109848 -24439 109856 -24395
rect 109948 -24439 109956 -24395
rect 110048 -24439 110056 -24395
rect 110148 -24439 110156 -24395
rect 110248 -24439 110256 -24395
rect 110348 -24439 110356 -24395
rect 110448 -24439 110456 -24395
rect 110548 -24439 110556 -24395
rect 110648 -24439 110656 -24395
rect 111148 -24439 111156 -24395
rect 111248 -24439 111256 -24395
rect 111348 -24439 111356 -24395
rect 111448 -24439 111456 -24395
rect 111548 -24439 111556 -24395
rect 111648 -24439 111656 -24395
rect 111748 -24439 111756 -24395
rect 111848 -24439 111856 -24395
rect 111948 -24439 111956 -24395
rect 112048 -24439 112056 -24395
rect 112148 -24439 112156 -24395
rect 112248 -24439 112256 -24395
rect 112348 -24439 112356 -24395
rect 112448 -24439 112456 -24395
rect 112548 -24439 112556 -24395
rect 112648 -24439 112656 -24395
rect 113148 -24439 113156 -24395
rect 113248 -24439 113256 -24395
rect 113348 -24439 113356 -24395
rect 113448 -24439 113456 -24395
rect 113548 -24439 113556 -24395
rect 113648 -24439 113656 -24395
rect 113748 -24439 113756 -24395
rect 113848 -24439 113856 -24395
rect 113948 -24439 113956 -24395
rect 114048 -24439 114056 -24395
rect 114148 -24439 114156 -24395
rect 114248 -24439 114256 -24395
rect 114348 -24439 114356 -24395
rect 114448 -24439 114456 -24395
rect 114548 -24439 114556 -24395
rect 114648 -24439 114656 -24395
rect 115148 -24439 115156 -24395
rect 115248 -24439 115256 -24395
rect 115348 -24439 115356 -24395
rect 115448 -24439 115456 -24395
rect 115548 -24439 115556 -24395
rect 115648 -24439 115656 -24395
rect 115748 -24439 115756 -24395
rect 115848 -24439 115856 -24395
rect 115948 -24439 115956 -24395
rect 116048 -24439 116056 -24395
rect 116148 -24439 116156 -24395
rect 116248 -24439 116256 -24395
rect 116348 -24439 116356 -24395
rect 116448 -24439 116456 -24395
rect 116548 -24439 116556 -24395
rect 116648 -24439 116656 -24395
rect 109104 -24495 109148 -24487
rect 109204 -24495 109248 -24487
rect 109304 -24495 109348 -24487
rect 109404 -24495 109448 -24487
rect 109504 -24495 109548 -24487
rect 109604 -24495 109648 -24487
rect 109704 -24495 109748 -24487
rect 109804 -24495 109848 -24487
rect 109904 -24495 109948 -24487
rect 110004 -24495 110048 -24487
rect 110104 -24495 110148 -24487
rect 110204 -24495 110248 -24487
rect 110304 -24495 110348 -24487
rect 110404 -24495 110448 -24487
rect 110504 -24495 110548 -24487
rect 110604 -24495 110648 -24487
rect 111104 -24495 111148 -24487
rect 111204 -24495 111248 -24487
rect 111304 -24495 111348 -24487
rect 111404 -24495 111448 -24487
rect 111504 -24495 111548 -24487
rect 111604 -24495 111648 -24487
rect 111704 -24495 111748 -24487
rect 111804 -24495 111848 -24487
rect 111904 -24495 111948 -24487
rect 112004 -24495 112048 -24487
rect 112104 -24495 112148 -24487
rect 112204 -24495 112248 -24487
rect 112304 -24495 112348 -24487
rect 112404 -24495 112448 -24487
rect 112504 -24495 112548 -24487
rect 112604 -24495 112648 -24487
rect 113104 -24495 113148 -24487
rect 113204 -24495 113248 -24487
rect 113304 -24495 113348 -24487
rect 113404 -24495 113448 -24487
rect 113504 -24495 113548 -24487
rect 113604 -24495 113648 -24487
rect 113704 -24495 113748 -24487
rect 113804 -24495 113848 -24487
rect 113904 -24495 113948 -24487
rect 114004 -24495 114048 -24487
rect 114104 -24495 114148 -24487
rect 114204 -24495 114248 -24487
rect 114304 -24495 114348 -24487
rect 114404 -24495 114448 -24487
rect 114504 -24495 114548 -24487
rect 114604 -24495 114648 -24487
rect 115104 -24495 115148 -24487
rect 115204 -24495 115248 -24487
rect 115304 -24495 115348 -24487
rect 115404 -24495 115448 -24487
rect 115504 -24495 115548 -24487
rect 115604 -24495 115648 -24487
rect 115704 -24495 115748 -24487
rect 115804 -24495 115848 -24487
rect 115904 -24495 115948 -24487
rect 116004 -24495 116048 -24487
rect 116104 -24495 116148 -24487
rect 116204 -24495 116248 -24487
rect 116304 -24495 116348 -24487
rect 116404 -24495 116448 -24487
rect 116504 -24495 116548 -24487
rect 116604 -24495 116648 -24487
rect 80849 -24526 80893 -24518
rect 80949 -24526 80993 -24518
rect 81049 -24526 81093 -24518
rect 81149 -24526 81193 -24518
rect 81249 -24526 81293 -24518
rect 81349 -24526 81393 -24518
rect 81449 -24526 81493 -24518
rect 81549 -24526 81593 -24518
rect 81649 -24526 81693 -24518
rect 81749 -24526 81793 -24518
rect 81849 -24526 81893 -24518
rect 81949 -24526 81993 -24518
rect 82049 -24526 82093 -24518
rect 82149 -24526 82193 -24518
rect 82249 -24526 82293 -24518
rect 82349 -24526 82393 -24518
rect 82849 -24526 82893 -24518
rect 82949 -24526 82993 -24518
rect 83049 -24526 83093 -24518
rect 83149 -24526 83193 -24518
rect 83249 -24526 83293 -24518
rect 83349 -24526 83393 -24518
rect 83449 -24526 83493 -24518
rect 83549 -24526 83593 -24518
rect 83649 -24526 83693 -24518
rect 83749 -24526 83793 -24518
rect 83849 -24526 83893 -24518
rect 83949 -24526 83993 -24518
rect 84049 -24526 84093 -24518
rect 84149 -24526 84193 -24518
rect 84249 -24526 84293 -24518
rect 84349 -24526 84393 -24518
rect 84849 -24526 84893 -24518
rect 84949 -24526 84993 -24518
rect 85049 -24526 85093 -24518
rect 85149 -24526 85193 -24518
rect 85249 -24526 85293 -24518
rect 85349 -24526 85393 -24518
rect 85449 -24526 85493 -24518
rect 85549 -24526 85593 -24518
rect 85649 -24526 85693 -24518
rect 85749 -24526 85793 -24518
rect 85849 -24526 85893 -24518
rect 85949 -24526 85993 -24518
rect 86049 -24526 86093 -24518
rect 86149 -24526 86193 -24518
rect 86249 -24526 86293 -24518
rect 86349 -24526 86393 -24518
rect 86849 -24526 86893 -24518
rect 86949 -24526 86993 -24518
rect 87049 -24526 87093 -24518
rect 87149 -24526 87193 -24518
rect 87249 -24526 87293 -24518
rect 87349 -24526 87393 -24518
rect 87449 -24526 87493 -24518
rect 87549 -24526 87593 -24518
rect 87649 -24526 87693 -24518
rect 87749 -24526 87793 -24518
rect 87849 -24526 87893 -24518
rect 87949 -24526 87993 -24518
rect 88049 -24526 88093 -24518
rect 88149 -24526 88193 -24518
rect 88249 -24526 88293 -24518
rect 88349 -24526 88393 -24518
rect 80893 -24570 80901 -24526
rect 80993 -24570 81001 -24526
rect 81093 -24570 81101 -24526
rect 81193 -24570 81201 -24526
rect 81293 -24570 81301 -24526
rect 81393 -24570 81401 -24526
rect 81493 -24570 81501 -24526
rect 81593 -24570 81601 -24526
rect 81693 -24570 81701 -24526
rect 81793 -24570 81801 -24526
rect 81893 -24570 81901 -24526
rect 81993 -24570 82001 -24526
rect 82093 -24570 82101 -24526
rect 82193 -24570 82201 -24526
rect 82293 -24570 82301 -24526
rect 82393 -24570 82401 -24526
rect 82893 -24570 82901 -24526
rect 82993 -24570 83001 -24526
rect 83093 -24570 83101 -24526
rect 83193 -24570 83201 -24526
rect 83293 -24570 83301 -24526
rect 83393 -24570 83401 -24526
rect 83493 -24570 83501 -24526
rect 83593 -24570 83601 -24526
rect 83693 -24570 83701 -24526
rect 83793 -24570 83801 -24526
rect 83893 -24570 83901 -24526
rect 83993 -24570 84001 -24526
rect 84093 -24570 84101 -24526
rect 84193 -24570 84201 -24526
rect 84293 -24570 84301 -24526
rect 84393 -24570 84401 -24526
rect 84893 -24570 84901 -24526
rect 84993 -24570 85001 -24526
rect 85093 -24570 85101 -24526
rect 85193 -24570 85201 -24526
rect 85293 -24570 85301 -24526
rect 85393 -24570 85401 -24526
rect 85493 -24570 85501 -24526
rect 85593 -24570 85601 -24526
rect 85693 -24570 85701 -24526
rect 85793 -24570 85801 -24526
rect 85893 -24570 85901 -24526
rect 85993 -24570 86001 -24526
rect 86093 -24570 86101 -24526
rect 86193 -24570 86201 -24526
rect 86293 -24570 86301 -24526
rect 86393 -24570 86401 -24526
rect 86893 -24570 86901 -24526
rect 86993 -24570 87001 -24526
rect 87093 -24570 87101 -24526
rect 87193 -24570 87201 -24526
rect 87293 -24570 87301 -24526
rect 87393 -24570 87401 -24526
rect 87493 -24570 87501 -24526
rect 87593 -24570 87601 -24526
rect 87693 -24570 87701 -24526
rect 87793 -24570 87801 -24526
rect 87893 -24570 87901 -24526
rect 87993 -24570 88001 -24526
rect 88093 -24570 88101 -24526
rect 88193 -24570 88201 -24526
rect 88293 -24570 88301 -24526
rect 88393 -24570 88401 -24526
rect 109148 -24539 109156 -24495
rect 109248 -24539 109256 -24495
rect 109348 -24539 109356 -24495
rect 109448 -24539 109456 -24495
rect 109548 -24539 109556 -24495
rect 109648 -24539 109656 -24495
rect 109748 -24539 109756 -24495
rect 109848 -24539 109856 -24495
rect 109948 -24539 109956 -24495
rect 110048 -24539 110056 -24495
rect 110148 -24539 110156 -24495
rect 110248 -24539 110256 -24495
rect 110348 -24539 110356 -24495
rect 110448 -24539 110456 -24495
rect 110548 -24539 110556 -24495
rect 110648 -24539 110656 -24495
rect 111148 -24539 111156 -24495
rect 111248 -24539 111256 -24495
rect 111348 -24539 111356 -24495
rect 111448 -24539 111456 -24495
rect 111548 -24539 111556 -24495
rect 111648 -24539 111656 -24495
rect 111748 -24539 111756 -24495
rect 111848 -24539 111856 -24495
rect 111948 -24539 111956 -24495
rect 112048 -24539 112056 -24495
rect 112148 -24539 112156 -24495
rect 112248 -24539 112256 -24495
rect 112348 -24539 112356 -24495
rect 112448 -24539 112456 -24495
rect 112548 -24539 112556 -24495
rect 112648 -24539 112656 -24495
rect 113148 -24539 113156 -24495
rect 113248 -24539 113256 -24495
rect 113348 -24539 113356 -24495
rect 113448 -24539 113456 -24495
rect 113548 -24539 113556 -24495
rect 113648 -24539 113656 -24495
rect 113748 -24539 113756 -24495
rect 113848 -24539 113856 -24495
rect 113948 -24539 113956 -24495
rect 114048 -24539 114056 -24495
rect 114148 -24539 114156 -24495
rect 114248 -24539 114256 -24495
rect 114348 -24539 114356 -24495
rect 114448 -24539 114456 -24495
rect 114548 -24539 114556 -24495
rect 114648 -24539 114656 -24495
rect 115148 -24539 115156 -24495
rect 115248 -24539 115256 -24495
rect 115348 -24539 115356 -24495
rect 115448 -24539 115456 -24495
rect 115548 -24539 115556 -24495
rect 115648 -24539 115656 -24495
rect 115748 -24539 115756 -24495
rect 115848 -24539 115856 -24495
rect 115948 -24539 115956 -24495
rect 116048 -24539 116056 -24495
rect 116148 -24539 116156 -24495
rect 116248 -24539 116256 -24495
rect 116348 -24539 116356 -24495
rect 116448 -24539 116456 -24495
rect 116548 -24539 116556 -24495
rect 116648 -24539 116656 -24495
rect 109104 -24595 109148 -24587
rect 109204 -24595 109248 -24587
rect 109304 -24595 109348 -24587
rect 109404 -24595 109448 -24587
rect 109504 -24595 109548 -24587
rect 109604 -24595 109648 -24587
rect 109704 -24595 109748 -24587
rect 109804 -24595 109848 -24587
rect 109904 -24595 109948 -24587
rect 110004 -24595 110048 -24587
rect 110104 -24595 110148 -24587
rect 110204 -24595 110248 -24587
rect 110304 -24595 110348 -24587
rect 110404 -24595 110448 -24587
rect 110504 -24595 110548 -24587
rect 110604 -24595 110648 -24587
rect 111104 -24595 111148 -24587
rect 111204 -24595 111248 -24587
rect 111304 -24595 111348 -24587
rect 111404 -24595 111448 -24587
rect 111504 -24595 111548 -24587
rect 111604 -24595 111648 -24587
rect 111704 -24595 111748 -24587
rect 111804 -24595 111848 -24587
rect 111904 -24595 111948 -24587
rect 112004 -24595 112048 -24587
rect 112104 -24595 112148 -24587
rect 112204 -24595 112248 -24587
rect 112304 -24595 112348 -24587
rect 112404 -24595 112448 -24587
rect 112504 -24595 112548 -24587
rect 112604 -24595 112648 -24587
rect 113104 -24595 113148 -24587
rect 113204 -24595 113248 -24587
rect 113304 -24595 113348 -24587
rect 113404 -24595 113448 -24587
rect 113504 -24595 113548 -24587
rect 113604 -24595 113648 -24587
rect 113704 -24595 113748 -24587
rect 113804 -24595 113848 -24587
rect 113904 -24595 113948 -24587
rect 114004 -24595 114048 -24587
rect 114104 -24595 114148 -24587
rect 114204 -24595 114248 -24587
rect 114304 -24595 114348 -24587
rect 114404 -24595 114448 -24587
rect 114504 -24595 114548 -24587
rect 114604 -24595 114648 -24587
rect 115104 -24595 115148 -24587
rect 115204 -24595 115248 -24587
rect 115304 -24595 115348 -24587
rect 115404 -24595 115448 -24587
rect 115504 -24595 115548 -24587
rect 115604 -24595 115648 -24587
rect 115704 -24595 115748 -24587
rect 115804 -24595 115848 -24587
rect 115904 -24595 115948 -24587
rect 116004 -24595 116048 -24587
rect 116104 -24595 116148 -24587
rect 116204 -24595 116248 -24587
rect 116304 -24595 116348 -24587
rect 116404 -24595 116448 -24587
rect 116504 -24595 116548 -24587
rect 116604 -24595 116648 -24587
rect 80849 -24626 80893 -24618
rect 80949 -24626 80993 -24618
rect 81049 -24626 81093 -24618
rect 81149 -24626 81193 -24618
rect 81249 -24626 81293 -24618
rect 81349 -24626 81393 -24618
rect 81449 -24626 81493 -24618
rect 81549 -24626 81593 -24618
rect 81649 -24626 81693 -24618
rect 81749 -24626 81793 -24618
rect 81849 -24626 81893 -24618
rect 81949 -24626 81993 -24618
rect 82049 -24626 82093 -24618
rect 82149 -24626 82193 -24618
rect 82249 -24626 82293 -24618
rect 82349 -24626 82393 -24618
rect 82849 -24626 82893 -24618
rect 82949 -24626 82993 -24618
rect 83049 -24626 83093 -24618
rect 83149 -24626 83193 -24618
rect 83249 -24626 83293 -24618
rect 83349 -24626 83393 -24618
rect 83449 -24626 83493 -24618
rect 83549 -24626 83593 -24618
rect 83649 -24626 83693 -24618
rect 83749 -24626 83793 -24618
rect 83849 -24626 83893 -24618
rect 83949 -24626 83993 -24618
rect 84049 -24626 84093 -24618
rect 84149 -24626 84193 -24618
rect 84249 -24626 84293 -24618
rect 84349 -24626 84393 -24618
rect 84849 -24626 84893 -24618
rect 84949 -24626 84993 -24618
rect 85049 -24626 85093 -24618
rect 85149 -24626 85193 -24618
rect 85249 -24626 85293 -24618
rect 85349 -24626 85393 -24618
rect 85449 -24626 85493 -24618
rect 85549 -24626 85593 -24618
rect 85649 -24626 85693 -24618
rect 85749 -24626 85793 -24618
rect 85849 -24626 85893 -24618
rect 85949 -24626 85993 -24618
rect 86049 -24626 86093 -24618
rect 86149 -24626 86193 -24618
rect 86249 -24626 86293 -24618
rect 86349 -24626 86393 -24618
rect 86849 -24626 86893 -24618
rect 86949 -24626 86993 -24618
rect 87049 -24626 87093 -24618
rect 87149 -24626 87193 -24618
rect 87249 -24626 87293 -24618
rect 87349 -24626 87393 -24618
rect 87449 -24626 87493 -24618
rect 87549 -24626 87593 -24618
rect 87649 -24626 87693 -24618
rect 87749 -24626 87793 -24618
rect 87849 -24626 87893 -24618
rect 87949 -24626 87993 -24618
rect 88049 -24626 88093 -24618
rect 88149 -24626 88193 -24618
rect 88249 -24626 88293 -24618
rect 88349 -24626 88393 -24618
rect 80893 -24670 80901 -24626
rect 80993 -24670 81001 -24626
rect 81093 -24670 81101 -24626
rect 81193 -24670 81201 -24626
rect 81293 -24670 81301 -24626
rect 81393 -24670 81401 -24626
rect 81493 -24670 81501 -24626
rect 81593 -24670 81601 -24626
rect 81693 -24670 81701 -24626
rect 81793 -24670 81801 -24626
rect 81893 -24670 81901 -24626
rect 81993 -24670 82001 -24626
rect 82093 -24670 82101 -24626
rect 82193 -24670 82201 -24626
rect 82293 -24670 82301 -24626
rect 82393 -24670 82401 -24626
rect 82893 -24670 82901 -24626
rect 82993 -24670 83001 -24626
rect 83093 -24670 83101 -24626
rect 83193 -24670 83201 -24626
rect 83293 -24670 83301 -24626
rect 83393 -24670 83401 -24626
rect 83493 -24670 83501 -24626
rect 83593 -24670 83601 -24626
rect 83693 -24670 83701 -24626
rect 83793 -24670 83801 -24626
rect 83893 -24670 83901 -24626
rect 83993 -24670 84001 -24626
rect 84093 -24670 84101 -24626
rect 84193 -24670 84201 -24626
rect 84293 -24670 84301 -24626
rect 84393 -24670 84401 -24626
rect 84893 -24670 84901 -24626
rect 84993 -24670 85001 -24626
rect 85093 -24670 85101 -24626
rect 85193 -24670 85201 -24626
rect 85293 -24670 85301 -24626
rect 85393 -24670 85401 -24626
rect 85493 -24670 85501 -24626
rect 85593 -24670 85601 -24626
rect 85693 -24670 85701 -24626
rect 85793 -24670 85801 -24626
rect 85893 -24670 85901 -24626
rect 85993 -24670 86001 -24626
rect 86093 -24670 86101 -24626
rect 86193 -24670 86201 -24626
rect 86293 -24670 86301 -24626
rect 86393 -24670 86401 -24626
rect 86893 -24670 86901 -24626
rect 86993 -24670 87001 -24626
rect 87093 -24670 87101 -24626
rect 87193 -24670 87201 -24626
rect 87293 -24670 87301 -24626
rect 87393 -24670 87401 -24626
rect 87493 -24670 87501 -24626
rect 87593 -24670 87601 -24626
rect 87693 -24670 87701 -24626
rect 87793 -24670 87801 -24626
rect 87893 -24670 87901 -24626
rect 87993 -24670 88001 -24626
rect 88093 -24670 88101 -24626
rect 88193 -24670 88201 -24626
rect 88293 -24670 88301 -24626
rect 88393 -24670 88401 -24626
rect 109148 -24639 109156 -24595
rect 109248 -24639 109256 -24595
rect 109348 -24639 109356 -24595
rect 109448 -24639 109456 -24595
rect 109548 -24639 109556 -24595
rect 109648 -24639 109656 -24595
rect 109748 -24639 109756 -24595
rect 109848 -24639 109856 -24595
rect 109948 -24639 109956 -24595
rect 110048 -24639 110056 -24595
rect 110148 -24639 110156 -24595
rect 110248 -24639 110256 -24595
rect 110348 -24639 110356 -24595
rect 110448 -24639 110456 -24595
rect 110548 -24639 110556 -24595
rect 110648 -24639 110656 -24595
rect 111148 -24639 111156 -24595
rect 111248 -24639 111256 -24595
rect 111348 -24639 111356 -24595
rect 111448 -24639 111456 -24595
rect 111548 -24639 111556 -24595
rect 111648 -24639 111656 -24595
rect 111748 -24639 111756 -24595
rect 111848 -24639 111856 -24595
rect 111948 -24639 111956 -24595
rect 112048 -24639 112056 -24595
rect 112148 -24639 112156 -24595
rect 112248 -24639 112256 -24595
rect 112348 -24639 112356 -24595
rect 112448 -24639 112456 -24595
rect 112548 -24639 112556 -24595
rect 112648 -24639 112656 -24595
rect 113148 -24639 113156 -24595
rect 113248 -24639 113256 -24595
rect 113348 -24639 113356 -24595
rect 113448 -24639 113456 -24595
rect 113548 -24639 113556 -24595
rect 113648 -24639 113656 -24595
rect 113748 -24639 113756 -24595
rect 113848 -24639 113856 -24595
rect 113948 -24639 113956 -24595
rect 114048 -24639 114056 -24595
rect 114148 -24639 114156 -24595
rect 114248 -24639 114256 -24595
rect 114348 -24639 114356 -24595
rect 114448 -24639 114456 -24595
rect 114548 -24639 114556 -24595
rect 114648 -24639 114656 -24595
rect 115148 -24639 115156 -24595
rect 115248 -24639 115256 -24595
rect 115348 -24639 115356 -24595
rect 115448 -24639 115456 -24595
rect 115548 -24639 115556 -24595
rect 115648 -24639 115656 -24595
rect 115748 -24639 115756 -24595
rect 115848 -24639 115856 -24595
rect 115948 -24639 115956 -24595
rect 116048 -24639 116056 -24595
rect 116148 -24639 116156 -24595
rect 116248 -24639 116256 -24595
rect 116348 -24639 116356 -24595
rect 116448 -24639 116456 -24595
rect 116548 -24639 116556 -24595
rect 116648 -24639 116656 -24595
rect 109104 -24695 109148 -24687
rect 109204 -24695 109248 -24687
rect 109304 -24695 109348 -24687
rect 109404 -24695 109448 -24687
rect 109504 -24695 109548 -24687
rect 109604 -24695 109648 -24687
rect 109704 -24695 109748 -24687
rect 109804 -24695 109848 -24687
rect 109904 -24695 109948 -24687
rect 110004 -24695 110048 -24687
rect 110104 -24695 110148 -24687
rect 110204 -24695 110248 -24687
rect 110304 -24695 110348 -24687
rect 110404 -24695 110448 -24687
rect 110504 -24695 110548 -24687
rect 110604 -24695 110648 -24687
rect 111104 -24695 111148 -24687
rect 111204 -24695 111248 -24687
rect 111304 -24695 111348 -24687
rect 111404 -24695 111448 -24687
rect 111504 -24695 111548 -24687
rect 111604 -24695 111648 -24687
rect 111704 -24695 111748 -24687
rect 111804 -24695 111848 -24687
rect 111904 -24695 111948 -24687
rect 112004 -24695 112048 -24687
rect 112104 -24695 112148 -24687
rect 112204 -24695 112248 -24687
rect 112304 -24695 112348 -24687
rect 112404 -24695 112448 -24687
rect 112504 -24695 112548 -24687
rect 112604 -24695 112648 -24687
rect 113104 -24695 113148 -24687
rect 113204 -24695 113248 -24687
rect 113304 -24695 113348 -24687
rect 113404 -24695 113448 -24687
rect 113504 -24695 113548 -24687
rect 113604 -24695 113648 -24687
rect 113704 -24695 113748 -24687
rect 113804 -24695 113848 -24687
rect 113904 -24695 113948 -24687
rect 114004 -24695 114048 -24687
rect 114104 -24695 114148 -24687
rect 114204 -24695 114248 -24687
rect 114304 -24695 114348 -24687
rect 114404 -24695 114448 -24687
rect 114504 -24695 114548 -24687
rect 114604 -24695 114648 -24687
rect 115104 -24695 115148 -24687
rect 115204 -24695 115248 -24687
rect 115304 -24695 115348 -24687
rect 115404 -24695 115448 -24687
rect 115504 -24695 115548 -24687
rect 115604 -24695 115648 -24687
rect 115704 -24695 115748 -24687
rect 115804 -24695 115848 -24687
rect 115904 -24695 115948 -24687
rect 116004 -24695 116048 -24687
rect 116104 -24695 116148 -24687
rect 116204 -24695 116248 -24687
rect 116304 -24695 116348 -24687
rect 116404 -24695 116448 -24687
rect 116504 -24695 116548 -24687
rect 116604 -24695 116648 -24687
rect 80849 -24726 80893 -24718
rect 80949 -24726 80993 -24718
rect 81049 -24726 81093 -24718
rect 81149 -24726 81193 -24718
rect 81249 -24726 81293 -24718
rect 81349 -24726 81393 -24718
rect 81449 -24726 81493 -24718
rect 81549 -24726 81593 -24718
rect 81649 -24726 81693 -24718
rect 81749 -24726 81793 -24718
rect 81849 -24726 81893 -24718
rect 81949 -24726 81993 -24718
rect 82049 -24726 82093 -24718
rect 82149 -24726 82193 -24718
rect 82249 -24726 82293 -24718
rect 82349 -24726 82393 -24718
rect 82849 -24726 82893 -24718
rect 82949 -24726 82993 -24718
rect 83049 -24726 83093 -24718
rect 83149 -24726 83193 -24718
rect 83249 -24726 83293 -24718
rect 83349 -24726 83393 -24718
rect 83449 -24726 83493 -24718
rect 83549 -24726 83593 -24718
rect 83649 -24726 83693 -24718
rect 83749 -24726 83793 -24718
rect 83849 -24726 83893 -24718
rect 83949 -24726 83993 -24718
rect 84049 -24726 84093 -24718
rect 84149 -24726 84193 -24718
rect 84249 -24726 84293 -24718
rect 84349 -24726 84393 -24718
rect 84849 -24726 84893 -24718
rect 84949 -24726 84993 -24718
rect 85049 -24726 85093 -24718
rect 85149 -24726 85193 -24718
rect 85249 -24726 85293 -24718
rect 85349 -24726 85393 -24718
rect 85449 -24726 85493 -24718
rect 85549 -24726 85593 -24718
rect 85649 -24726 85693 -24718
rect 85749 -24726 85793 -24718
rect 85849 -24726 85893 -24718
rect 85949 -24726 85993 -24718
rect 86049 -24726 86093 -24718
rect 86149 -24726 86193 -24718
rect 86249 -24726 86293 -24718
rect 86349 -24726 86393 -24718
rect 86849 -24726 86893 -24718
rect 86949 -24726 86993 -24718
rect 87049 -24726 87093 -24718
rect 87149 -24726 87193 -24718
rect 87249 -24726 87293 -24718
rect 87349 -24726 87393 -24718
rect 87449 -24726 87493 -24718
rect 87549 -24726 87593 -24718
rect 87649 -24726 87693 -24718
rect 87749 -24726 87793 -24718
rect 87849 -24726 87893 -24718
rect 87949 -24726 87993 -24718
rect 88049 -24726 88093 -24718
rect 88149 -24726 88193 -24718
rect 88249 -24726 88293 -24718
rect 88349 -24726 88393 -24718
rect 80893 -24770 80901 -24726
rect 80993 -24770 81001 -24726
rect 81093 -24770 81101 -24726
rect 81193 -24770 81201 -24726
rect 81293 -24770 81301 -24726
rect 81393 -24770 81401 -24726
rect 81493 -24770 81501 -24726
rect 81593 -24770 81601 -24726
rect 81693 -24770 81701 -24726
rect 81793 -24770 81801 -24726
rect 81893 -24770 81901 -24726
rect 81993 -24770 82001 -24726
rect 82093 -24770 82101 -24726
rect 82193 -24770 82201 -24726
rect 82293 -24770 82301 -24726
rect 82393 -24770 82401 -24726
rect 82893 -24770 82901 -24726
rect 82993 -24770 83001 -24726
rect 83093 -24770 83101 -24726
rect 83193 -24770 83201 -24726
rect 83293 -24770 83301 -24726
rect 83393 -24770 83401 -24726
rect 83493 -24770 83501 -24726
rect 83593 -24770 83601 -24726
rect 83693 -24770 83701 -24726
rect 83793 -24770 83801 -24726
rect 83893 -24770 83901 -24726
rect 83993 -24770 84001 -24726
rect 84093 -24770 84101 -24726
rect 84193 -24770 84201 -24726
rect 84293 -24770 84301 -24726
rect 84393 -24770 84401 -24726
rect 84893 -24770 84901 -24726
rect 84993 -24770 85001 -24726
rect 85093 -24770 85101 -24726
rect 85193 -24770 85201 -24726
rect 85293 -24770 85301 -24726
rect 85393 -24770 85401 -24726
rect 85493 -24770 85501 -24726
rect 85593 -24770 85601 -24726
rect 85693 -24770 85701 -24726
rect 85793 -24770 85801 -24726
rect 85893 -24770 85901 -24726
rect 85993 -24770 86001 -24726
rect 86093 -24770 86101 -24726
rect 86193 -24770 86201 -24726
rect 86293 -24770 86301 -24726
rect 86393 -24770 86401 -24726
rect 86893 -24770 86901 -24726
rect 86993 -24770 87001 -24726
rect 87093 -24770 87101 -24726
rect 87193 -24770 87201 -24726
rect 87293 -24770 87301 -24726
rect 87393 -24770 87401 -24726
rect 87493 -24770 87501 -24726
rect 87593 -24770 87601 -24726
rect 87693 -24770 87701 -24726
rect 87793 -24770 87801 -24726
rect 87893 -24770 87901 -24726
rect 87993 -24770 88001 -24726
rect 88093 -24770 88101 -24726
rect 88193 -24770 88201 -24726
rect 88293 -24770 88301 -24726
rect 88393 -24770 88401 -24726
rect 109148 -24739 109156 -24695
rect 109248 -24739 109256 -24695
rect 109348 -24739 109356 -24695
rect 109448 -24739 109456 -24695
rect 109548 -24739 109556 -24695
rect 109648 -24739 109656 -24695
rect 109748 -24739 109756 -24695
rect 109848 -24739 109856 -24695
rect 109948 -24739 109956 -24695
rect 110048 -24739 110056 -24695
rect 110148 -24739 110156 -24695
rect 110248 -24739 110256 -24695
rect 110348 -24739 110356 -24695
rect 110448 -24739 110456 -24695
rect 110548 -24739 110556 -24695
rect 110648 -24739 110656 -24695
rect 111148 -24739 111156 -24695
rect 111248 -24739 111256 -24695
rect 111348 -24739 111356 -24695
rect 111448 -24739 111456 -24695
rect 111548 -24739 111556 -24695
rect 111648 -24739 111656 -24695
rect 111748 -24739 111756 -24695
rect 111848 -24739 111856 -24695
rect 111948 -24739 111956 -24695
rect 112048 -24739 112056 -24695
rect 112148 -24739 112156 -24695
rect 112248 -24739 112256 -24695
rect 112348 -24739 112356 -24695
rect 112448 -24739 112456 -24695
rect 112548 -24739 112556 -24695
rect 112648 -24739 112656 -24695
rect 113148 -24739 113156 -24695
rect 113248 -24739 113256 -24695
rect 113348 -24739 113356 -24695
rect 113448 -24739 113456 -24695
rect 113548 -24739 113556 -24695
rect 113648 -24739 113656 -24695
rect 113748 -24739 113756 -24695
rect 113848 -24739 113856 -24695
rect 113948 -24739 113956 -24695
rect 114048 -24739 114056 -24695
rect 114148 -24739 114156 -24695
rect 114248 -24739 114256 -24695
rect 114348 -24739 114356 -24695
rect 114448 -24739 114456 -24695
rect 114548 -24739 114556 -24695
rect 114648 -24739 114656 -24695
rect 115148 -24739 115156 -24695
rect 115248 -24739 115256 -24695
rect 115348 -24739 115356 -24695
rect 115448 -24739 115456 -24695
rect 115548 -24739 115556 -24695
rect 115648 -24739 115656 -24695
rect 115748 -24739 115756 -24695
rect 115848 -24739 115856 -24695
rect 115948 -24739 115956 -24695
rect 116048 -24739 116056 -24695
rect 116148 -24739 116156 -24695
rect 116248 -24739 116256 -24695
rect 116348 -24739 116356 -24695
rect 116448 -24739 116456 -24695
rect 116548 -24739 116556 -24695
rect 116648 -24739 116656 -24695
rect 109104 -24795 109148 -24787
rect 109204 -24795 109248 -24787
rect 109304 -24795 109348 -24787
rect 109404 -24795 109448 -24787
rect 109504 -24795 109548 -24787
rect 109604 -24795 109648 -24787
rect 109704 -24795 109748 -24787
rect 109804 -24795 109848 -24787
rect 109904 -24795 109948 -24787
rect 110004 -24795 110048 -24787
rect 110104 -24795 110148 -24787
rect 110204 -24795 110248 -24787
rect 110304 -24795 110348 -24787
rect 110404 -24795 110448 -24787
rect 110504 -24795 110548 -24787
rect 110604 -24795 110648 -24787
rect 111104 -24795 111148 -24787
rect 111204 -24795 111248 -24787
rect 111304 -24795 111348 -24787
rect 111404 -24795 111448 -24787
rect 111504 -24795 111548 -24787
rect 111604 -24795 111648 -24787
rect 111704 -24795 111748 -24787
rect 111804 -24795 111848 -24787
rect 111904 -24795 111948 -24787
rect 112004 -24795 112048 -24787
rect 112104 -24795 112148 -24787
rect 112204 -24795 112248 -24787
rect 112304 -24795 112348 -24787
rect 112404 -24795 112448 -24787
rect 112504 -24795 112548 -24787
rect 112604 -24795 112648 -24787
rect 113104 -24795 113148 -24787
rect 113204 -24795 113248 -24787
rect 113304 -24795 113348 -24787
rect 113404 -24795 113448 -24787
rect 113504 -24795 113548 -24787
rect 113604 -24795 113648 -24787
rect 113704 -24795 113748 -24787
rect 113804 -24795 113848 -24787
rect 113904 -24795 113948 -24787
rect 114004 -24795 114048 -24787
rect 114104 -24795 114148 -24787
rect 114204 -24795 114248 -24787
rect 114304 -24795 114348 -24787
rect 114404 -24795 114448 -24787
rect 114504 -24795 114548 -24787
rect 114604 -24795 114648 -24787
rect 115104 -24795 115148 -24787
rect 115204 -24795 115248 -24787
rect 115304 -24795 115348 -24787
rect 115404 -24795 115448 -24787
rect 115504 -24795 115548 -24787
rect 115604 -24795 115648 -24787
rect 115704 -24795 115748 -24787
rect 115804 -24795 115848 -24787
rect 115904 -24795 115948 -24787
rect 116004 -24795 116048 -24787
rect 116104 -24795 116148 -24787
rect 116204 -24795 116248 -24787
rect 116304 -24795 116348 -24787
rect 116404 -24795 116448 -24787
rect 116504 -24795 116548 -24787
rect 116604 -24795 116648 -24787
rect 80849 -24826 80893 -24818
rect 80949 -24826 80993 -24818
rect 81049 -24826 81093 -24818
rect 81149 -24826 81193 -24818
rect 81249 -24826 81293 -24818
rect 81349 -24826 81393 -24818
rect 81449 -24826 81493 -24818
rect 81549 -24826 81593 -24818
rect 81649 -24826 81693 -24818
rect 81749 -24826 81793 -24818
rect 81849 -24826 81893 -24818
rect 81949 -24826 81993 -24818
rect 82049 -24826 82093 -24818
rect 82149 -24826 82193 -24818
rect 82249 -24826 82293 -24818
rect 82349 -24826 82393 -24818
rect 82849 -24826 82893 -24818
rect 82949 -24826 82993 -24818
rect 83049 -24826 83093 -24818
rect 83149 -24826 83193 -24818
rect 83249 -24826 83293 -24818
rect 83349 -24826 83393 -24818
rect 83449 -24826 83493 -24818
rect 83549 -24826 83593 -24818
rect 83649 -24826 83693 -24818
rect 83749 -24826 83793 -24818
rect 83849 -24826 83893 -24818
rect 83949 -24826 83993 -24818
rect 84049 -24826 84093 -24818
rect 84149 -24826 84193 -24818
rect 84249 -24826 84293 -24818
rect 84349 -24826 84393 -24818
rect 84849 -24826 84893 -24818
rect 84949 -24826 84993 -24818
rect 85049 -24826 85093 -24818
rect 85149 -24826 85193 -24818
rect 85249 -24826 85293 -24818
rect 85349 -24826 85393 -24818
rect 85449 -24826 85493 -24818
rect 85549 -24826 85593 -24818
rect 85649 -24826 85693 -24818
rect 85749 -24826 85793 -24818
rect 85849 -24826 85893 -24818
rect 85949 -24826 85993 -24818
rect 86049 -24826 86093 -24818
rect 86149 -24826 86193 -24818
rect 86249 -24826 86293 -24818
rect 86349 -24826 86393 -24818
rect 86849 -24826 86893 -24818
rect 86949 -24826 86993 -24818
rect 87049 -24826 87093 -24818
rect 87149 -24826 87193 -24818
rect 87249 -24826 87293 -24818
rect 87349 -24826 87393 -24818
rect 87449 -24826 87493 -24818
rect 87549 -24826 87593 -24818
rect 87649 -24826 87693 -24818
rect 87749 -24826 87793 -24818
rect 87849 -24826 87893 -24818
rect 87949 -24826 87993 -24818
rect 88049 -24826 88093 -24818
rect 88149 -24826 88193 -24818
rect 88249 -24826 88293 -24818
rect 88349 -24826 88393 -24818
rect 80893 -24870 80901 -24826
rect 80993 -24870 81001 -24826
rect 81093 -24870 81101 -24826
rect 81193 -24870 81201 -24826
rect 81293 -24870 81301 -24826
rect 81393 -24870 81401 -24826
rect 81493 -24870 81501 -24826
rect 81593 -24870 81601 -24826
rect 81693 -24870 81701 -24826
rect 81793 -24870 81801 -24826
rect 81893 -24870 81901 -24826
rect 81993 -24870 82001 -24826
rect 82093 -24870 82101 -24826
rect 82193 -24870 82201 -24826
rect 82293 -24870 82301 -24826
rect 82393 -24870 82401 -24826
rect 82893 -24870 82901 -24826
rect 82993 -24870 83001 -24826
rect 83093 -24870 83101 -24826
rect 83193 -24870 83201 -24826
rect 83293 -24870 83301 -24826
rect 83393 -24870 83401 -24826
rect 83493 -24870 83501 -24826
rect 83593 -24870 83601 -24826
rect 83693 -24870 83701 -24826
rect 83793 -24870 83801 -24826
rect 83893 -24870 83901 -24826
rect 83993 -24870 84001 -24826
rect 84093 -24870 84101 -24826
rect 84193 -24870 84201 -24826
rect 84293 -24870 84301 -24826
rect 84393 -24870 84401 -24826
rect 84893 -24870 84901 -24826
rect 84993 -24870 85001 -24826
rect 85093 -24870 85101 -24826
rect 85193 -24870 85201 -24826
rect 85293 -24870 85301 -24826
rect 85393 -24870 85401 -24826
rect 85493 -24870 85501 -24826
rect 85593 -24870 85601 -24826
rect 85693 -24870 85701 -24826
rect 85793 -24870 85801 -24826
rect 85893 -24870 85901 -24826
rect 85993 -24870 86001 -24826
rect 86093 -24870 86101 -24826
rect 86193 -24870 86201 -24826
rect 86293 -24870 86301 -24826
rect 86393 -24870 86401 -24826
rect 86893 -24870 86901 -24826
rect 86993 -24870 87001 -24826
rect 87093 -24870 87101 -24826
rect 87193 -24870 87201 -24826
rect 87293 -24870 87301 -24826
rect 87393 -24870 87401 -24826
rect 87493 -24870 87501 -24826
rect 87593 -24870 87601 -24826
rect 87693 -24870 87701 -24826
rect 87793 -24870 87801 -24826
rect 87893 -24870 87901 -24826
rect 87993 -24870 88001 -24826
rect 88093 -24870 88101 -24826
rect 88193 -24870 88201 -24826
rect 88293 -24870 88301 -24826
rect 88393 -24870 88401 -24826
rect 109148 -24839 109156 -24795
rect 109248 -24839 109256 -24795
rect 109348 -24839 109356 -24795
rect 109448 -24839 109456 -24795
rect 109548 -24839 109556 -24795
rect 109648 -24839 109656 -24795
rect 109748 -24839 109756 -24795
rect 109848 -24839 109856 -24795
rect 109948 -24839 109956 -24795
rect 110048 -24839 110056 -24795
rect 110148 -24839 110156 -24795
rect 110248 -24839 110256 -24795
rect 110348 -24839 110356 -24795
rect 110448 -24839 110456 -24795
rect 110548 -24839 110556 -24795
rect 110648 -24839 110656 -24795
rect 111148 -24839 111156 -24795
rect 111248 -24839 111256 -24795
rect 111348 -24839 111356 -24795
rect 111448 -24839 111456 -24795
rect 111548 -24839 111556 -24795
rect 111648 -24839 111656 -24795
rect 111748 -24839 111756 -24795
rect 111848 -24839 111856 -24795
rect 111948 -24839 111956 -24795
rect 112048 -24839 112056 -24795
rect 112148 -24839 112156 -24795
rect 112248 -24839 112256 -24795
rect 112348 -24839 112356 -24795
rect 112448 -24839 112456 -24795
rect 112548 -24839 112556 -24795
rect 112648 -24839 112656 -24795
rect 113148 -24839 113156 -24795
rect 113248 -24839 113256 -24795
rect 113348 -24839 113356 -24795
rect 113448 -24839 113456 -24795
rect 113548 -24839 113556 -24795
rect 113648 -24839 113656 -24795
rect 113748 -24839 113756 -24795
rect 113848 -24839 113856 -24795
rect 113948 -24839 113956 -24795
rect 114048 -24839 114056 -24795
rect 114148 -24839 114156 -24795
rect 114248 -24839 114256 -24795
rect 114348 -24839 114356 -24795
rect 114448 -24839 114456 -24795
rect 114548 -24839 114556 -24795
rect 114648 -24839 114656 -24795
rect 115148 -24839 115156 -24795
rect 115248 -24839 115256 -24795
rect 115348 -24839 115356 -24795
rect 115448 -24839 115456 -24795
rect 115548 -24839 115556 -24795
rect 115648 -24839 115656 -24795
rect 115748 -24839 115756 -24795
rect 115848 -24839 115856 -24795
rect 115948 -24839 115956 -24795
rect 116048 -24839 116056 -24795
rect 116148 -24839 116156 -24795
rect 116248 -24839 116256 -24795
rect 116348 -24839 116356 -24795
rect 116448 -24839 116456 -24795
rect 116548 -24839 116556 -24795
rect 116648 -24839 116656 -24795
rect 109104 -24895 109148 -24887
rect 109204 -24895 109248 -24887
rect 109304 -24895 109348 -24887
rect 109404 -24895 109448 -24887
rect 109504 -24895 109548 -24887
rect 109604 -24895 109648 -24887
rect 109704 -24895 109748 -24887
rect 109804 -24895 109848 -24887
rect 109904 -24895 109948 -24887
rect 110004 -24895 110048 -24887
rect 110104 -24895 110148 -24887
rect 110204 -24895 110248 -24887
rect 110304 -24895 110348 -24887
rect 110404 -24895 110448 -24887
rect 110504 -24895 110548 -24887
rect 110604 -24895 110648 -24887
rect 111104 -24895 111148 -24887
rect 111204 -24895 111248 -24887
rect 111304 -24895 111348 -24887
rect 111404 -24895 111448 -24887
rect 111504 -24895 111548 -24887
rect 111604 -24895 111648 -24887
rect 111704 -24895 111748 -24887
rect 111804 -24895 111848 -24887
rect 111904 -24895 111948 -24887
rect 112004 -24895 112048 -24887
rect 112104 -24895 112148 -24887
rect 112204 -24895 112248 -24887
rect 112304 -24895 112348 -24887
rect 112404 -24895 112448 -24887
rect 112504 -24895 112548 -24887
rect 112604 -24895 112648 -24887
rect 113104 -24895 113148 -24887
rect 113204 -24895 113248 -24887
rect 113304 -24895 113348 -24887
rect 113404 -24895 113448 -24887
rect 113504 -24895 113548 -24887
rect 113604 -24895 113648 -24887
rect 113704 -24895 113748 -24887
rect 113804 -24895 113848 -24887
rect 113904 -24895 113948 -24887
rect 114004 -24895 114048 -24887
rect 114104 -24895 114148 -24887
rect 114204 -24895 114248 -24887
rect 114304 -24895 114348 -24887
rect 114404 -24895 114448 -24887
rect 114504 -24895 114548 -24887
rect 114604 -24895 114648 -24887
rect 115104 -24895 115148 -24887
rect 115204 -24895 115248 -24887
rect 115304 -24895 115348 -24887
rect 115404 -24895 115448 -24887
rect 115504 -24895 115548 -24887
rect 115604 -24895 115648 -24887
rect 115704 -24895 115748 -24887
rect 115804 -24895 115848 -24887
rect 115904 -24895 115948 -24887
rect 116004 -24895 116048 -24887
rect 116104 -24895 116148 -24887
rect 116204 -24895 116248 -24887
rect 116304 -24895 116348 -24887
rect 116404 -24895 116448 -24887
rect 116504 -24895 116548 -24887
rect 116604 -24895 116648 -24887
rect 80849 -24926 80893 -24918
rect 80949 -24926 80993 -24918
rect 81049 -24926 81093 -24918
rect 81149 -24926 81193 -24918
rect 81249 -24926 81293 -24918
rect 81349 -24926 81393 -24918
rect 81449 -24926 81493 -24918
rect 81549 -24926 81593 -24918
rect 81649 -24926 81693 -24918
rect 81749 -24926 81793 -24918
rect 81849 -24926 81893 -24918
rect 81949 -24926 81993 -24918
rect 82049 -24926 82093 -24918
rect 82149 -24926 82193 -24918
rect 82249 -24926 82293 -24918
rect 82349 -24926 82393 -24918
rect 82849 -24926 82893 -24918
rect 82949 -24926 82993 -24918
rect 83049 -24926 83093 -24918
rect 83149 -24926 83193 -24918
rect 83249 -24926 83293 -24918
rect 83349 -24926 83393 -24918
rect 83449 -24926 83493 -24918
rect 83549 -24926 83593 -24918
rect 83649 -24926 83693 -24918
rect 83749 -24926 83793 -24918
rect 83849 -24926 83893 -24918
rect 83949 -24926 83993 -24918
rect 84049 -24926 84093 -24918
rect 84149 -24926 84193 -24918
rect 84249 -24926 84293 -24918
rect 84349 -24926 84393 -24918
rect 84849 -24926 84893 -24918
rect 84949 -24926 84993 -24918
rect 85049 -24926 85093 -24918
rect 85149 -24926 85193 -24918
rect 85249 -24926 85293 -24918
rect 85349 -24926 85393 -24918
rect 85449 -24926 85493 -24918
rect 85549 -24926 85593 -24918
rect 85649 -24926 85693 -24918
rect 85749 -24926 85793 -24918
rect 85849 -24926 85893 -24918
rect 85949 -24926 85993 -24918
rect 86049 -24926 86093 -24918
rect 86149 -24926 86193 -24918
rect 86249 -24926 86293 -24918
rect 86349 -24926 86393 -24918
rect 86849 -24926 86893 -24918
rect 86949 -24926 86993 -24918
rect 87049 -24926 87093 -24918
rect 87149 -24926 87193 -24918
rect 87249 -24926 87293 -24918
rect 87349 -24926 87393 -24918
rect 87449 -24926 87493 -24918
rect 87549 -24926 87593 -24918
rect 87649 -24926 87693 -24918
rect 87749 -24926 87793 -24918
rect 87849 -24926 87893 -24918
rect 87949 -24926 87993 -24918
rect 88049 -24926 88093 -24918
rect 88149 -24926 88193 -24918
rect 88249 -24926 88293 -24918
rect 88349 -24926 88393 -24918
rect 80893 -24970 80901 -24926
rect 80993 -24970 81001 -24926
rect 81093 -24970 81101 -24926
rect 81193 -24970 81201 -24926
rect 81293 -24970 81301 -24926
rect 81393 -24970 81401 -24926
rect 81493 -24970 81501 -24926
rect 81593 -24970 81601 -24926
rect 81693 -24970 81701 -24926
rect 81793 -24970 81801 -24926
rect 81893 -24970 81901 -24926
rect 81993 -24970 82001 -24926
rect 82093 -24970 82101 -24926
rect 82193 -24970 82201 -24926
rect 82293 -24970 82301 -24926
rect 82393 -24970 82401 -24926
rect 82893 -24970 82901 -24926
rect 82993 -24970 83001 -24926
rect 83093 -24970 83101 -24926
rect 83193 -24970 83201 -24926
rect 83293 -24970 83301 -24926
rect 83393 -24970 83401 -24926
rect 83493 -24970 83501 -24926
rect 83593 -24970 83601 -24926
rect 83693 -24970 83701 -24926
rect 83793 -24970 83801 -24926
rect 83893 -24970 83901 -24926
rect 83993 -24970 84001 -24926
rect 84093 -24970 84101 -24926
rect 84193 -24970 84201 -24926
rect 84293 -24970 84301 -24926
rect 84393 -24970 84401 -24926
rect 84893 -24970 84901 -24926
rect 84993 -24970 85001 -24926
rect 85093 -24970 85101 -24926
rect 85193 -24970 85201 -24926
rect 85293 -24970 85301 -24926
rect 85393 -24970 85401 -24926
rect 85493 -24970 85501 -24926
rect 85593 -24970 85601 -24926
rect 85693 -24970 85701 -24926
rect 85793 -24970 85801 -24926
rect 85893 -24970 85901 -24926
rect 85993 -24970 86001 -24926
rect 86093 -24970 86101 -24926
rect 86193 -24970 86201 -24926
rect 86293 -24970 86301 -24926
rect 86393 -24970 86401 -24926
rect 86893 -24970 86901 -24926
rect 86993 -24970 87001 -24926
rect 87093 -24970 87101 -24926
rect 87193 -24970 87201 -24926
rect 87293 -24970 87301 -24926
rect 87393 -24970 87401 -24926
rect 87493 -24970 87501 -24926
rect 87593 -24970 87601 -24926
rect 87693 -24970 87701 -24926
rect 87793 -24970 87801 -24926
rect 87893 -24970 87901 -24926
rect 87993 -24970 88001 -24926
rect 88093 -24970 88101 -24926
rect 88193 -24970 88201 -24926
rect 88293 -24970 88301 -24926
rect 88393 -24970 88401 -24926
rect 109148 -24939 109156 -24895
rect 109248 -24939 109256 -24895
rect 109348 -24939 109356 -24895
rect 109448 -24939 109456 -24895
rect 109548 -24939 109556 -24895
rect 109648 -24939 109656 -24895
rect 109748 -24939 109756 -24895
rect 109848 -24939 109856 -24895
rect 109948 -24939 109956 -24895
rect 110048 -24939 110056 -24895
rect 110148 -24939 110156 -24895
rect 110248 -24939 110256 -24895
rect 110348 -24939 110356 -24895
rect 110448 -24939 110456 -24895
rect 110548 -24939 110556 -24895
rect 110648 -24939 110656 -24895
rect 111148 -24939 111156 -24895
rect 111248 -24939 111256 -24895
rect 111348 -24939 111356 -24895
rect 111448 -24939 111456 -24895
rect 111548 -24939 111556 -24895
rect 111648 -24939 111656 -24895
rect 111748 -24939 111756 -24895
rect 111848 -24939 111856 -24895
rect 111948 -24939 111956 -24895
rect 112048 -24939 112056 -24895
rect 112148 -24939 112156 -24895
rect 112248 -24939 112256 -24895
rect 112348 -24939 112356 -24895
rect 112448 -24939 112456 -24895
rect 112548 -24939 112556 -24895
rect 112648 -24939 112656 -24895
rect 113148 -24939 113156 -24895
rect 113248 -24939 113256 -24895
rect 113348 -24939 113356 -24895
rect 113448 -24939 113456 -24895
rect 113548 -24939 113556 -24895
rect 113648 -24939 113656 -24895
rect 113748 -24939 113756 -24895
rect 113848 -24939 113856 -24895
rect 113948 -24939 113956 -24895
rect 114048 -24939 114056 -24895
rect 114148 -24939 114156 -24895
rect 114248 -24939 114256 -24895
rect 114348 -24939 114356 -24895
rect 114448 -24939 114456 -24895
rect 114548 -24939 114556 -24895
rect 114648 -24939 114656 -24895
rect 115148 -24939 115156 -24895
rect 115248 -24939 115256 -24895
rect 115348 -24939 115356 -24895
rect 115448 -24939 115456 -24895
rect 115548 -24939 115556 -24895
rect 115648 -24939 115656 -24895
rect 115748 -24939 115756 -24895
rect 115848 -24939 115856 -24895
rect 115948 -24939 115956 -24895
rect 116048 -24939 116056 -24895
rect 116148 -24939 116156 -24895
rect 116248 -24939 116256 -24895
rect 116348 -24939 116356 -24895
rect 116448 -24939 116456 -24895
rect 116548 -24939 116556 -24895
rect 116648 -24939 116656 -24895
rect 109104 -24995 109148 -24987
rect 109204 -24995 109248 -24987
rect 109304 -24995 109348 -24987
rect 109404 -24995 109448 -24987
rect 109504 -24995 109548 -24987
rect 109604 -24995 109648 -24987
rect 109704 -24995 109748 -24987
rect 109804 -24995 109848 -24987
rect 109904 -24995 109948 -24987
rect 110004 -24995 110048 -24987
rect 110104 -24995 110148 -24987
rect 110204 -24995 110248 -24987
rect 110304 -24995 110348 -24987
rect 110404 -24995 110448 -24987
rect 110504 -24995 110548 -24987
rect 110604 -24995 110648 -24987
rect 111104 -24995 111148 -24987
rect 111204 -24995 111248 -24987
rect 111304 -24995 111348 -24987
rect 111404 -24995 111448 -24987
rect 111504 -24995 111548 -24987
rect 111604 -24995 111648 -24987
rect 111704 -24995 111748 -24987
rect 111804 -24995 111848 -24987
rect 111904 -24995 111948 -24987
rect 112004 -24995 112048 -24987
rect 112104 -24995 112148 -24987
rect 112204 -24995 112248 -24987
rect 112304 -24995 112348 -24987
rect 112404 -24995 112448 -24987
rect 112504 -24995 112548 -24987
rect 112604 -24995 112648 -24987
rect 113104 -24995 113148 -24987
rect 113204 -24995 113248 -24987
rect 113304 -24995 113348 -24987
rect 113404 -24995 113448 -24987
rect 113504 -24995 113548 -24987
rect 113604 -24995 113648 -24987
rect 113704 -24995 113748 -24987
rect 113804 -24995 113848 -24987
rect 113904 -24995 113948 -24987
rect 114004 -24995 114048 -24987
rect 114104 -24995 114148 -24987
rect 114204 -24995 114248 -24987
rect 114304 -24995 114348 -24987
rect 114404 -24995 114448 -24987
rect 114504 -24995 114548 -24987
rect 114604 -24995 114648 -24987
rect 115104 -24995 115148 -24987
rect 115204 -24995 115248 -24987
rect 115304 -24995 115348 -24987
rect 115404 -24995 115448 -24987
rect 115504 -24995 115548 -24987
rect 115604 -24995 115648 -24987
rect 115704 -24995 115748 -24987
rect 115804 -24995 115848 -24987
rect 115904 -24995 115948 -24987
rect 116004 -24995 116048 -24987
rect 116104 -24995 116148 -24987
rect 116204 -24995 116248 -24987
rect 116304 -24995 116348 -24987
rect 116404 -24995 116448 -24987
rect 116504 -24995 116548 -24987
rect 116604 -24995 116648 -24987
rect 80849 -25026 80893 -25018
rect 80949 -25026 80993 -25018
rect 81049 -25026 81093 -25018
rect 81149 -25026 81193 -25018
rect 81249 -25026 81293 -25018
rect 81349 -25026 81393 -25018
rect 81449 -25026 81493 -25018
rect 81549 -25026 81593 -25018
rect 81649 -25026 81693 -25018
rect 81749 -25026 81793 -25018
rect 81849 -25026 81893 -25018
rect 81949 -25026 81993 -25018
rect 82049 -25026 82093 -25018
rect 82149 -25026 82193 -25018
rect 82249 -25026 82293 -25018
rect 82349 -25026 82393 -25018
rect 82849 -25026 82893 -25018
rect 82949 -25026 82993 -25018
rect 83049 -25026 83093 -25018
rect 83149 -25026 83193 -25018
rect 83249 -25026 83293 -25018
rect 83349 -25026 83393 -25018
rect 83449 -25026 83493 -25018
rect 83549 -25026 83593 -25018
rect 83649 -25026 83693 -25018
rect 83749 -25026 83793 -25018
rect 83849 -25026 83893 -25018
rect 83949 -25026 83993 -25018
rect 84049 -25026 84093 -25018
rect 84149 -25026 84193 -25018
rect 84249 -25026 84293 -25018
rect 84349 -25026 84393 -25018
rect 84849 -25026 84893 -25018
rect 84949 -25026 84993 -25018
rect 85049 -25026 85093 -25018
rect 85149 -25026 85193 -25018
rect 85249 -25026 85293 -25018
rect 85349 -25026 85393 -25018
rect 85449 -25026 85493 -25018
rect 85549 -25026 85593 -25018
rect 85649 -25026 85693 -25018
rect 85749 -25026 85793 -25018
rect 85849 -25026 85893 -25018
rect 85949 -25026 85993 -25018
rect 86049 -25026 86093 -25018
rect 86149 -25026 86193 -25018
rect 86249 -25026 86293 -25018
rect 86349 -25026 86393 -25018
rect 86849 -25026 86893 -25018
rect 86949 -25026 86993 -25018
rect 87049 -25026 87093 -25018
rect 87149 -25026 87193 -25018
rect 87249 -25026 87293 -25018
rect 87349 -25026 87393 -25018
rect 87449 -25026 87493 -25018
rect 87549 -25026 87593 -25018
rect 87649 -25026 87693 -25018
rect 87749 -25026 87793 -25018
rect 87849 -25026 87893 -25018
rect 87949 -25026 87993 -25018
rect 88049 -25026 88093 -25018
rect 88149 -25026 88193 -25018
rect 88249 -25026 88293 -25018
rect 88349 -25026 88393 -25018
rect 80893 -25070 80901 -25026
rect 80993 -25070 81001 -25026
rect 81093 -25070 81101 -25026
rect 81193 -25070 81201 -25026
rect 81293 -25070 81301 -25026
rect 81393 -25070 81401 -25026
rect 81493 -25070 81501 -25026
rect 81593 -25070 81601 -25026
rect 81693 -25070 81701 -25026
rect 81793 -25070 81801 -25026
rect 81893 -25070 81901 -25026
rect 81993 -25070 82001 -25026
rect 82093 -25070 82101 -25026
rect 82193 -25070 82201 -25026
rect 82293 -25070 82301 -25026
rect 82393 -25070 82401 -25026
rect 82893 -25070 82901 -25026
rect 82993 -25070 83001 -25026
rect 83093 -25070 83101 -25026
rect 83193 -25070 83201 -25026
rect 83293 -25070 83301 -25026
rect 83393 -25070 83401 -25026
rect 83493 -25070 83501 -25026
rect 83593 -25070 83601 -25026
rect 83693 -25070 83701 -25026
rect 83793 -25070 83801 -25026
rect 83893 -25070 83901 -25026
rect 83993 -25070 84001 -25026
rect 84093 -25070 84101 -25026
rect 84193 -25070 84201 -25026
rect 84293 -25070 84301 -25026
rect 84393 -25070 84401 -25026
rect 84893 -25070 84901 -25026
rect 84993 -25070 85001 -25026
rect 85093 -25070 85101 -25026
rect 85193 -25070 85201 -25026
rect 85293 -25070 85301 -25026
rect 85393 -25070 85401 -25026
rect 85493 -25070 85501 -25026
rect 85593 -25070 85601 -25026
rect 85693 -25070 85701 -25026
rect 85793 -25070 85801 -25026
rect 85893 -25070 85901 -25026
rect 85993 -25070 86001 -25026
rect 86093 -25070 86101 -25026
rect 86193 -25070 86201 -25026
rect 86293 -25070 86301 -25026
rect 86393 -25070 86401 -25026
rect 86893 -25070 86901 -25026
rect 86993 -25070 87001 -25026
rect 87093 -25070 87101 -25026
rect 87193 -25070 87201 -25026
rect 87293 -25070 87301 -25026
rect 87393 -25070 87401 -25026
rect 87493 -25070 87501 -25026
rect 87593 -25070 87601 -25026
rect 87693 -25070 87701 -25026
rect 87793 -25070 87801 -25026
rect 87893 -25070 87901 -25026
rect 87993 -25070 88001 -25026
rect 88093 -25070 88101 -25026
rect 88193 -25070 88201 -25026
rect 88293 -25070 88301 -25026
rect 88393 -25070 88401 -25026
rect 109148 -25039 109156 -24995
rect 109248 -25039 109256 -24995
rect 109348 -25039 109356 -24995
rect 109448 -25039 109456 -24995
rect 109548 -25039 109556 -24995
rect 109648 -25039 109656 -24995
rect 109748 -25039 109756 -24995
rect 109848 -25039 109856 -24995
rect 109948 -25039 109956 -24995
rect 110048 -25039 110056 -24995
rect 110148 -25039 110156 -24995
rect 110248 -25039 110256 -24995
rect 110348 -25039 110356 -24995
rect 110448 -25039 110456 -24995
rect 110548 -25039 110556 -24995
rect 110648 -25039 110656 -24995
rect 111148 -25039 111156 -24995
rect 111248 -25039 111256 -24995
rect 111348 -25039 111356 -24995
rect 111448 -25039 111456 -24995
rect 111548 -25039 111556 -24995
rect 111648 -25039 111656 -24995
rect 111748 -25039 111756 -24995
rect 111848 -25039 111856 -24995
rect 111948 -25039 111956 -24995
rect 112048 -25039 112056 -24995
rect 112148 -25039 112156 -24995
rect 112248 -25039 112256 -24995
rect 112348 -25039 112356 -24995
rect 112448 -25039 112456 -24995
rect 112548 -25039 112556 -24995
rect 112648 -25039 112656 -24995
rect 113148 -25039 113156 -24995
rect 113248 -25039 113256 -24995
rect 113348 -25039 113356 -24995
rect 113448 -25039 113456 -24995
rect 113548 -25039 113556 -24995
rect 113648 -25039 113656 -24995
rect 113748 -25039 113756 -24995
rect 113848 -25039 113856 -24995
rect 113948 -25039 113956 -24995
rect 114048 -25039 114056 -24995
rect 114148 -25039 114156 -24995
rect 114248 -25039 114256 -24995
rect 114348 -25039 114356 -24995
rect 114448 -25039 114456 -24995
rect 114548 -25039 114556 -24995
rect 114648 -25039 114656 -24995
rect 115148 -25039 115156 -24995
rect 115248 -25039 115256 -24995
rect 115348 -25039 115356 -24995
rect 115448 -25039 115456 -24995
rect 115548 -25039 115556 -24995
rect 115648 -25039 115656 -24995
rect 115748 -25039 115756 -24995
rect 115848 -25039 115856 -24995
rect 115948 -25039 115956 -24995
rect 116048 -25039 116056 -24995
rect 116148 -25039 116156 -24995
rect 116248 -25039 116256 -24995
rect 116348 -25039 116356 -24995
rect 116448 -25039 116456 -24995
rect 116548 -25039 116556 -24995
rect 116648 -25039 116656 -24995
rect 109104 -25095 109148 -25087
rect 109204 -25095 109248 -25087
rect 109304 -25095 109348 -25087
rect 109404 -25095 109448 -25087
rect 109504 -25095 109548 -25087
rect 109604 -25095 109648 -25087
rect 109704 -25095 109748 -25087
rect 109804 -25095 109848 -25087
rect 109904 -25095 109948 -25087
rect 110004 -25095 110048 -25087
rect 110104 -25095 110148 -25087
rect 110204 -25095 110248 -25087
rect 110304 -25095 110348 -25087
rect 110404 -25095 110448 -25087
rect 110504 -25095 110548 -25087
rect 110604 -25095 110648 -25087
rect 111104 -25095 111148 -25087
rect 111204 -25095 111248 -25087
rect 111304 -25095 111348 -25087
rect 111404 -25095 111448 -25087
rect 111504 -25095 111548 -25087
rect 111604 -25095 111648 -25087
rect 111704 -25095 111748 -25087
rect 111804 -25095 111848 -25087
rect 111904 -25095 111948 -25087
rect 112004 -25095 112048 -25087
rect 112104 -25095 112148 -25087
rect 112204 -25095 112248 -25087
rect 112304 -25095 112348 -25087
rect 112404 -25095 112448 -25087
rect 112504 -25095 112548 -25087
rect 112604 -25095 112648 -25087
rect 113104 -25095 113148 -25087
rect 113204 -25095 113248 -25087
rect 113304 -25095 113348 -25087
rect 113404 -25095 113448 -25087
rect 113504 -25095 113548 -25087
rect 113604 -25095 113648 -25087
rect 113704 -25095 113748 -25087
rect 113804 -25095 113848 -25087
rect 113904 -25095 113948 -25087
rect 114004 -25095 114048 -25087
rect 114104 -25095 114148 -25087
rect 114204 -25095 114248 -25087
rect 114304 -25095 114348 -25087
rect 114404 -25095 114448 -25087
rect 114504 -25095 114548 -25087
rect 114604 -25095 114648 -25087
rect 115104 -25095 115148 -25087
rect 115204 -25095 115248 -25087
rect 115304 -25095 115348 -25087
rect 115404 -25095 115448 -25087
rect 115504 -25095 115548 -25087
rect 115604 -25095 115648 -25087
rect 115704 -25095 115748 -25087
rect 115804 -25095 115848 -25087
rect 115904 -25095 115948 -25087
rect 116004 -25095 116048 -25087
rect 116104 -25095 116148 -25087
rect 116204 -25095 116248 -25087
rect 116304 -25095 116348 -25087
rect 116404 -25095 116448 -25087
rect 116504 -25095 116548 -25087
rect 116604 -25095 116648 -25087
rect 80849 -25126 80893 -25118
rect 80949 -25126 80993 -25118
rect 81049 -25126 81093 -25118
rect 81149 -25126 81193 -25118
rect 81249 -25126 81293 -25118
rect 81349 -25126 81393 -25118
rect 81449 -25126 81493 -25118
rect 81549 -25126 81593 -25118
rect 81649 -25126 81693 -25118
rect 81749 -25126 81793 -25118
rect 81849 -25126 81893 -25118
rect 81949 -25126 81993 -25118
rect 82049 -25126 82093 -25118
rect 82149 -25126 82193 -25118
rect 82249 -25126 82293 -25118
rect 82349 -25126 82393 -25118
rect 82849 -25126 82893 -25118
rect 82949 -25126 82993 -25118
rect 83049 -25126 83093 -25118
rect 83149 -25126 83193 -25118
rect 83249 -25126 83293 -25118
rect 83349 -25126 83393 -25118
rect 83449 -25126 83493 -25118
rect 83549 -25126 83593 -25118
rect 83649 -25126 83693 -25118
rect 83749 -25126 83793 -25118
rect 83849 -25126 83893 -25118
rect 83949 -25126 83993 -25118
rect 84049 -25126 84093 -25118
rect 84149 -25126 84193 -25118
rect 84249 -25126 84293 -25118
rect 84349 -25126 84393 -25118
rect 84849 -25126 84893 -25118
rect 84949 -25126 84993 -25118
rect 85049 -25126 85093 -25118
rect 85149 -25126 85193 -25118
rect 85249 -25126 85293 -25118
rect 85349 -25126 85393 -25118
rect 85449 -25126 85493 -25118
rect 85549 -25126 85593 -25118
rect 85649 -25126 85693 -25118
rect 85749 -25126 85793 -25118
rect 85849 -25126 85893 -25118
rect 85949 -25126 85993 -25118
rect 86049 -25126 86093 -25118
rect 86149 -25126 86193 -25118
rect 86249 -25126 86293 -25118
rect 86349 -25126 86393 -25118
rect 86849 -25126 86893 -25118
rect 86949 -25126 86993 -25118
rect 87049 -25126 87093 -25118
rect 87149 -25126 87193 -25118
rect 87249 -25126 87293 -25118
rect 87349 -25126 87393 -25118
rect 87449 -25126 87493 -25118
rect 87549 -25126 87593 -25118
rect 87649 -25126 87693 -25118
rect 87749 -25126 87793 -25118
rect 87849 -25126 87893 -25118
rect 87949 -25126 87993 -25118
rect 88049 -25126 88093 -25118
rect 88149 -25126 88193 -25118
rect 88249 -25126 88293 -25118
rect 88349 -25126 88393 -25118
rect 80893 -25170 80901 -25126
rect 80993 -25170 81001 -25126
rect 81093 -25170 81101 -25126
rect 81193 -25170 81201 -25126
rect 81293 -25170 81301 -25126
rect 81393 -25170 81401 -25126
rect 81493 -25170 81501 -25126
rect 81593 -25170 81601 -25126
rect 81693 -25170 81701 -25126
rect 81793 -25170 81801 -25126
rect 81893 -25170 81901 -25126
rect 81993 -25170 82001 -25126
rect 82093 -25170 82101 -25126
rect 82193 -25170 82201 -25126
rect 82293 -25170 82301 -25126
rect 82393 -25170 82401 -25126
rect 82893 -25170 82901 -25126
rect 82993 -25170 83001 -25126
rect 83093 -25170 83101 -25126
rect 83193 -25170 83201 -25126
rect 83293 -25170 83301 -25126
rect 83393 -25170 83401 -25126
rect 83493 -25170 83501 -25126
rect 83593 -25170 83601 -25126
rect 83693 -25170 83701 -25126
rect 83793 -25170 83801 -25126
rect 83893 -25170 83901 -25126
rect 83993 -25170 84001 -25126
rect 84093 -25170 84101 -25126
rect 84193 -25170 84201 -25126
rect 84293 -25170 84301 -25126
rect 84393 -25170 84401 -25126
rect 84893 -25170 84901 -25126
rect 84993 -25170 85001 -25126
rect 85093 -25170 85101 -25126
rect 85193 -25170 85201 -25126
rect 85293 -25170 85301 -25126
rect 85393 -25170 85401 -25126
rect 85493 -25170 85501 -25126
rect 85593 -25170 85601 -25126
rect 85693 -25170 85701 -25126
rect 85793 -25170 85801 -25126
rect 85893 -25170 85901 -25126
rect 85993 -25170 86001 -25126
rect 86093 -25170 86101 -25126
rect 86193 -25170 86201 -25126
rect 86293 -25170 86301 -25126
rect 86393 -25170 86401 -25126
rect 86893 -25170 86901 -25126
rect 86993 -25170 87001 -25126
rect 87093 -25170 87101 -25126
rect 87193 -25170 87201 -25126
rect 87293 -25170 87301 -25126
rect 87393 -25170 87401 -25126
rect 87493 -25170 87501 -25126
rect 87593 -25170 87601 -25126
rect 87693 -25170 87701 -25126
rect 87793 -25170 87801 -25126
rect 87893 -25170 87901 -25126
rect 87993 -25170 88001 -25126
rect 88093 -25170 88101 -25126
rect 88193 -25170 88201 -25126
rect 88293 -25170 88301 -25126
rect 88393 -25170 88401 -25126
rect 109148 -25139 109156 -25095
rect 109248 -25139 109256 -25095
rect 109348 -25139 109356 -25095
rect 109448 -25139 109456 -25095
rect 109548 -25139 109556 -25095
rect 109648 -25139 109656 -25095
rect 109748 -25139 109756 -25095
rect 109848 -25139 109856 -25095
rect 109948 -25139 109956 -25095
rect 110048 -25139 110056 -25095
rect 110148 -25139 110156 -25095
rect 110248 -25139 110256 -25095
rect 110348 -25139 110356 -25095
rect 110448 -25139 110456 -25095
rect 110548 -25139 110556 -25095
rect 110648 -25139 110656 -25095
rect 111148 -25139 111156 -25095
rect 111248 -25139 111256 -25095
rect 111348 -25139 111356 -25095
rect 111448 -25139 111456 -25095
rect 111548 -25139 111556 -25095
rect 111648 -25139 111656 -25095
rect 111748 -25139 111756 -25095
rect 111848 -25139 111856 -25095
rect 111948 -25139 111956 -25095
rect 112048 -25139 112056 -25095
rect 112148 -25139 112156 -25095
rect 112248 -25139 112256 -25095
rect 112348 -25139 112356 -25095
rect 112448 -25139 112456 -25095
rect 112548 -25139 112556 -25095
rect 112648 -25139 112656 -25095
rect 113148 -25139 113156 -25095
rect 113248 -25139 113256 -25095
rect 113348 -25139 113356 -25095
rect 113448 -25139 113456 -25095
rect 113548 -25139 113556 -25095
rect 113648 -25139 113656 -25095
rect 113748 -25139 113756 -25095
rect 113848 -25139 113856 -25095
rect 113948 -25139 113956 -25095
rect 114048 -25139 114056 -25095
rect 114148 -25139 114156 -25095
rect 114248 -25139 114256 -25095
rect 114348 -25139 114356 -25095
rect 114448 -25139 114456 -25095
rect 114548 -25139 114556 -25095
rect 114648 -25139 114656 -25095
rect 115148 -25139 115156 -25095
rect 115248 -25139 115256 -25095
rect 115348 -25139 115356 -25095
rect 115448 -25139 115456 -25095
rect 115548 -25139 115556 -25095
rect 115648 -25139 115656 -25095
rect 115748 -25139 115756 -25095
rect 115848 -25139 115856 -25095
rect 115948 -25139 115956 -25095
rect 116048 -25139 116056 -25095
rect 116148 -25139 116156 -25095
rect 116248 -25139 116256 -25095
rect 116348 -25139 116356 -25095
rect 116448 -25139 116456 -25095
rect 116548 -25139 116556 -25095
rect 116648 -25139 116656 -25095
rect 109104 -25195 109148 -25187
rect 109204 -25195 109248 -25187
rect 109304 -25195 109348 -25187
rect 109404 -25195 109448 -25187
rect 109504 -25195 109548 -25187
rect 109604 -25195 109648 -25187
rect 109704 -25195 109748 -25187
rect 109804 -25195 109848 -25187
rect 109904 -25195 109948 -25187
rect 110004 -25195 110048 -25187
rect 110104 -25195 110148 -25187
rect 110204 -25195 110248 -25187
rect 110304 -25195 110348 -25187
rect 110404 -25195 110448 -25187
rect 110504 -25195 110548 -25187
rect 110604 -25195 110648 -25187
rect 111104 -25195 111148 -25187
rect 111204 -25195 111248 -25187
rect 111304 -25195 111348 -25187
rect 111404 -25195 111448 -25187
rect 111504 -25195 111548 -25187
rect 111604 -25195 111648 -25187
rect 111704 -25195 111748 -25187
rect 111804 -25195 111848 -25187
rect 111904 -25195 111948 -25187
rect 112004 -25195 112048 -25187
rect 112104 -25195 112148 -25187
rect 112204 -25195 112248 -25187
rect 112304 -25195 112348 -25187
rect 112404 -25195 112448 -25187
rect 112504 -25195 112548 -25187
rect 112604 -25195 112648 -25187
rect 113104 -25195 113148 -25187
rect 113204 -25195 113248 -25187
rect 113304 -25195 113348 -25187
rect 113404 -25195 113448 -25187
rect 113504 -25195 113548 -25187
rect 113604 -25195 113648 -25187
rect 113704 -25195 113748 -25187
rect 113804 -25195 113848 -25187
rect 113904 -25195 113948 -25187
rect 114004 -25195 114048 -25187
rect 114104 -25195 114148 -25187
rect 114204 -25195 114248 -25187
rect 114304 -25195 114348 -25187
rect 114404 -25195 114448 -25187
rect 114504 -25195 114548 -25187
rect 114604 -25195 114648 -25187
rect 115104 -25195 115148 -25187
rect 115204 -25195 115248 -25187
rect 115304 -25195 115348 -25187
rect 115404 -25195 115448 -25187
rect 115504 -25195 115548 -25187
rect 115604 -25195 115648 -25187
rect 115704 -25195 115748 -25187
rect 115804 -25195 115848 -25187
rect 115904 -25195 115948 -25187
rect 116004 -25195 116048 -25187
rect 116104 -25195 116148 -25187
rect 116204 -25195 116248 -25187
rect 116304 -25195 116348 -25187
rect 116404 -25195 116448 -25187
rect 116504 -25195 116548 -25187
rect 116604 -25195 116648 -25187
rect 80849 -25226 80893 -25218
rect 80949 -25226 80993 -25218
rect 81049 -25226 81093 -25218
rect 81149 -25226 81193 -25218
rect 81249 -25226 81293 -25218
rect 81349 -25226 81393 -25218
rect 81449 -25226 81493 -25218
rect 81549 -25226 81593 -25218
rect 81649 -25226 81693 -25218
rect 81749 -25226 81793 -25218
rect 81849 -25226 81893 -25218
rect 81949 -25226 81993 -25218
rect 82049 -25226 82093 -25218
rect 82149 -25226 82193 -25218
rect 82249 -25226 82293 -25218
rect 82349 -25226 82393 -25218
rect 82849 -25226 82893 -25218
rect 82949 -25226 82993 -25218
rect 83049 -25226 83093 -25218
rect 83149 -25226 83193 -25218
rect 83249 -25226 83293 -25218
rect 83349 -25226 83393 -25218
rect 83449 -25226 83493 -25218
rect 83549 -25226 83593 -25218
rect 83649 -25226 83693 -25218
rect 83749 -25226 83793 -25218
rect 83849 -25226 83893 -25218
rect 83949 -25226 83993 -25218
rect 84049 -25226 84093 -25218
rect 84149 -25226 84193 -25218
rect 84249 -25226 84293 -25218
rect 84349 -25226 84393 -25218
rect 84849 -25226 84893 -25218
rect 84949 -25226 84993 -25218
rect 85049 -25226 85093 -25218
rect 85149 -25226 85193 -25218
rect 85249 -25226 85293 -25218
rect 85349 -25226 85393 -25218
rect 85449 -25226 85493 -25218
rect 85549 -25226 85593 -25218
rect 85649 -25226 85693 -25218
rect 85749 -25226 85793 -25218
rect 85849 -25226 85893 -25218
rect 85949 -25226 85993 -25218
rect 86049 -25226 86093 -25218
rect 86149 -25226 86193 -25218
rect 86249 -25226 86293 -25218
rect 86349 -25226 86393 -25218
rect 86849 -25226 86893 -25218
rect 86949 -25226 86993 -25218
rect 87049 -25226 87093 -25218
rect 87149 -25226 87193 -25218
rect 87249 -25226 87293 -25218
rect 87349 -25226 87393 -25218
rect 87449 -25226 87493 -25218
rect 87549 -25226 87593 -25218
rect 87649 -25226 87693 -25218
rect 87749 -25226 87793 -25218
rect 87849 -25226 87893 -25218
rect 87949 -25226 87993 -25218
rect 88049 -25226 88093 -25218
rect 88149 -25226 88193 -25218
rect 88249 -25226 88293 -25218
rect 88349 -25226 88393 -25218
rect 80893 -25270 80901 -25226
rect 80993 -25270 81001 -25226
rect 81093 -25270 81101 -25226
rect 81193 -25270 81201 -25226
rect 81293 -25270 81301 -25226
rect 81393 -25270 81401 -25226
rect 81493 -25270 81501 -25226
rect 81593 -25270 81601 -25226
rect 81693 -25270 81701 -25226
rect 81793 -25270 81801 -25226
rect 81893 -25270 81901 -25226
rect 81993 -25270 82001 -25226
rect 82093 -25270 82101 -25226
rect 82193 -25270 82201 -25226
rect 82293 -25270 82301 -25226
rect 82393 -25270 82401 -25226
rect 82893 -25270 82901 -25226
rect 82993 -25270 83001 -25226
rect 83093 -25270 83101 -25226
rect 83193 -25270 83201 -25226
rect 83293 -25270 83301 -25226
rect 83393 -25270 83401 -25226
rect 83493 -25270 83501 -25226
rect 83593 -25270 83601 -25226
rect 83693 -25270 83701 -25226
rect 83793 -25270 83801 -25226
rect 83893 -25270 83901 -25226
rect 83993 -25270 84001 -25226
rect 84093 -25270 84101 -25226
rect 84193 -25270 84201 -25226
rect 84293 -25270 84301 -25226
rect 84393 -25270 84401 -25226
rect 84893 -25270 84901 -25226
rect 84993 -25270 85001 -25226
rect 85093 -25270 85101 -25226
rect 85193 -25270 85201 -25226
rect 85293 -25270 85301 -25226
rect 85393 -25270 85401 -25226
rect 85493 -25270 85501 -25226
rect 85593 -25270 85601 -25226
rect 85693 -25270 85701 -25226
rect 85793 -25270 85801 -25226
rect 85893 -25270 85901 -25226
rect 85993 -25270 86001 -25226
rect 86093 -25270 86101 -25226
rect 86193 -25270 86201 -25226
rect 86293 -25270 86301 -25226
rect 86393 -25270 86401 -25226
rect 86893 -25270 86901 -25226
rect 86993 -25270 87001 -25226
rect 87093 -25270 87101 -25226
rect 87193 -25270 87201 -25226
rect 87293 -25270 87301 -25226
rect 87393 -25270 87401 -25226
rect 87493 -25270 87501 -25226
rect 87593 -25270 87601 -25226
rect 87693 -25270 87701 -25226
rect 87793 -25270 87801 -25226
rect 87893 -25270 87901 -25226
rect 87993 -25270 88001 -25226
rect 88093 -25270 88101 -25226
rect 88193 -25270 88201 -25226
rect 88293 -25270 88301 -25226
rect 88393 -25270 88401 -25226
rect 109148 -25239 109156 -25195
rect 109248 -25239 109256 -25195
rect 109348 -25239 109356 -25195
rect 109448 -25239 109456 -25195
rect 109548 -25239 109556 -25195
rect 109648 -25239 109656 -25195
rect 109748 -25239 109756 -25195
rect 109848 -25239 109856 -25195
rect 109948 -25239 109956 -25195
rect 110048 -25239 110056 -25195
rect 110148 -25239 110156 -25195
rect 110248 -25239 110256 -25195
rect 110348 -25239 110356 -25195
rect 110448 -25239 110456 -25195
rect 110548 -25239 110556 -25195
rect 110648 -25239 110656 -25195
rect 111148 -25239 111156 -25195
rect 111248 -25239 111256 -25195
rect 111348 -25239 111356 -25195
rect 111448 -25239 111456 -25195
rect 111548 -25239 111556 -25195
rect 111648 -25239 111656 -25195
rect 111748 -25239 111756 -25195
rect 111848 -25239 111856 -25195
rect 111948 -25239 111956 -25195
rect 112048 -25239 112056 -25195
rect 112148 -25239 112156 -25195
rect 112248 -25239 112256 -25195
rect 112348 -25239 112356 -25195
rect 112448 -25239 112456 -25195
rect 112548 -25239 112556 -25195
rect 112648 -25239 112656 -25195
rect 113148 -25239 113156 -25195
rect 113248 -25239 113256 -25195
rect 113348 -25239 113356 -25195
rect 113448 -25239 113456 -25195
rect 113548 -25239 113556 -25195
rect 113648 -25239 113656 -25195
rect 113748 -25239 113756 -25195
rect 113848 -25239 113856 -25195
rect 113948 -25239 113956 -25195
rect 114048 -25239 114056 -25195
rect 114148 -25239 114156 -25195
rect 114248 -25239 114256 -25195
rect 114348 -25239 114356 -25195
rect 114448 -25239 114456 -25195
rect 114548 -25239 114556 -25195
rect 114648 -25239 114656 -25195
rect 115148 -25239 115156 -25195
rect 115248 -25239 115256 -25195
rect 115348 -25239 115356 -25195
rect 115448 -25239 115456 -25195
rect 115548 -25239 115556 -25195
rect 115648 -25239 115656 -25195
rect 115748 -25239 115756 -25195
rect 115848 -25239 115856 -25195
rect 115948 -25239 115956 -25195
rect 116048 -25239 116056 -25195
rect 116148 -25239 116156 -25195
rect 116248 -25239 116256 -25195
rect 116348 -25239 116356 -25195
rect 116448 -25239 116456 -25195
rect 116548 -25239 116556 -25195
rect 116648 -25239 116656 -25195
rect 109104 -25295 109148 -25287
rect 109204 -25295 109248 -25287
rect 109304 -25295 109348 -25287
rect 109404 -25295 109448 -25287
rect 109504 -25295 109548 -25287
rect 109604 -25295 109648 -25287
rect 109704 -25295 109748 -25287
rect 109804 -25295 109848 -25287
rect 109904 -25295 109948 -25287
rect 110004 -25295 110048 -25287
rect 110104 -25295 110148 -25287
rect 110204 -25295 110248 -25287
rect 110304 -25295 110348 -25287
rect 110404 -25295 110448 -25287
rect 110504 -25295 110548 -25287
rect 110604 -25295 110648 -25287
rect 111104 -25295 111148 -25287
rect 111204 -25295 111248 -25287
rect 111304 -25295 111348 -25287
rect 111404 -25295 111448 -25287
rect 111504 -25295 111548 -25287
rect 111604 -25295 111648 -25287
rect 111704 -25295 111748 -25287
rect 111804 -25295 111848 -25287
rect 111904 -25295 111948 -25287
rect 112004 -25295 112048 -25287
rect 112104 -25295 112148 -25287
rect 112204 -25295 112248 -25287
rect 112304 -25295 112348 -25287
rect 112404 -25295 112448 -25287
rect 112504 -25295 112548 -25287
rect 112604 -25295 112648 -25287
rect 113104 -25295 113148 -25287
rect 113204 -25295 113248 -25287
rect 113304 -25295 113348 -25287
rect 113404 -25295 113448 -25287
rect 113504 -25295 113548 -25287
rect 113604 -25295 113648 -25287
rect 113704 -25295 113748 -25287
rect 113804 -25295 113848 -25287
rect 113904 -25295 113948 -25287
rect 114004 -25295 114048 -25287
rect 114104 -25295 114148 -25287
rect 114204 -25295 114248 -25287
rect 114304 -25295 114348 -25287
rect 114404 -25295 114448 -25287
rect 114504 -25295 114548 -25287
rect 114604 -25295 114648 -25287
rect 115104 -25295 115148 -25287
rect 115204 -25295 115248 -25287
rect 115304 -25295 115348 -25287
rect 115404 -25295 115448 -25287
rect 115504 -25295 115548 -25287
rect 115604 -25295 115648 -25287
rect 115704 -25295 115748 -25287
rect 115804 -25295 115848 -25287
rect 115904 -25295 115948 -25287
rect 116004 -25295 116048 -25287
rect 116104 -25295 116148 -25287
rect 116204 -25295 116248 -25287
rect 116304 -25295 116348 -25287
rect 116404 -25295 116448 -25287
rect 116504 -25295 116548 -25287
rect 116604 -25295 116648 -25287
rect 80849 -25326 80893 -25318
rect 80949 -25326 80993 -25318
rect 81049 -25326 81093 -25318
rect 81149 -25326 81193 -25318
rect 81249 -25326 81293 -25318
rect 81349 -25326 81393 -25318
rect 81449 -25326 81493 -25318
rect 81549 -25326 81593 -25318
rect 81649 -25326 81693 -25318
rect 81749 -25326 81793 -25318
rect 81849 -25326 81893 -25318
rect 81949 -25326 81993 -25318
rect 82049 -25326 82093 -25318
rect 82149 -25326 82193 -25318
rect 82249 -25326 82293 -25318
rect 82349 -25326 82393 -25318
rect 82849 -25326 82893 -25318
rect 82949 -25326 82993 -25318
rect 83049 -25326 83093 -25318
rect 83149 -25326 83193 -25318
rect 83249 -25326 83293 -25318
rect 83349 -25326 83393 -25318
rect 83449 -25326 83493 -25318
rect 83549 -25326 83593 -25318
rect 83649 -25326 83693 -25318
rect 83749 -25326 83793 -25318
rect 83849 -25326 83893 -25318
rect 83949 -25326 83993 -25318
rect 84049 -25326 84093 -25318
rect 84149 -25326 84193 -25318
rect 84249 -25326 84293 -25318
rect 84349 -25326 84393 -25318
rect 84849 -25326 84893 -25318
rect 84949 -25326 84993 -25318
rect 85049 -25326 85093 -25318
rect 85149 -25326 85193 -25318
rect 85249 -25326 85293 -25318
rect 85349 -25326 85393 -25318
rect 85449 -25326 85493 -25318
rect 85549 -25326 85593 -25318
rect 85649 -25326 85693 -25318
rect 85749 -25326 85793 -25318
rect 85849 -25326 85893 -25318
rect 85949 -25326 85993 -25318
rect 86049 -25326 86093 -25318
rect 86149 -25326 86193 -25318
rect 86249 -25326 86293 -25318
rect 86349 -25326 86393 -25318
rect 86849 -25326 86893 -25318
rect 86949 -25326 86993 -25318
rect 87049 -25326 87093 -25318
rect 87149 -25326 87193 -25318
rect 87249 -25326 87293 -25318
rect 87349 -25326 87393 -25318
rect 87449 -25326 87493 -25318
rect 87549 -25326 87593 -25318
rect 87649 -25326 87693 -25318
rect 87749 -25326 87793 -25318
rect 87849 -25326 87893 -25318
rect 87949 -25326 87993 -25318
rect 88049 -25326 88093 -25318
rect 88149 -25326 88193 -25318
rect 88249 -25326 88293 -25318
rect 88349 -25326 88393 -25318
rect 80893 -25370 80901 -25326
rect 80993 -25370 81001 -25326
rect 81093 -25370 81101 -25326
rect 81193 -25370 81201 -25326
rect 81293 -25370 81301 -25326
rect 81393 -25370 81401 -25326
rect 81493 -25370 81501 -25326
rect 81593 -25370 81601 -25326
rect 81693 -25370 81701 -25326
rect 81793 -25370 81801 -25326
rect 81893 -25370 81901 -25326
rect 81993 -25370 82001 -25326
rect 82093 -25370 82101 -25326
rect 82193 -25370 82201 -25326
rect 82293 -25370 82301 -25326
rect 82393 -25370 82401 -25326
rect 82893 -25370 82901 -25326
rect 82993 -25370 83001 -25326
rect 83093 -25370 83101 -25326
rect 83193 -25370 83201 -25326
rect 83293 -25370 83301 -25326
rect 83393 -25370 83401 -25326
rect 83493 -25370 83501 -25326
rect 83593 -25370 83601 -25326
rect 83693 -25370 83701 -25326
rect 83793 -25370 83801 -25326
rect 83893 -25370 83901 -25326
rect 83993 -25370 84001 -25326
rect 84093 -25370 84101 -25326
rect 84193 -25370 84201 -25326
rect 84293 -25370 84301 -25326
rect 84393 -25370 84401 -25326
rect 84893 -25370 84901 -25326
rect 84993 -25370 85001 -25326
rect 85093 -25370 85101 -25326
rect 85193 -25370 85201 -25326
rect 85293 -25370 85301 -25326
rect 85393 -25370 85401 -25326
rect 85493 -25370 85501 -25326
rect 85593 -25370 85601 -25326
rect 85693 -25370 85701 -25326
rect 85793 -25370 85801 -25326
rect 85893 -25370 85901 -25326
rect 85993 -25370 86001 -25326
rect 86093 -25370 86101 -25326
rect 86193 -25370 86201 -25326
rect 86293 -25370 86301 -25326
rect 86393 -25370 86401 -25326
rect 86893 -25370 86901 -25326
rect 86993 -25370 87001 -25326
rect 87093 -25370 87101 -25326
rect 87193 -25370 87201 -25326
rect 87293 -25370 87301 -25326
rect 87393 -25370 87401 -25326
rect 87493 -25370 87501 -25326
rect 87593 -25370 87601 -25326
rect 87693 -25370 87701 -25326
rect 87793 -25370 87801 -25326
rect 87893 -25370 87901 -25326
rect 87993 -25370 88001 -25326
rect 88093 -25370 88101 -25326
rect 88193 -25370 88201 -25326
rect 88293 -25370 88301 -25326
rect 88393 -25370 88401 -25326
rect 109148 -25339 109156 -25295
rect 109248 -25339 109256 -25295
rect 109348 -25339 109356 -25295
rect 109448 -25339 109456 -25295
rect 109548 -25339 109556 -25295
rect 109648 -25339 109656 -25295
rect 109748 -25339 109756 -25295
rect 109848 -25339 109856 -25295
rect 109948 -25339 109956 -25295
rect 110048 -25339 110056 -25295
rect 110148 -25339 110156 -25295
rect 110248 -25339 110256 -25295
rect 110348 -25339 110356 -25295
rect 110448 -25339 110456 -25295
rect 110548 -25339 110556 -25295
rect 110648 -25339 110656 -25295
rect 111148 -25339 111156 -25295
rect 111248 -25339 111256 -25295
rect 111348 -25339 111356 -25295
rect 111448 -25339 111456 -25295
rect 111548 -25339 111556 -25295
rect 111648 -25339 111656 -25295
rect 111748 -25339 111756 -25295
rect 111848 -25339 111856 -25295
rect 111948 -25339 111956 -25295
rect 112048 -25339 112056 -25295
rect 112148 -25339 112156 -25295
rect 112248 -25339 112256 -25295
rect 112348 -25339 112356 -25295
rect 112448 -25339 112456 -25295
rect 112548 -25339 112556 -25295
rect 112648 -25339 112656 -25295
rect 113148 -25339 113156 -25295
rect 113248 -25339 113256 -25295
rect 113348 -25339 113356 -25295
rect 113448 -25339 113456 -25295
rect 113548 -25339 113556 -25295
rect 113648 -25339 113656 -25295
rect 113748 -25339 113756 -25295
rect 113848 -25339 113856 -25295
rect 113948 -25339 113956 -25295
rect 114048 -25339 114056 -25295
rect 114148 -25339 114156 -25295
rect 114248 -25339 114256 -25295
rect 114348 -25339 114356 -25295
rect 114448 -25339 114456 -25295
rect 114548 -25339 114556 -25295
rect 114648 -25339 114656 -25295
rect 115148 -25339 115156 -25295
rect 115248 -25339 115256 -25295
rect 115348 -25339 115356 -25295
rect 115448 -25339 115456 -25295
rect 115548 -25339 115556 -25295
rect 115648 -25339 115656 -25295
rect 115748 -25339 115756 -25295
rect 115848 -25339 115856 -25295
rect 115948 -25339 115956 -25295
rect 116048 -25339 116056 -25295
rect 116148 -25339 116156 -25295
rect 116248 -25339 116256 -25295
rect 116348 -25339 116356 -25295
rect 116448 -25339 116456 -25295
rect 116548 -25339 116556 -25295
rect 116648 -25339 116656 -25295
rect 109104 -25395 109148 -25387
rect 109204 -25395 109248 -25387
rect 109304 -25395 109348 -25387
rect 109404 -25395 109448 -25387
rect 109504 -25395 109548 -25387
rect 109604 -25395 109648 -25387
rect 109704 -25395 109748 -25387
rect 109804 -25395 109848 -25387
rect 109904 -25395 109948 -25387
rect 110004 -25395 110048 -25387
rect 110104 -25395 110148 -25387
rect 110204 -25395 110248 -25387
rect 110304 -25395 110348 -25387
rect 110404 -25395 110448 -25387
rect 110504 -25395 110548 -25387
rect 110604 -25395 110648 -25387
rect 111104 -25395 111148 -25387
rect 111204 -25395 111248 -25387
rect 111304 -25395 111348 -25387
rect 111404 -25395 111448 -25387
rect 111504 -25395 111548 -25387
rect 111604 -25395 111648 -25387
rect 111704 -25395 111748 -25387
rect 111804 -25395 111848 -25387
rect 111904 -25395 111948 -25387
rect 112004 -25395 112048 -25387
rect 112104 -25395 112148 -25387
rect 112204 -25395 112248 -25387
rect 112304 -25395 112348 -25387
rect 112404 -25395 112448 -25387
rect 112504 -25395 112548 -25387
rect 112604 -25395 112648 -25387
rect 113104 -25395 113148 -25387
rect 113204 -25395 113248 -25387
rect 113304 -25395 113348 -25387
rect 113404 -25395 113448 -25387
rect 113504 -25395 113548 -25387
rect 113604 -25395 113648 -25387
rect 113704 -25395 113748 -25387
rect 113804 -25395 113848 -25387
rect 113904 -25395 113948 -25387
rect 114004 -25395 114048 -25387
rect 114104 -25395 114148 -25387
rect 114204 -25395 114248 -25387
rect 114304 -25395 114348 -25387
rect 114404 -25395 114448 -25387
rect 114504 -25395 114548 -25387
rect 114604 -25395 114648 -25387
rect 115104 -25395 115148 -25387
rect 115204 -25395 115248 -25387
rect 115304 -25395 115348 -25387
rect 115404 -25395 115448 -25387
rect 115504 -25395 115548 -25387
rect 115604 -25395 115648 -25387
rect 115704 -25395 115748 -25387
rect 115804 -25395 115848 -25387
rect 115904 -25395 115948 -25387
rect 116004 -25395 116048 -25387
rect 116104 -25395 116148 -25387
rect 116204 -25395 116248 -25387
rect 116304 -25395 116348 -25387
rect 116404 -25395 116448 -25387
rect 116504 -25395 116548 -25387
rect 116604 -25395 116648 -25387
rect 80849 -25426 80893 -25418
rect 80949 -25426 80993 -25418
rect 81049 -25426 81093 -25418
rect 81149 -25426 81193 -25418
rect 81249 -25426 81293 -25418
rect 81349 -25426 81393 -25418
rect 81449 -25426 81493 -25418
rect 81549 -25426 81593 -25418
rect 81649 -25426 81693 -25418
rect 81749 -25426 81793 -25418
rect 81849 -25426 81893 -25418
rect 81949 -25426 81993 -25418
rect 82049 -25426 82093 -25418
rect 82149 -25426 82193 -25418
rect 82249 -25426 82293 -25418
rect 82349 -25426 82393 -25418
rect 82849 -25426 82893 -25418
rect 82949 -25426 82993 -25418
rect 83049 -25426 83093 -25418
rect 83149 -25426 83193 -25418
rect 83249 -25426 83293 -25418
rect 83349 -25426 83393 -25418
rect 83449 -25426 83493 -25418
rect 83549 -25426 83593 -25418
rect 83649 -25426 83693 -25418
rect 83749 -25426 83793 -25418
rect 83849 -25426 83893 -25418
rect 83949 -25426 83993 -25418
rect 84049 -25426 84093 -25418
rect 84149 -25426 84193 -25418
rect 84249 -25426 84293 -25418
rect 84349 -25426 84393 -25418
rect 84849 -25426 84893 -25418
rect 84949 -25426 84993 -25418
rect 85049 -25426 85093 -25418
rect 85149 -25426 85193 -25418
rect 85249 -25426 85293 -25418
rect 85349 -25426 85393 -25418
rect 85449 -25426 85493 -25418
rect 85549 -25426 85593 -25418
rect 85649 -25426 85693 -25418
rect 85749 -25426 85793 -25418
rect 85849 -25426 85893 -25418
rect 85949 -25426 85993 -25418
rect 86049 -25426 86093 -25418
rect 86149 -25426 86193 -25418
rect 86249 -25426 86293 -25418
rect 86349 -25426 86393 -25418
rect 86849 -25426 86893 -25418
rect 86949 -25426 86993 -25418
rect 87049 -25426 87093 -25418
rect 87149 -25426 87193 -25418
rect 87249 -25426 87293 -25418
rect 87349 -25426 87393 -25418
rect 87449 -25426 87493 -25418
rect 87549 -25426 87593 -25418
rect 87649 -25426 87693 -25418
rect 87749 -25426 87793 -25418
rect 87849 -25426 87893 -25418
rect 87949 -25426 87993 -25418
rect 88049 -25426 88093 -25418
rect 88149 -25426 88193 -25418
rect 88249 -25426 88293 -25418
rect 88349 -25426 88393 -25418
rect 80893 -25470 80901 -25426
rect 80993 -25470 81001 -25426
rect 81093 -25470 81101 -25426
rect 81193 -25470 81201 -25426
rect 81293 -25470 81301 -25426
rect 81393 -25470 81401 -25426
rect 81493 -25470 81501 -25426
rect 81593 -25470 81601 -25426
rect 81693 -25470 81701 -25426
rect 81793 -25470 81801 -25426
rect 81893 -25470 81901 -25426
rect 81993 -25470 82001 -25426
rect 82093 -25470 82101 -25426
rect 82193 -25470 82201 -25426
rect 82293 -25470 82301 -25426
rect 82393 -25470 82401 -25426
rect 82893 -25470 82901 -25426
rect 82993 -25470 83001 -25426
rect 83093 -25470 83101 -25426
rect 83193 -25470 83201 -25426
rect 83293 -25470 83301 -25426
rect 83393 -25470 83401 -25426
rect 83493 -25470 83501 -25426
rect 83593 -25470 83601 -25426
rect 83693 -25470 83701 -25426
rect 83793 -25470 83801 -25426
rect 83893 -25470 83901 -25426
rect 83993 -25470 84001 -25426
rect 84093 -25470 84101 -25426
rect 84193 -25470 84201 -25426
rect 84293 -25470 84301 -25426
rect 84393 -25470 84401 -25426
rect 84893 -25470 84901 -25426
rect 84993 -25470 85001 -25426
rect 85093 -25470 85101 -25426
rect 85193 -25470 85201 -25426
rect 85293 -25470 85301 -25426
rect 85393 -25470 85401 -25426
rect 85493 -25470 85501 -25426
rect 85593 -25470 85601 -25426
rect 85693 -25470 85701 -25426
rect 85793 -25470 85801 -25426
rect 85893 -25470 85901 -25426
rect 85993 -25470 86001 -25426
rect 86093 -25470 86101 -25426
rect 86193 -25470 86201 -25426
rect 86293 -25470 86301 -25426
rect 86393 -25470 86401 -25426
rect 86893 -25470 86901 -25426
rect 86993 -25470 87001 -25426
rect 87093 -25470 87101 -25426
rect 87193 -25470 87201 -25426
rect 87293 -25470 87301 -25426
rect 87393 -25470 87401 -25426
rect 87493 -25470 87501 -25426
rect 87593 -25470 87601 -25426
rect 87693 -25470 87701 -25426
rect 87793 -25470 87801 -25426
rect 87893 -25470 87901 -25426
rect 87993 -25470 88001 -25426
rect 88093 -25470 88101 -25426
rect 88193 -25470 88201 -25426
rect 88293 -25470 88301 -25426
rect 88393 -25470 88401 -25426
rect 109148 -25439 109156 -25395
rect 109248 -25439 109256 -25395
rect 109348 -25439 109356 -25395
rect 109448 -25439 109456 -25395
rect 109548 -25439 109556 -25395
rect 109648 -25439 109656 -25395
rect 109748 -25439 109756 -25395
rect 109848 -25439 109856 -25395
rect 109948 -25439 109956 -25395
rect 110048 -25439 110056 -25395
rect 110148 -25439 110156 -25395
rect 110248 -25439 110256 -25395
rect 110348 -25439 110356 -25395
rect 110448 -25439 110456 -25395
rect 110548 -25439 110556 -25395
rect 110648 -25439 110656 -25395
rect 111148 -25439 111156 -25395
rect 111248 -25439 111256 -25395
rect 111348 -25439 111356 -25395
rect 111448 -25439 111456 -25395
rect 111548 -25439 111556 -25395
rect 111648 -25439 111656 -25395
rect 111748 -25439 111756 -25395
rect 111848 -25439 111856 -25395
rect 111948 -25439 111956 -25395
rect 112048 -25439 112056 -25395
rect 112148 -25439 112156 -25395
rect 112248 -25439 112256 -25395
rect 112348 -25439 112356 -25395
rect 112448 -25439 112456 -25395
rect 112548 -25439 112556 -25395
rect 112648 -25439 112656 -25395
rect 113148 -25439 113156 -25395
rect 113248 -25439 113256 -25395
rect 113348 -25439 113356 -25395
rect 113448 -25439 113456 -25395
rect 113548 -25439 113556 -25395
rect 113648 -25439 113656 -25395
rect 113748 -25439 113756 -25395
rect 113848 -25439 113856 -25395
rect 113948 -25439 113956 -25395
rect 114048 -25439 114056 -25395
rect 114148 -25439 114156 -25395
rect 114248 -25439 114256 -25395
rect 114348 -25439 114356 -25395
rect 114448 -25439 114456 -25395
rect 114548 -25439 114556 -25395
rect 114648 -25439 114656 -25395
rect 115148 -25439 115156 -25395
rect 115248 -25439 115256 -25395
rect 115348 -25439 115356 -25395
rect 115448 -25439 115456 -25395
rect 115548 -25439 115556 -25395
rect 115648 -25439 115656 -25395
rect 115748 -25439 115756 -25395
rect 115848 -25439 115856 -25395
rect 115948 -25439 115956 -25395
rect 116048 -25439 116056 -25395
rect 116148 -25439 116156 -25395
rect 116248 -25439 116256 -25395
rect 116348 -25439 116356 -25395
rect 116448 -25439 116456 -25395
rect 116548 -25439 116556 -25395
rect 116648 -25439 116656 -25395
rect 109104 -25495 109148 -25487
rect 109204 -25495 109248 -25487
rect 109304 -25495 109348 -25487
rect 109404 -25495 109448 -25487
rect 109504 -25495 109548 -25487
rect 109604 -25495 109648 -25487
rect 109704 -25495 109748 -25487
rect 109804 -25495 109848 -25487
rect 109904 -25495 109948 -25487
rect 110004 -25495 110048 -25487
rect 110104 -25495 110148 -25487
rect 110204 -25495 110248 -25487
rect 110304 -25495 110348 -25487
rect 110404 -25495 110448 -25487
rect 110504 -25495 110548 -25487
rect 110604 -25495 110648 -25487
rect 111104 -25495 111148 -25487
rect 111204 -25495 111248 -25487
rect 111304 -25495 111348 -25487
rect 111404 -25495 111448 -25487
rect 111504 -25495 111548 -25487
rect 111604 -25495 111648 -25487
rect 111704 -25495 111748 -25487
rect 111804 -25495 111848 -25487
rect 111904 -25495 111948 -25487
rect 112004 -25495 112048 -25487
rect 112104 -25495 112148 -25487
rect 112204 -25495 112248 -25487
rect 112304 -25495 112348 -25487
rect 112404 -25495 112448 -25487
rect 112504 -25495 112548 -25487
rect 112604 -25495 112648 -25487
rect 113104 -25495 113148 -25487
rect 113204 -25495 113248 -25487
rect 113304 -25495 113348 -25487
rect 113404 -25495 113448 -25487
rect 113504 -25495 113548 -25487
rect 113604 -25495 113648 -25487
rect 113704 -25495 113748 -25487
rect 113804 -25495 113848 -25487
rect 113904 -25495 113948 -25487
rect 114004 -25495 114048 -25487
rect 114104 -25495 114148 -25487
rect 114204 -25495 114248 -25487
rect 114304 -25495 114348 -25487
rect 114404 -25495 114448 -25487
rect 114504 -25495 114548 -25487
rect 114604 -25495 114648 -25487
rect 115104 -25495 115148 -25487
rect 115204 -25495 115248 -25487
rect 115304 -25495 115348 -25487
rect 115404 -25495 115448 -25487
rect 115504 -25495 115548 -25487
rect 115604 -25495 115648 -25487
rect 115704 -25495 115748 -25487
rect 115804 -25495 115848 -25487
rect 115904 -25495 115948 -25487
rect 116004 -25495 116048 -25487
rect 116104 -25495 116148 -25487
rect 116204 -25495 116248 -25487
rect 116304 -25495 116348 -25487
rect 116404 -25495 116448 -25487
rect 116504 -25495 116548 -25487
rect 116604 -25495 116648 -25487
rect 80849 -25526 80893 -25518
rect 80949 -25526 80993 -25518
rect 81049 -25526 81093 -25518
rect 81149 -25526 81193 -25518
rect 81249 -25526 81293 -25518
rect 81349 -25526 81393 -25518
rect 81449 -25526 81493 -25518
rect 81549 -25526 81593 -25518
rect 81649 -25526 81693 -25518
rect 81749 -25526 81793 -25518
rect 81849 -25526 81893 -25518
rect 81949 -25526 81993 -25518
rect 82049 -25526 82093 -25518
rect 82149 -25526 82193 -25518
rect 82249 -25526 82293 -25518
rect 82349 -25526 82393 -25518
rect 82849 -25526 82893 -25518
rect 82949 -25526 82993 -25518
rect 83049 -25526 83093 -25518
rect 83149 -25526 83193 -25518
rect 83249 -25526 83293 -25518
rect 83349 -25526 83393 -25518
rect 83449 -25526 83493 -25518
rect 83549 -25526 83593 -25518
rect 83649 -25526 83693 -25518
rect 83749 -25526 83793 -25518
rect 83849 -25526 83893 -25518
rect 83949 -25526 83993 -25518
rect 84049 -25526 84093 -25518
rect 84149 -25526 84193 -25518
rect 84249 -25526 84293 -25518
rect 84349 -25526 84393 -25518
rect 84849 -25526 84893 -25518
rect 84949 -25526 84993 -25518
rect 85049 -25526 85093 -25518
rect 85149 -25526 85193 -25518
rect 85249 -25526 85293 -25518
rect 85349 -25526 85393 -25518
rect 85449 -25526 85493 -25518
rect 85549 -25526 85593 -25518
rect 85649 -25526 85693 -25518
rect 85749 -25526 85793 -25518
rect 85849 -25526 85893 -25518
rect 85949 -25526 85993 -25518
rect 86049 -25526 86093 -25518
rect 86149 -25526 86193 -25518
rect 86249 -25526 86293 -25518
rect 86349 -25526 86393 -25518
rect 86849 -25526 86893 -25518
rect 86949 -25526 86993 -25518
rect 87049 -25526 87093 -25518
rect 87149 -25526 87193 -25518
rect 87249 -25526 87293 -25518
rect 87349 -25526 87393 -25518
rect 87449 -25526 87493 -25518
rect 87549 -25526 87593 -25518
rect 87649 -25526 87693 -25518
rect 87749 -25526 87793 -25518
rect 87849 -25526 87893 -25518
rect 87949 -25526 87993 -25518
rect 88049 -25526 88093 -25518
rect 88149 -25526 88193 -25518
rect 88249 -25526 88293 -25518
rect 88349 -25526 88393 -25518
rect 80893 -25570 80901 -25526
rect 80993 -25570 81001 -25526
rect 81093 -25570 81101 -25526
rect 81193 -25570 81201 -25526
rect 81293 -25570 81301 -25526
rect 81393 -25570 81401 -25526
rect 81493 -25570 81501 -25526
rect 81593 -25570 81601 -25526
rect 81693 -25570 81701 -25526
rect 81793 -25570 81801 -25526
rect 81893 -25570 81901 -25526
rect 81993 -25570 82001 -25526
rect 82093 -25570 82101 -25526
rect 82193 -25570 82201 -25526
rect 82293 -25570 82301 -25526
rect 82393 -25570 82401 -25526
rect 82893 -25570 82901 -25526
rect 82993 -25570 83001 -25526
rect 83093 -25570 83101 -25526
rect 83193 -25570 83201 -25526
rect 83293 -25570 83301 -25526
rect 83393 -25570 83401 -25526
rect 83493 -25570 83501 -25526
rect 83593 -25570 83601 -25526
rect 83693 -25570 83701 -25526
rect 83793 -25570 83801 -25526
rect 83893 -25570 83901 -25526
rect 83993 -25570 84001 -25526
rect 84093 -25570 84101 -25526
rect 84193 -25570 84201 -25526
rect 84293 -25570 84301 -25526
rect 84393 -25570 84401 -25526
rect 84893 -25570 84901 -25526
rect 84993 -25570 85001 -25526
rect 85093 -25570 85101 -25526
rect 85193 -25570 85201 -25526
rect 85293 -25570 85301 -25526
rect 85393 -25570 85401 -25526
rect 85493 -25570 85501 -25526
rect 85593 -25570 85601 -25526
rect 85693 -25570 85701 -25526
rect 85793 -25570 85801 -25526
rect 85893 -25570 85901 -25526
rect 85993 -25570 86001 -25526
rect 86093 -25570 86101 -25526
rect 86193 -25570 86201 -25526
rect 86293 -25570 86301 -25526
rect 86393 -25570 86401 -25526
rect 86893 -25570 86901 -25526
rect 86993 -25570 87001 -25526
rect 87093 -25570 87101 -25526
rect 87193 -25570 87201 -25526
rect 87293 -25570 87301 -25526
rect 87393 -25570 87401 -25526
rect 87493 -25570 87501 -25526
rect 87593 -25570 87601 -25526
rect 87693 -25570 87701 -25526
rect 87793 -25570 87801 -25526
rect 87893 -25570 87901 -25526
rect 87993 -25570 88001 -25526
rect 88093 -25570 88101 -25526
rect 88193 -25570 88201 -25526
rect 88293 -25570 88301 -25526
rect 88393 -25570 88401 -25526
rect 109148 -25539 109156 -25495
rect 109248 -25539 109256 -25495
rect 109348 -25539 109356 -25495
rect 109448 -25539 109456 -25495
rect 109548 -25539 109556 -25495
rect 109648 -25539 109656 -25495
rect 109748 -25539 109756 -25495
rect 109848 -25539 109856 -25495
rect 109948 -25539 109956 -25495
rect 110048 -25539 110056 -25495
rect 110148 -25539 110156 -25495
rect 110248 -25539 110256 -25495
rect 110348 -25539 110356 -25495
rect 110448 -25539 110456 -25495
rect 110548 -25539 110556 -25495
rect 110648 -25539 110656 -25495
rect 111148 -25539 111156 -25495
rect 111248 -25539 111256 -25495
rect 111348 -25539 111356 -25495
rect 111448 -25539 111456 -25495
rect 111548 -25539 111556 -25495
rect 111648 -25539 111656 -25495
rect 111748 -25539 111756 -25495
rect 111848 -25539 111856 -25495
rect 111948 -25539 111956 -25495
rect 112048 -25539 112056 -25495
rect 112148 -25539 112156 -25495
rect 112248 -25539 112256 -25495
rect 112348 -25539 112356 -25495
rect 112448 -25539 112456 -25495
rect 112548 -25539 112556 -25495
rect 112648 -25539 112656 -25495
rect 113148 -25539 113156 -25495
rect 113248 -25539 113256 -25495
rect 113348 -25539 113356 -25495
rect 113448 -25539 113456 -25495
rect 113548 -25539 113556 -25495
rect 113648 -25539 113656 -25495
rect 113748 -25539 113756 -25495
rect 113848 -25539 113856 -25495
rect 113948 -25539 113956 -25495
rect 114048 -25539 114056 -25495
rect 114148 -25539 114156 -25495
rect 114248 -25539 114256 -25495
rect 114348 -25539 114356 -25495
rect 114448 -25539 114456 -25495
rect 114548 -25539 114556 -25495
rect 114648 -25539 114656 -25495
rect 115148 -25539 115156 -25495
rect 115248 -25539 115256 -25495
rect 115348 -25539 115356 -25495
rect 115448 -25539 115456 -25495
rect 115548 -25539 115556 -25495
rect 115648 -25539 115656 -25495
rect 115748 -25539 115756 -25495
rect 115848 -25539 115856 -25495
rect 115948 -25539 115956 -25495
rect 116048 -25539 116056 -25495
rect 116148 -25539 116156 -25495
rect 116248 -25539 116256 -25495
rect 116348 -25539 116356 -25495
rect 116448 -25539 116456 -25495
rect 116548 -25539 116556 -25495
rect 116648 -25539 116656 -25495
rect 109104 -25595 109148 -25587
rect 109204 -25595 109248 -25587
rect 109304 -25595 109348 -25587
rect 109404 -25595 109448 -25587
rect 109504 -25595 109548 -25587
rect 109604 -25595 109648 -25587
rect 109704 -25595 109748 -25587
rect 109804 -25595 109848 -25587
rect 109904 -25595 109948 -25587
rect 110004 -25595 110048 -25587
rect 110104 -25595 110148 -25587
rect 110204 -25595 110248 -25587
rect 110304 -25595 110348 -25587
rect 110404 -25595 110448 -25587
rect 110504 -25595 110548 -25587
rect 110604 -25595 110648 -25587
rect 111104 -25595 111148 -25587
rect 111204 -25595 111248 -25587
rect 111304 -25595 111348 -25587
rect 111404 -25595 111448 -25587
rect 111504 -25595 111548 -25587
rect 111604 -25595 111648 -25587
rect 111704 -25595 111748 -25587
rect 111804 -25595 111848 -25587
rect 111904 -25595 111948 -25587
rect 112004 -25595 112048 -25587
rect 112104 -25595 112148 -25587
rect 112204 -25595 112248 -25587
rect 112304 -25595 112348 -25587
rect 112404 -25595 112448 -25587
rect 112504 -25595 112548 -25587
rect 112604 -25595 112648 -25587
rect 113104 -25595 113148 -25587
rect 113204 -25595 113248 -25587
rect 113304 -25595 113348 -25587
rect 113404 -25595 113448 -25587
rect 113504 -25595 113548 -25587
rect 113604 -25595 113648 -25587
rect 113704 -25595 113748 -25587
rect 113804 -25595 113848 -25587
rect 113904 -25595 113948 -25587
rect 114004 -25595 114048 -25587
rect 114104 -25595 114148 -25587
rect 114204 -25595 114248 -25587
rect 114304 -25595 114348 -25587
rect 114404 -25595 114448 -25587
rect 114504 -25595 114548 -25587
rect 114604 -25595 114648 -25587
rect 115104 -25595 115148 -25587
rect 115204 -25595 115248 -25587
rect 115304 -25595 115348 -25587
rect 115404 -25595 115448 -25587
rect 115504 -25595 115548 -25587
rect 115604 -25595 115648 -25587
rect 115704 -25595 115748 -25587
rect 115804 -25595 115848 -25587
rect 115904 -25595 115948 -25587
rect 116004 -25595 116048 -25587
rect 116104 -25595 116148 -25587
rect 116204 -25595 116248 -25587
rect 116304 -25595 116348 -25587
rect 116404 -25595 116448 -25587
rect 116504 -25595 116548 -25587
rect 116604 -25595 116648 -25587
rect 109148 -25639 109156 -25595
rect 109248 -25639 109256 -25595
rect 109348 -25639 109356 -25595
rect 109448 -25639 109456 -25595
rect 109548 -25639 109556 -25595
rect 109648 -25639 109656 -25595
rect 109748 -25639 109756 -25595
rect 109848 -25639 109856 -25595
rect 109948 -25639 109956 -25595
rect 110048 -25639 110056 -25595
rect 110148 -25639 110156 -25595
rect 110248 -25639 110256 -25595
rect 110348 -25639 110356 -25595
rect 110448 -25639 110456 -25595
rect 110548 -25639 110556 -25595
rect 110648 -25639 110656 -25595
rect 111148 -25639 111156 -25595
rect 111248 -25639 111256 -25595
rect 111348 -25639 111356 -25595
rect 111448 -25639 111456 -25595
rect 111548 -25639 111556 -25595
rect 111648 -25639 111656 -25595
rect 111748 -25639 111756 -25595
rect 111848 -25639 111856 -25595
rect 111948 -25639 111956 -25595
rect 112048 -25639 112056 -25595
rect 112148 -25639 112156 -25595
rect 112248 -25639 112256 -25595
rect 112348 -25639 112356 -25595
rect 112448 -25639 112456 -25595
rect 112548 -25639 112556 -25595
rect 112648 -25639 112656 -25595
rect 113148 -25639 113156 -25595
rect 113248 -25639 113256 -25595
rect 113348 -25639 113356 -25595
rect 113448 -25639 113456 -25595
rect 113548 -25639 113556 -25595
rect 113648 -25639 113656 -25595
rect 113748 -25639 113756 -25595
rect 113848 -25639 113856 -25595
rect 113948 -25639 113956 -25595
rect 114048 -25639 114056 -25595
rect 114148 -25639 114156 -25595
rect 114248 -25639 114256 -25595
rect 114348 -25639 114356 -25595
rect 114448 -25639 114456 -25595
rect 114548 -25639 114556 -25595
rect 114648 -25639 114656 -25595
rect 115148 -25639 115156 -25595
rect 115248 -25639 115256 -25595
rect 115348 -25639 115356 -25595
rect 115448 -25639 115456 -25595
rect 115548 -25639 115556 -25595
rect 115648 -25639 115656 -25595
rect 115748 -25639 115756 -25595
rect 115848 -25639 115856 -25595
rect 115948 -25639 115956 -25595
rect 116048 -25639 116056 -25595
rect 116148 -25639 116156 -25595
rect 116248 -25639 116256 -25595
rect 116348 -25639 116356 -25595
rect 116448 -25639 116456 -25595
rect 116548 -25639 116556 -25595
rect 116648 -25639 116656 -25595
rect 109104 -25695 109148 -25687
rect 109204 -25695 109248 -25687
rect 109304 -25695 109348 -25687
rect 109404 -25695 109448 -25687
rect 109504 -25695 109548 -25687
rect 109604 -25695 109648 -25687
rect 109704 -25695 109748 -25687
rect 109804 -25695 109848 -25687
rect 109904 -25695 109948 -25687
rect 110004 -25695 110048 -25687
rect 110104 -25695 110148 -25687
rect 110204 -25695 110248 -25687
rect 110304 -25695 110348 -25687
rect 110404 -25695 110448 -25687
rect 110504 -25695 110548 -25687
rect 110604 -25695 110648 -25687
rect 111104 -25695 111148 -25687
rect 111204 -25695 111248 -25687
rect 111304 -25695 111348 -25687
rect 111404 -25695 111448 -25687
rect 111504 -25695 111548 -25687
rect 111604 -25695 111648 -25687
rect 111704 -25695 111748 -25687
rect 111804 -25695 111848 -25687
rect 111904 -25695 111948 -25687
rect 112004 -25695 112048 -25687
rect 112104 -25695 112148 -25687
rect 112204 -25695 112248 -25687
rect 112304 -25695 112348 -25687
rect 112404 -25695 112448 -25687
rect 112504 -25695 112548 -25687
rect 112604 -25695 112648 -25687
rect 113104 -25695 113148 -25687
rect 113204 -25695 113248 -25687
rect 113304 -25695 113348 -25687
rect 113404 -25695 113448 -25687
rect 113504 -25695 113548 -25687
rect 113604 -25695 113648 -25687
rect 113704 -25695 113748 -25687
rect 113804 -25695 113848 -25687
rect 113904 -25695 113948 -25687
rect 114004 -25695 114048 -25687
rect 114104 -25695 114148 -25687
rect 114204 -25695 114248 -25687
rect 114304 -25695 114348 -25687
rect 114404 -25695 114448 -25687
rect 114504 -25695 114548 -25687
rect 114604 -25695 114648 -25687
rect 115104 -25695 115148 -25687
rect 115204 -25695 115248 -25687
rect 115304 -25695 115348 -25687
rect 115404 -25695 115448 -25687
rect 115504 -25695 115548 -25687
rect 115604 -25695 115648 -25687
rect 115704 -25695 115748 -25687
rect 115804 -25695 115848 -25687
rect 115904 -25695 115948 -25687
rect 116004 -25695 116048 -25687
rect 116104 -25695 116148 -25687
rect 116204 -25695 116248 -25687
rect 116304 -25695 116348 -25687
rect 116404 -25695 116448 -25687
rect 116504 -25695 116548 -25687
rect 116604 -25695 116648 -25687
rect 109148 -25739 109156 -25695
rect 109248 -25739 109256 -25695
rect 109348 -25739 109356 -25695
rect 109448 -25739 109456 -25695
rect 109548 -25739 109556 -25695
rect 109648 -25739 109656 -25695
rect 109748 -25739 109756 -25695
rect 109848 -25739 109856 -25695
rect 109948 -25739 109956 -25695
rect 110048 -25739 110056 -25695
rect 110148 -25739 110156 -25695
rect 110248 -25739 110256 -25695
rect 110348 -25739 110356 -25695
rect 110448 -25739 110456 -25695
rect 110548 -25739 110556 -25695
rect 110648 -25739 110656 -25695
rect 111148 -25739 111156 -25695
rect 111248 -25739 111256 -25695
rect 111348 -25739 111356 -25695
rect 111448 -25739 111456 -25695
rect 111548 -25739 111556 -25695
rect 111648 -25739 111656 -25695
rect 111748 -25739 111756 -25695
rect 111848 -25739 111856 -25695
rect 111948 -25739 111956 -25695
rect 112048 -25739 112056 -25695
rect 112148 -25739 112156 -25695
rect 112248 -25739 112256 -25695
rect 112348 -25739 112356 -25695
rect 112448 -25739 112456 -25695
rect 112548 -25739 112556 -25695
rect 112648 -25739 112656 -25695
rect 113148 -25739 113156 -25695
rect 113248 -25739 113256 -25695
rect 113348 -25739 113356 -25695
rect 113448 -25739 113456 -25695
rect 113548 -25739 113556 -25695
rect 113648 -25739 113656 -25695
rect 113748 -25739 113756 -25695
rect 113848 -25739 113856 -25695
rect 113948 -25739 113956 -25695
rect 114048 -25739 114056 -25695
rect 114148 -25739 114156 -25695
rect 114248 -25739 114256 -25695
rect 114348 -25739 114356 -25695
rect 114448 -25739 114456 -25695
rect 114548 -25739 114556 -25695
rect 114648 -25739 114656 -25695
rect 115148 -25739 115156 -25695
rect 115248 -25739 115256 -25695
rect 115348 -25739 115356 -25695
rect 115448 -25739 115456 -25695
rect 115548 -25739 115556 -25695
rect 115648 -25739 115656 -25695
rect 115748 -25739 115756 -25695
rect 115848 -25739 115856 -25695
rect 115948 -25739 115956 -25695
rect 116048 -25739 116056 -25695
rect 116148 -25739 116156 -25695
rect 116248 -25739 116256 -25695
rect 116348 -25739 116356 -25695
rect 116448 -25739 116456 -25695
rect 116548 -25739 116556 -25695
rect 116648 -25739 116656 -25695
rect -109180 -48119 -109178 -28119
rect -109114 -48119 -109112 -28119
rect -77180 -48119 -77178 -28119
rect -77114 -48119 -77112 -28119
rect -45180 -48119 -45178 -28119
rect -45114 -48119 -45112 -28119
rect -13180 -48119 -13178 -28119
rect -13114 -48119 -13112 -28119
rect 18820 -48119 18822 -28119
rect 18886 -48119 18888 -28119
rect 50820 -48119 50822 -28119
rect 50886 -48119 50888 -28119
rect 82820 -48119 82822 -28119
rect 82886 -48119 82888 -28119
rect 114820 -48119 114822 -28119
rect 114886 -48119 114888 -28119
rect 146820 -48119 146822 -28119
rect 146886 -48119 146888 -28119
rect 109305 -51137 109349 -51129
rect 109405 -51137 109449 -51129
rect 109505 -51137 109549 -51129
rect 109605 -51137 109649 -51129
rect 109705 -51137 109749 -51129
rect 109805 -51137 109849 -51129
rect 109905 -51137 109949 -51129
rect 110005 -51137 110049 -51129
rect 110105 -51137 110149 -51129
rect 110205 -51137 110249 -51129
rect 110305 -51137 110349 -51129
rect 110405 -51137 110449 -51129
rect 110505 -51137 110549 -51129
rect 110605 -51137 110649 -51129
rect 110705 -51137 110749 -51129
rect 110805 -51137 110849 -51129
rect 111305 -51137 111349 -51129
rect 111405 -51137 111449 -51129
rect 111505 -51137 111549 -51129
rect 111605 -51137 111649 -51129
rect 111705 -51137 111749 -51129
rect 111805 -51137 111849 -51129
rect 111905 -51137 111949 -51129
rect 112005 -51137 112049 -51129
rect 112105 -51137 112149 -51129
rect 112205 -51137 112249 -51129
rect 112305 -51137 112349 -51129
rect 112405 -51137 112449 -51129
rect 112505 -51137 112549 -51129
rect 112605 -51137 112649 -51129
rect 112705 -51137 112749 -51129
rect 112805 -51137 112849 -51129
rect 113305 -51137 113349 -51129
rect 113405 -51137 113449 -51129
rect 113505 -51137 113549 -51129
rect 113605 -51137 113649 -51129
rect 113705 -51137 113749 -51129
rect 113805 -51137 113849 -51129
rect 113905 -51137 113949 -51129
rect 114005 -51137 114049 -51129
rect 114105 -51137 114149 -51129
rect 114205 -51137 114249 -51129
rect 114305 -51137 114349 -51129
rect 114405 -51137 114449 -51129
rect 114505 -51137 114549 -51129
rect 114605 -51137 114649 -51129
rect 114705 -51137 114749 -51129
rect 114805 -51137 114849 -51129
rect 115305 -51137 115349 -51129
rect 115405 -51137 115449 -51129
rect 115505 -51137 115549 -51129
rect 115605 -51137 115649 -51129
rect 115705 -51137 115749 -51129
rect 115805 -51137 115849 -51129
rect 115905 -51137 115949 -51129
rect 116005 -51137 116049 -51129
rect 116105 -51137 116149 -51129
rect 116205 -51137 116249 -51129
rect 116305 -51137 116349 -51129
rect 116405 -51137 116449 -51129
rect 116505 -51137 116549 -51129
rect 116605 -51137 116649 -51129
rect 116705 -51137 116749 -51129
rect 116805 -51137 116849 -51129
rect 109349 -51181 109357 -51137
rect 109449 -51181 109457 -51137
rect 109549 -51181 109557 -51137
rect 109649 -51181 109657 -51137
rect 109749 -51181 109757 -51137
rect 109849 -51181 109857 -51137
rect 109949 -51181 109957 -51137
rect 110049 -51181 110057 -51137
rect 110149 -51181 110157 -51137
rect 110249 -51181 110257 -51137
rect 110349 -51181 110357 -51137
rect 110449 -51181 110457 -51137
rect 110549 -51181 110557 -51137
rect 110649 -51181 110657 -51137
rect 110749 -51181 110757 -51137
rect 110849 -51181 110857 -51137
rect 111349 -51181 111357 -51137
rect 111449 -51181 111457 -51137
rect 111549 -51181 111557 -51137
rect 111649 -51181 111657 -51137
rect 111749 -51181 111757 -51137
rect 111849 -51181 111857 -51137
rect 111949 -51181 111957 -51137
rect 112049 -51181 112057 -51137
rect 112149 -51181 112157 -51137
rect 112249 -51181 112257 -51137
rect 112349 -51181 112357 -51137
rect 112449 -51181 112457 -51137
rect 112549 -51181 112557 -51137
rect 112649 -51181 112657 -51137
rect 112749 -51181 112757 -51137
rect 112849 -51181 112857 -51137
rect 113349 -51181 113357 -51137
rect 113449 -51181 113457 -51137
rect 113549 -51181 113557 -51137
rect 113649 -51181 113657 -51137
rect 113749 -51181 113757 -51137
rect 113849 -51181 113857 -51137
rect 113949 -51181 113957 -51137
rect 114049 -51181 114057 -51137
rect 114149 -51181 114157 -51137
rect 114249 -51181 114257 -51137
rect 114349 -51181 114357 -51137
rect 114449 -51181 114457 -51137
rect 114549 -51181 114557 -51137
rect 114649 -51181 114657 -51137
rect 114749 -51181 114757 -51137
rect 114849 -51181 114857 -51137
rect 115349 -51181 115357 -51137
rect 115449 -51181 115457 -51137
rect 115549 -51181 115557 -51137
rect 115649 -51181 115657 -51137
rect 115749 -51181 115757 -51137
rect 115849 -51181 115857 -51137
rect 115949 -51181 115957 -51137
rect 116049 -51181 116057 -51137
rect 116149 -51181 116157 -51137
rect 116249 -51181 116257 -51137
rect 116349 -51181 116357 -51137
rect 116449 -51181 116457 -51137
rect 116549 -51181 116557 -51137
rect 116649 -51181 116657 -51137
rect 116749 -51181 116757 -51137
rect 116849 -51181 116857 -51137
rect 109305 -51237 109349 -51229
rect 109405 -51237 109449 -51229
rect 109505 -51237 109549 -51229
rect 109605 -51237 109649 -51229
rect 109705 -51237 109749 -51229
rect 109805 -51237 109849 -51229
rect 109905 -51237 109949 -51229
rect 110005 -51237 110049 -51229
rect 110105 -51237 110149 -51229
rect 110205 -51237 110249 -51229
rect 110305 -51237 110349 -51229
rect 110405 -51237 110449 -51229
rect 110505 -51237 110549 -51229
rect 110605 -51237 110649 -51229
rect 110705 -51237 110749 -51229
rect 110805 -51237 110849 -51229
rect 111305 -51237 111349 -51229
rect 111405 -51237 111449 -51229
rect 111505 -51237 111549 -51229
rect 111605 -51237 111649 -51229
rect 111705 -51237 111749 -51229
rect 111805 -51237 111849 -51229
rect 111905 -51237 111949 -51229
rect 112005 -51237 112049 -51229
rect 112105 -51237 112149 -51229
rect 112205 -51237 112249 -51229
rect 112305 -51237 112349 -51229
rect 112405 -51237 112449 -51229
rect 112505 -51237 112549 -51229
rect 112605 -51237 112649 -51229
rect 112705 -51237 112749 -51229
rect 112805 -51237 112849 -51229
rect 113305 -51237 113349 -51229
rect 113405 -51237 113449 -51229
rect 113505 -51237 113549 -51229
rect 113605 -51237 113649 -51229
rect 113705 -51237 113749 -51229
rect 113805 -51237 113849 -51229
rect 113905 -51237 113949 -51229
rect 114005 -51237 114049 -51229
rect 114105 -51237 114149 -51229
rect 114205 -51237 114249 -51229
rect 114305 -51237 114349 -51229
rect 114405 -51237 114449 -51229
rect 114505 -51237 114549 -51229
rect 114605 -51237 114649 -51229
rect 114705 -51237 114749 -51229
rect 114805 -51237 114849 -51229
rect 115305 -51237 115349 -51229
rect 115405 -51237 115449 -51229
rect 115505 -51237 115549 -51229
rect 115605 -51237 115649 -51229
rect 115705 -51237 115749 -51229
rect 115805 -51237 115849 -51229
rect 115905 -51237 115949 -51229
rect 116005 -51237 116049 -51229
rect 116105 -51237 116149 -51229
rect 116205 -51237 116249 -51229
rect 116305 -51237 116349 -51229
rect 116405 -51237 116449 -51229
rect 116505 -51237 116549 -51229
rect 116605 -51237 116649 -51229
rect 116705 -51237 116749 -51229
rect 116805 -51237 116849 -51229
rect 109349 -51281 109357 -51237
rect 109449 -51281 109457 -51237
rect 109549 -51281 109557 -51237
rect 109649 -51281 109657 -51237
rect 109749 -51281 109757 -51237
rect 109849 -51281 109857 -51237
rect 109949 -51281 109957 -51237
rect 110049 -51281 110057 -51237
rect 110149 -51281 110157 -51237
rect 110249 -51281 110257 -51237
rect 110349 -51281 110357 -51237
rect 110449 -51281 110457 -51237
rect 110549 -51281 110557 -51237
rect 110649 -51281 110657 -51237
rect 110749 -51281 110757 -51237
rect 110849 -51281 110857 -51237
rect 111349 -51281 111357 -51237
rect 111449 -51281 111457 -51237
rect 111549 -51281 111557 -51237
rect 111649 -51281 111657 -51237
rect 111749 -51281 111757 -51237
rect 111849 -51281 111857 -51237
rect 111949 -51281 111957 -51237
rect 112049 -51281 112057 -51237
rect 112149 -51281 112157 -51237
rect 112249 -51281 112257 -51237
rect 112349 -51281 112357 -51237
rect 112449 -51281 112457 -51237
rect 112549 -51281 112557 -51237
rect 112649 -51281 112657 -51237
rect 112749 -51281 112757 -51237
rect 112849 -51281 112857 -51237
rect 113349 -51281 113357 -51237
rect 113449 -51281 113457 -51237
rect 113549 -51281 113557 -51237
rect 113649 -51281 113657 -51237
rect 113749 -51281 113757 -51237
rect 113849 -51281 113857 -51237
rect 113949 -51281 113957 -51237
rect 114049 -51281 114057 -51237
rect 114149 -51281 114157 -51237
rect 114249 -51281 114257 -51237
rect 114349 -51281 114357 -51237
rect 114449 -51281 114457 -51237
rect 114549 -51281 114557 -51237
rect 114649 -51281 114657 -51237
rect 114749 -51281 114757 -51237
rect 114849 -51281 114857 -51237
rect 115349 -51281 115357 -51237
rect 115449 -51281 115457 -51237
rect 115549 -51281 115557 -51237
rect 115649 -51281 115657 -51237
rect 115749 -51281 115757 -51237
rect 115849 -51281 115857 -51237
rect 115949 -51281 115957 -51237
rect 116049 -51281 116057 -51237
rect 116149 -51281 116157 -51237
rect 116249 -51281 116257 -51237
rect 116349 -51281 116357 -51237
rect 116449 -51281 116457 -51237
rect 116549 -51281 116557 -51237
rect 116649 -51281 116657 -51237
rect 116749 -51281 116757 -51237
rect 116849 -51281 116857 -51237
rect 109305 -51337 109349 -51329
rect 109405 -51337 109449 -51329
rect 109505 -51337 109549 -51329
rect 109605 -51337 109649 -51329
rect 109705 -51337 109749 -51329
rect 109805 -51337 109849 -51329
rect 109905 -51337 109949 -51329
rect 110005 -51337 110049 -51329
rect 110105 -51337 110149 -51329
rect 110205 -51337 110249 -51329
rect 110305 -51337 110349 -51329
rect 110405 -51337 110449 -51329
rect 110505 -51337 110549 -51329
rect 110605 -51337 110649 -51329
rect 110705 -51337 110749 -51329
rect 110805 -51337 110849 -51329
rect 111305 -51337 111349 -51329
rect 111405 -51337 111449 -51329
rect 111505 -51337 111549 -51329
rect 111605 -51337 111649 -51329
rect 111705 -51337 111749 -51329
rect 111805 -51337 111849 -51329
rect 111905 -51337 111949 -51329
rect 112005 -51337 112049 -51329
rect 112105 -51337 112149 -51329
rect 112205 -51337 112249 -51329
rect 112305 -51337 112349 -51329
rect 112405 -51337 112449 -51329
rect 112505 -51337 112549 -51329
rect 112605 -51337 112649 -51329
rect 112705 -51337 112749 -51329
rect 112805 -51337 112849 -51329
rect 113305 -51337 113349 -51329
rect 113405 -51337 113449 -51329
rect 113505 -51337 113549 -51329
rect 113605 -51337 113649 -51329
rect 113705 -51337 113749 -51329
rect 113805 -51337 113849 -51329
rect 113905 -51337 113949 -51329
rect 114005 -51337 114049 -51329
rect 114105 -51337 114149 -51329
rect 114205 -51337 114249 -51329
rect 114305 -51337 114349 -51329
rect 114405 -51337 114449 -51329
rect 114505 -51337 114549 -51329
rect 114605 -51337 114649 -51329
rect 114705 -51337 114749 -51329
rect 114805 -51337 114849 -51329
rect 115305 -51337 115349 -51329
rect 115405 -51337 115449 -51329
rect 115505 -51337 115549 -51329
rect 115605 -51337 115649 -51329
rect 115705 -51337 115749 -51329
rect 115805 -51337 115849 -51329
rect 115905 -51337 115949 -51329
rect 116005 -51337 116049 -51329
rect 116105 -51337 116149 -51329
rect 116205 -51337 116249 -51329
rect 116305 -51337 116349 -51329
rect 116405 -51337 116449 -51329
rect 116505 -51337 116549 -51329
rect 116605 -51337 116649 -51329
rect 116705 -51337 116749 -51329
rect 116805 -51337 116849 -51329
rect 109349 -51381 109357 -51337
rect 109449 -51381 109457 -51337
rect 109549 -51381 109557 -51337
rect 109649 -51381 109657 -51337
rect 109749 -51381 109757 -51337
rect 109849 -51381 109857 -51337
rect 109949 -51381 109957 -51337
rect 110049 -51381 110057 -51337
rect 110149 -51381 110157 -51337
rect 110249 -51381 110257 -51337
rect 110349 -51381 110357 -51337
rect 110449 -51381 110457 -51337
rect 110549 -51381 110557 -51337
rect 110649 -51381 110657 -51337
rect 110749 -51381 110757 -51337
rect 110849 -51381 110857 -51337
rect 111349 -51381 111357 -51337
rect 111449 -51381 111457 -51337
rect 111549 -51381 111557 -51337
rect 111649 -51381 111657 -51337
rect 111749 -51381 111757 -51337
rect 111849 -51381 111857 -51337
rect 111949 -51381 111957 -51337
rect 112049 -51381 112057 -51337
rect 112149 -51381 112157 -51337
rect 112249 -51381 112257 -51337
rect 112349 -51381 112357 -51337
rect 112449 -51381 112457 -51337
rect 112549 -51381 112557 -51337
rect 112649 -51381 112657 -51337
rect 112749 -51381 112757 -51337
rect 112849 -51381 112857 -51337
rect 113349 -51381 113357 -51337
rect 113449 -51381 113457 -51337
rect 113549 -51381 113557 -51337
rect 113649 -51381 113657 -51337
rect 113749 -51381 113757 -51337
rect 113849 -51381 113857 -51337
rect 113949 -51381 113957 -51337
rect 114049 -51381 114057 -51337
rect 114149 -51381 114157 -51337
rect 114249 -51381 114257 -51337
rect 114349 -51381 114357 -51337
rect 114449 -51381 114457 -51337
rect 114549 -51381 114557 -51337
rect 114649 -51381 114657 -51337
rect 114749 -51381 114757 -51337
rect 114849 -51381 114857 -51337
rect 115349 -51381 115357 -51337
rect 115449 -51381 115457 -51337
rect 115549 -51381 115557 -51337
rect 115649 -51381 115657 -51337
rect 115749 -51381 115757 -51337
rect 115849 -51381 115857 -51337
rect 115949 -51381 115957 -51337
rect 116049 -51381 116057 -51337
rect 116149 -51381 116157 -51337
rect 116249 -51381 116257 -51337
rect 116349 -51381 116357 -51337
rect 116449 -51381 116457 -51337
rect 116549 -51381 116557 -51337
rect 116649 -51381 116657 -51337
rect 116749 -51381 116757 -51337
rect 116849 -51381 116857 -51337
rect 109305 -51437 109349 -51429
rect 109405 -51437 109449 -51429
rect 109505 -51437 109549 -51429
rect 109605 -51437 109649 -51429
rect 109705 -51437 109749 -51429
rect 109805 -51437 109849 -51429
rect 109905 -51437 109949 -51429
rect 110005 -51437 110049 -51429
rect 110105 -51437 110149 -51429
rect 110205 -51437 110249 -51429
rect 110305 -51437 110349 -51429
rect 110405 -51437 110449 -51429
rect 110505 -51437 110549 -51429
rect 110605 -51437 110649 -51429
rect 110705 -51437 110749 -51429
rect 110805 -51437 110849 -51429
rect 111305 -51437 111349 -51429
rect 111405 -51437 111449 -51429
rect 111505 -51437 111549 -51429
rect 111605 -51437 111649 -51429
rect 111705 -51437 111749 -51429
rect 111805 -51437 111849 -51429
rect 111905 -51437 111949 -51429
rect 112005 -51437 112049 -51429
rect 112105 -51437 112149 -51429
rect 112205 -51437 112249 -51429
rect 112305 -51437 112349 -51429
rect 112405 -51437 112449 -51429
rect 112505 -51437 112549 -51429
rect 112605 -51437 112649 -51429
rect 112705 -51437 112749 -51429
rect 112805 -51437 112849 -51429
rect 113305 -51437 113349 -51429
rect 113405 -51437 113449 -51429
rect 113505 -51437 113549 -51429
rect 113605 -51437 113649 -51429
rect 113705 -51437 113749 -51429
rect 113805 -51437 113849 -51429
rect 113905 -51437 113949 -51429
rect 114005 -51437 114049 -51429
rect 114105 -51437 114149 -51429
rect 114205 -51437 114249 -51429
rect 114305 -51437 114349 -51429
rect 114405 -51437 114449 -51429
rect 114505 -51437 114549 -51429
rect 114605 -51437 114649 -51429
rect 114705 -51437 114749 -51429
rect 114805 -51437 114849 -51429
rect 115305 -51437 115349 -51429
rect 115405 -51437 115449 -51429
rect 115505 -51437 115549 -51429
rect 115605 -51437 115649 -51429
rect 115705 -51437 115749 -51429
rect 115805 -51437 115849 -51429
rect 115905 -51437 115949 -51429
rect 116005 -51437 116049 -51429
rect 116105 -51437 116149 -51429
rect 116205 -51437 116249 -51429
rect 116305 -51437 116349 -51429
rect 116405 -51437 116449 -51429
rect 116505 -51437 116549 -51429
rect 116605 -51437 116649 -51429
rect 116705 -51437 116749 -51429
rect 116805 -51437 116849 -51429
rect 109349 -51481 109357 -51437
rect 109449 -51481 109457 -51437
rect 109549 -51481 109557 -51437
rect 109649 -51481 109657 -51437
rect 109749 -51481 109757 -51437
rect 109849 -51481 109857 -51437
rect 109949 -51481 109957 -51437
rect 110049 -51481 110057 -51437
rect 110149 -51481 110157 -51437
rect 110249 -51481 110257 -51437
rect 110349 -51481 110357 -51437
rect 110449 -51481 110457 -51437
rect 110549 -51481 110557 -51437
rect 110649 -51481 110657 -51437
rect 110749 -51481 110757 -51437
rect 110849 -51481 110857 -51437
rect 111349 -51481 111357 -51437
rect 111449 -51481 111457 -51437
rect 111549 -51481 111557 -51437
rect 111649 -51481 111657 -51437
rect 111749 -51481 111757 -51437
rect 111849 -51481 111857 -51437
rect 111949 -51481 111957 -51437
rect 112049 -51481 112057 -51437
rect 112149 -51481 112157 -51437
rect 112249 -51481 112257 -51437
rect 112349 -51481 112357 -51437
rect 112449 -51481 112457 -51437
rect 112549 -51481 112557 -51437
rect 112649 -51481 112657 -51437
rect 112749 -51481 112757 -51437
rect 112849 -51481 112857 -51437
rect 113349 -51481 113357 -51437
rect 113449 -51481 113457 -51437
rect 113549 -51481 113557 -51437
rect 113649 -51481 113657 -51437
rect 113749 -51481 113757 -51437
rect 113849 -51481 113857 -51437
rect 113949 -51481 113957 -51437
rect 114049 -51481 114057 -51437
rect 114149 -51481 114157 -51437
rect 114249 -51481 114257 -51437
rect 114349 -51481 114357 -51437
rect 114449 -51481 114457 -51437
rect 114549 -51481 114557 -51437
rect 114649 -51481 114657 -51437
rect 114749 -51481 114757 -51437
rect 114849 -51481 114857 -51437
rect 115349 -51481 115357 -51437
rect 115449 -51481 115457 -51437
rect 115549 -51481 115557 -51437
rect 115649 -51481 115657 -51437
rect 115749 -51481 115757 -51437
rect 115849 -51481 115857 -51437
rect 115949 -51481 115957 -51437
rect 116049 -51481 116057 -51437
rect 116149 -51481 116157 -51437
rect 116249 -51481 116257 -51437
rect 116349 -51481 116357 -51437
rect 116449 -51481 116457 -51437
rect 116549 -51481 116557 -51437
rect 116649 -51481 116657 -51437
rect 116749 -51481 116757 -51437
rect 116849 -51481 116857 -51437
rect 109305 -51537 109349 -51529
rect 109405 -51537 109449 -51529
rect 109505 -51537 109549 -51529
rect 109605 -51537 109649 -51529
rect 109705 -51537 109749 -51529
rect 109805 -51537 109849 -51529
rect 109905 -51537 109949 -51529
rect 110005 -51537 110049 -51529
rect 110105 -51537 110149 -51529
rect 110205 -51537 110249 -51529
rect 110305 -51537 110349 -51529
rect 110405 -51537 110449 -51529
rect 110505 -51537 110549 -51529
rect 110605 -51537 110649 -51529
rect 110705 -51537 110749 -51529
rect 110805 -51537 110849 -51529
rect 111305 -51537 111349 -51529
rect 111405 -51537 111449 -51529
rect 111505 -51537 111549 -51529
rect 111605 -51537 111649 -51529
rect 111705 -51537 111749 -51529
rect 111805 -51537 111849 -51529
rect 111905 -51537 111949 -51529
rect 112005 -51537 112049 -51529
rect 112105 -51537 112149 -51529
rect 112205 -51537 112249 -51529
rect 112305 -51537 112349 -51529
rect 112405 -51537 112449 -51529
rect 112505 -51537 112549 -51529
rect 112605 -51537 112649 -51529
rect 112705 -51537 112749 -51529
rect 112805 -51537 112849 -51529
rect 113305 -51537 113349 -51529
rect 113405 -51537 113449 -51529
rect 113505 -51537 113549 -51529
rect 113605 -51537 113649 -51529
rect 113705 -51537 113749 -51529
rect 113805 -51537 113849 -51529
rect 113905 -51537 113949 -51529
rect 114005 -51537 114049 -51529
rect 114105 -51537 114149 -51529
rect 114205 -51537 114249 -51529
rect 114305 -51537 114349 -51529
rect 114405 -51537 114449 -51529
rect 114505 -51537 114549 -51529
rect 114605 -51537 114649 -51529
rect 114705 -51537 114749 -51529
rect 114805 -51537 114849 -51529
rect 115305 -51537 115349 -51529
rect 115405 -51537 115449 -51529
rect 115505 -51537 115549 -51529
rect 115605 -51537 115649 -51529
rect 115705 -51537 115749 -51529
rect 115805 -51537 115849 -51529
rect 115905 -51537 115949 -51529
rect 116005 -51537 116049 -51529
rect 116105 -51537 116149 -51529
rect 116205 -51537 116249 -51529
rect 116305 -51537 116349 -51529
rect 116405 -51537 116449 -51529
rect 116505 -51537 116549 -51529
rect 116605 -51537 116649 -51529
rect 116705 -51537 116749 -51529
rect 116805 -51537 116849 -51529
rect 109349 -51581 109357 -51537
rect 109449 -51581 109457 -51537
rect 109549 -51581 109557 -51537
rect 109649 -51581 109657 -51537
rect 109749 -51581 109757 -51537
rect 109849 -51581 109857 -51537
rect 109949 -51581 109957 -51537
rect 110049 -51581 110057 -51537
rect 110149 -51581 110157 -51537
rect 110249 -51581 110257 -51537
rect 110349 -51581 110357 -51537
rect 110449 -51581 110457 -51537
rect 110549 -51581 110557 -51537
rect 110649 -51581 110657 -51537
rect 110749 -51581 110757 -51537
rect 110849 -51581 110857 -51537
rect 111349 -51581 111357 -51537
rect 111449 -51581 111457 -51537
rect 111549 -51581 111557 -51537
rect 111649 -51581 111657 -51537
rect 111749 -51581 111757 -51537
rect 111849 -51581 111857 -51537
rect 111949 -51581 111957 -51537
rect 112049 -51581 112057 -51537
rect 112149 -51581 112157 -51537
rect 112249 -51581 112257 -51537
rect 112349 -51581 112357 -51537
rect 112449 -51581 112457 -51537
rect 112549 -51581 112557 -51537
rect 112649 -51581 112657 -51537
rect 112749 -51581 112757 -51537
rect 112849 -51581 112857 -51537
rect 113349 -51581 113357 -51537
rect 113449 -51581 113457 -51537
rect 113549 -51581 113557 -51537
rect 113649 -51581 113657 -51537
rect 113749 -51581 113757 -51537
rect 113849 -51581 113857 -51537
rect 113949 -51581 113957 -51537
rect 114049 -51581 114057 -51537
rect 114149 -51581 114157 -51537
rect 114249 -51581 114257 -51537
rect 114349 -51581 114357 -51537
rect 114449 -51581 114457 -51537
rect 114549 -51581 114557 -51537
rect 114649 -51581 114657 -51537
rect 114749 -51581 114757 -51537
rect 114849 -51581 114857 -51537
rect 115349 -51581 115357 -51537
rect 115449 -51581 115457 -51537
rect 115549 -51581 115557 -51537
rect 115649 -51581 115657 -51537
rect 115749 -51581 115757 -51537
rect 115849 -51581 115857 -51537
rect 115949 -51581 115957 -51537
rect 116049 -51581 116057 -51537
rect 116149 -51581 116157 -51537
rect 116249 -51581 116257 -51537
rect 116349 -51581 116357 -51537
rect 116449 -51581 116457 -51537
rect 116549 -51581 116557 -51537
rect 116649 -51581 116657 -51537
rect 116749 -51581 116757 -51537
rect 116849 -51581 116857 -51537
rect 109305 -51637 109349 -51629
rect 109405 -51637 109449 -51629
rect 109505 -51637 109549 -51629
rect 109605 -51637 109649 -51629
rect 109705 -51637 109749 -51629
rect 109805 -51637 109849 -51629
rect 109905 -51637 109949 -51629
rect 110005 -51637 110049 -51629
rect 110105 -51637 110149 -51629
rect 110205 -51637 110249 -51629
rect 110305 -51637 110349 -51629
rect 110405 -51637 110449 -51629
rect 110505 -51637 110549 -51629
rect 110605 -51637 110649 -51629
rect 110705 -51637 110749 -51629
rect 110805 -51637 110849 -51629
rect 111305 -51637 111349 -51629
rect 111405 -51637 111449 -51629
rect 111505 -51637 111549 -51629
rect 111605 -51637 111649 -51629
rect 111705 -51637 111749 -51629
rect 111805 -51637 111849 -51629
rect 111905 -51637 111949 -51629
rect 112005 -51637 112049 -51629
rect 112105 -51637 112149 -51629
rect 112205 -51637 112249 -51629
rect 112305 -51637 112349 -51629
rect 112405 -51637 112449 -51629
rect 112505 -51637 112549 -51629
rect 112605 -51637 112649 -51629
rect 112705 -51637 112749 -51629
rect 112805 -51637 112849 -51629
rect 113305 -51637 113349 -51629
rect 113405 -51637 113449 -51629
rect 113505 -51637 113549 -51629
rect 113605 -51637 113649 -51629
rect 113705 -51637 113749 -51629
rect 113805 -51637 113849 -51629
rect 113905 -51637 113949 -51629
rect 114005 -51637 114049 -51629
rect 114105 -51637 114149 -51629
rect 114205 -51637 114249 -51629
rect 114305 -51637 114349 -51629
rect 114405 -51637 114449 -51629
rect 114505 -51637 114549 -51629
rect 114605 -51637 114649 -51629
rect 114705 -51637 114749 -51629
rect 114805 -51637 114849 -51629
rect 115305 -51637 115349 -51629
rect 115405 -51637 115449 -51629
rect 115505 -51637 115549 -51629
rect 115605 -51637 115649 -51629
rect 115705 -51637 115749 -51629
rect 115805 -51637 115849 -51629
rect 115905 -51637 115949 -51629
rect 116005 -51637 116049 -51629
rect 116105 -51637 116149 -51629
rect 116205 -51637 116249 -51629
rect 116305 -51637 116349 -51629
rect 116405 -51637 116449 -51629
rect 116505 -51637 116549 -51629
rect 116605 -51637 116649 -51629
rect 116705 -51637 116749 -51629
rect 116805 -51637 116849 -51629
rect 109349 -51681 109357 -51637
rect 109449 -51681 109457 -51637
rect 109549 -51681 109557 -51637
rect 109649 -51681 109657 -51637
rect 109749 -51681 109757 -51637
rect 109849 -51681 109857 -51637
rect 109949 -51681 109957 -51637
rect 110049 -51681 110057 -51637
rect 110149 -51681 110157 -51637
rect 110249 -51681 110257 -51637
rect 110349 -51681 110357 -51637
rect 110449 -51681 110457 -51637
rect 110549 -51681 110557 -51637
rect 110649 -51681 110657 -51637
rect 110749 -51681 110757 -51637
rect 110849 -51681 110857 -51637
rect 111349 -51681 111357 -51637
rect 111449 -51681 111457 -51637
rect 111549 -51681 111557 -51637
rect 111649 -51681 111657 -51637
rect 111749 -51681 111757 -51637
rect 111849 -51681 111857 -51637
rect 111949 -51681 111957 -51637
rect 112049 -51681 112057 -51637
rect 112149 -51681 112157 -51637
rect 112249 -51681 112257 -51637
rect 112349 -51681 112357 -51637
rect 112449 -51681 112457 -51637
rect 112549 -51681 112557 -51637
rect 112649 -51681 112657 -51637
rect 112749 -51681 112757 -51637
rect 112849 -51681 112857 -51637
rect 113349 -51681 113357 -51637
rect 113449 -51681 113457 -51637
rect 113549 -51681 113557 -51637
rect 113649 -51681 113657 -51637
rect 113749 -51681 113757 -51637
rect 113849 -51681 113857 -51637
rect 113949 -51681 113957 -51637
rect 114049 -51681 114057 -51637
rect 114149 -51681 114157 -51637
rect 114249 -51681 114257 -51637
rect 114349 -51681 114357 -51637
rect 114449 -51681 114457 -51637
rect 114549 -51681 114557 -51637
rect 114649 -51681 114657 -51637
rect 114749 -51681 114757 -51637
rect 114849 -51681 114857 -51637
rect 115349 -51681 115357 -51637
rect 115449 -51681 115457 -51637
rect 115549 -51681 115557 -51637
rect 115649 -51681 115657 -51637
rect 115749 -51681 115757 -51637
rect 115849 -51681 115857 -51637
rect 115949 -51681 115957 -51637
rect 116049 -51681 116057 -51637
rect 116149 -51681 116157 -51637
rect 116249 -51681 116257 -51637
rect 116349 -51681 116357 -51637
rect 116449 -51681 116457 -51637
rect 116549 -51681 116557 -51637
rect 116649 -51681 116657 -51637
rect 116749 -51681 116757 -51637
rect 116849 -51681 116857 -51637
rect 109305 -51737 109349 -51729
rect 109405 -51737 109449 -51729
rect 109505 -51737 109549 -51729
rect 109605 -51737 109649 -51729
rect 109705 -51737 109749 -51729
rect 109805 -51737 109849 -51729
rect 109905 -51737 109949 -51729
rect 110005 -51737 110049 -51729
rect 110105 -51737 110149 -51729
rect 110205 -51737 110249 -51729
rect 110305 -51737 110349 -51729
rect 110405 -51737 110449 -51729
rect 110505 -51737 110549 -51729
rect 110605 -51737 110649 -51729
rect 110705 -51737 110749 -51729
rect 110805 -51737 110849 -51729
rect 111305 -51737 111349 -51729
rect 111405 -51737 111449 -51729
rect 111505 -51737 111549 -51729
rect 111605 -51737 111649 -51729
rect 111705 -51737 111749 -51729
rect 111805 -51737 111849 -51729
rect 111905 -51737 111949 -51729
rect 112005 -51737 112049 -51729
rect 112105 -51737 112149 -51729
rect 112205 -51737 112249 -51729
rect 112305 -51737 112349 -51729
rect 112405 -51737 112449 -51729
rect 112505 -51737 112549 -51729
rect 112605 -51737 112649 -51729
rect 112705 -51737 112749 -51729
rect 112805 -51737 112849 -51729
rect 113305 -51737 113349 -51729
rect 113405 -51737 113449 -51729
rect 113505 -51737 113549 -51729
rect 113605 -51737 113649 -51729
rect 113705 -51737 113749 -51729
rect 113805 -51737 113849 -51729
rect 113905 -51737 113949 -51729
rect 114005 -51737 114049 -51729
rect 114105 -51737 114149 -51729
rect 114205 -51737 114249 -51729
rect 114305 -51737 114349 -51729
rect 114405 -51737 114449 -51729
rect 114505 -51737 114549 -51729
rect 114605 -51737 114649 -51729
rect 114705 -51737 114749 -51729
rect 114805 -51737 114849 -51729
rect 115305 -51737 115349 -51729
rect 115405 -51737 115449 -51729
rect 115505 -51737 115549 -51729
rect 115605 -51737 115649 -51729
rect 115705 -51737 115749 -51729
rect 115805 -51737 115849 -51729
rect 115905 -51737 115949 -51729
rect 116005 -51737 116049 -51729
rect 116105 -51737 116149 -51729
rect 116205 -51737 116249 -51729
rect 116305 -51737 116349 -51729
rect 116405 -51737 116449 -51729
rect 116505 -51737 116549 -51729
rect 116605 -51737 116649 -51729
rect 116705 -51737 116749 -51729
rect 116805 -51737 116849 -51729
rect 109349 -51781 109357 -51737
rect 109449 -51781 109457 -51737
rect 109549 -51781 109557 -51737
rect 109649 -51781 109657 -51737
rect 109749 -51781 109757 -51737
rect 109849 -51781 109857 -51737
rect 109949 -51781 109957 -51737
rect 110049 -51781 110057 -51737
rect 110149 -51781 110157 -51737
rect 110249 -51781 110257 -51737
rect 110349 -51781 110357 -51737
rect 110449 -51781 110457 -51737
rect 110549 -51781 110557 -51737
rect 110649 -51781 110657 -51737
rect 110749 -51781 110757 -51737
rect 110849 -51781 110857 -51737
rect 111349 -51781 111357 -51737
rect 111449 -51781 111457 -51737
rect 111549 -51781 111557 -51737
rect 111649 -51781 111657 -51737
rect 111749 -51781 111757 -51737
rect 111849 -51781 111857 -51737
rect 111949 -51781 111957 -51737
rect 112049 -51781 112057 -51737
rect 112149 -51781 112157 -51737
rect 112249 -51781 112257 -51737
rect 112349 -51781 112357 -51737
rect 112449 -51781 112457 -51737
rect 112549 -51781 112557 -51737
rect 112649 -51781 112657 -51737
rect 112749 -51781 112757 -51737
rect 112849 -51781 112857 -51737
rect 113349 -51781 113357 -51737
rect 113449 -51781 113457 -51737
rect 113549 -51781 113557 -51737
rect 113649 -51781 113657 -51737
rect 113749 -51781 113757 -51737
rect 113849 -51781 113857 -51737
rect 113949 -51781 113957 -51737
rect 114049 -51781 114057 -51737
rect 114149 -51781 114157 -51737
rect 114249 -51781 114257 -51737
rect 114349 -51781 114357 -51737
rect 114449 -51781 114457 -51737
rect 114549 -51781 114557 -51737
rect 114649 -51781 114657 -51737
rect 114749 -51781 114757 -51737
rect 114849 -51781 114857 -51737
rect 115349 -51781 115357 -51737
rect 115449 -51781 115457 -51737
rect 115549 -51781 115557 -51737
rect 115649 -51781 115657 -51737
rect 115749 -51781 115757 -51737
rect 115849 -51781 115857 -51737
rect 115949 -51781 115957 -51737
rect 116049 -51781 116057 -51737
rect 116149 -51781 116157 -51737
rect 116249 -51781 116257 -51737
rect 116349 -51781 116357 -51737
rect 116449 -51781 116457 -51737
rect 116549 -51781 116557 -51737
rect 116649 -51781 116657 -51737
rect 116749 -51781 116757 -51737
rect 116849 -51781 116857 -51737
rect 109305 -51837 109349 -51829
rect 109405 -51837 109449 -51829
rect 109505 -51837 109549 -51829
rect 109605 -51837 109649 -51829
rect 109705 -51837 109749 -51829
rect 109805 -51837 109849 -51829
rect 109905 -51837 109949 -51829
rect 110005 -51837 110049 -51829
rect 110105 -51837 110149 -51829
rect 110205 -51837 110249 -51829
rect 110305 -51837 110349 -51829
rect 110405 -51837 110449 -51829
rect 110505 -51837 110549 -51829
rect 110605 -51837 110649 -51829
rect 110705 -51837 110749 -51829
rect 110805 -51837 110849 -51829
rect 111305 -51837 111349 -51829
rect 111405 -51837 111449 -51829
rect 111505 -51837 111549 -51829
rect 111605 -51837 111649 -51829
rect 111705 -51837 111749 -51829
rect 111805 -51837 111849 -51829
rect 111905 -51837 111949 -51829
rect 112005 -51837 112049 -51829
rect 112105 -51837 112149 -51829
rect 112205 -51837 112249 -51829
rect 112305 -51837 112349 -51829
rect 112405 -51837 112449 -51829
rect 112505 -51837 112549 -51829
rect 112605 -51837 112649 -51829
rect 112705 -51837 112749 -51829
rect 112805 -51837 112849 -51829
rect 113305 -51837 113349 -51829
rect 113405 -51837 113449 -51829
rect 113505 -51837 113549 -51829
rect 113605 -51837 113649 -51829
rect 113705 -51837 113749 -51829
rect 113805 -51837 113849 -51829
rect 113905 -51837 113949 -51829
rect 114005 -51837 114049 -51829
rect 114105 -51837 114149 -51829
rect 114205 -51837 114249 -51829
rect 114305 -51837 114349 -51829
rect 114405 -51837 114449 -51829
rect 114505 -51837 114549 -51829
rect 114605 -51837 114649 -51829
rect 114705 -51837 114749 -51829
rect 114805 -51837 114849 -51829
rect 115305 -51837 115349 -51829
rect 115405 -51837 115449 -51829
rect 115505 -51837 115549 -51829
rect 115605 -51837 115649 -51829
rect 115705 -51837 115749 -51829
rect 115805 -51837 115849 -51829
rect 115905 -51837 115949 -51829
rect 116005 -51837 116049 -51829
rect 116105 -51837 116149 -51829
rect 116205 -51837 116249 -51829
rect 116305 -51837 116349 -51829
rect 116405 -51837 116449 -51829
rect 116505 -51837 116549 -51829
rect 116605 -51837 116649 -51829
rect 116705 -51837 116749 -51829
rect 116805 -51837 116849 -51829
rect 109349 -51881 109357 -51837
rect 109449 -51881 109457 -51837
rect 109549 -51881 109557 -51837
rect 109649 -51881 109657 -51837
rect 109749 -51881 109757 -51837
rect 109849 -51881 109857 -51837
rect 109949 -51881 109957 -51837
rect 110049 -51881 110057 -51837
rect 110149 -51881 110157 -51837
rect 110249 -51881 110257 -51837
rect 110349 -51881 110357 -51837
rect 110449 -51881 110457 -51837
rect 110549 -51881 110557 -51837
rect 110649 -51881 110657 -51837
rect 110749 -51881 110757 -51837
rect 110849 -51881 110857 -51837
rect 111349 -51881 111357 -51837
rect 111449 -51881 111457 -51837
rect 111549 -51881 111557 -51837
rect 111649 -51881 111657 -51837
rect 111749 -51881 111757 -51837
rect 111849 -51881 111857 -51837
rect 111949 -51881 111957 -51837
rect 112049 -51881 112057 -51837
rect 112149 -51881 112157 -51837
rect 112249 -51881 112257 -51837
rect 112349 -51881 112357 -51837
rect 112449 -51881 112457 -51837
rect 112549 -51881 112557 -51837
rect 112649 -51881 112657 -51837
rect 112749 -51881 112757 -51837
rect 112849 -51881 112857 -51837
rect 113349 -51881 113357 -51837
rect 113449 -51881 113457 -51837
rect 113549 -51881 113557 -51837
rect 113649 -51881 113657 -51837
rect 113749 -51881 113757 -51837
rect 113849 -51881 113857 -51837
rect 113949 -51881 113957 -51837
rect 114049 -51881 114057 -51837
rect 114149 -51881 114157 -51837
rect 114249 -51881 114257 -51837
rect 114349 -51881 114357 -51837
rect 114449 -51881 114457 -51837
rect 114549 -51881 114557 -51837
rect 114649 -51881 114657 -51837
rect 114749 -51881 114757 -51837
rect 114849 -51881 114857 -51837
rect 115349 -51881 115357 -51837
rect 115449 -51881 115457 -51837
rect 115549 -51881 115557 -51837
rect 115649 -51881 115657 -51837
rect 115749 -51881 115757 -51837
rect 115849 -51881 115857 -51837
rect 115949 -51881 115957 -51837
rect 116049 -51881 116057 -51837
rect 116149 -51881 116157 -51837
rect 116249 -51881 116257 -51837
rect 116349 -51881 116357 -51837
rect 116449 -51881 116457 -51837
rect 116549 -51881 116557 -51837
rect 116649 -51881 116657 -51837
rect 116749 -51881 116757 -51837
rect 116849 -51881 116857 -51837
rect 109305 -51937 109349 -51929
rect 109405 -51937 109449 -51929
rect 109505 -51937 109549 -51929
rect 109605 -51937 109649 -51929
rect 109705 -51937 109749 -51929
rect 109805 -51937 109849 -51929
rect 109905 -51937 109949 -51929
rect 110005 -51937 110049 -51929
rect 110105 -51937 110149 -51929
rect 110205 -51937 110249 -51929
rect 110305 -51937 110349 -51929
rect 110405 -51937 110449 -51929
rect 110505 -51937 110549 -51929
rect 110605 -51937 110649 -51929
rect 110705 -51937 110749 -51929
rect 110805 -51937 110849 -51929
rect 111305 -51937 111349 -51929
rect 111405 -51937 111449 -51929
rect 111505 -51937 111549 -51929
rect 111605 -51937 111649 -51929
rect 111705 -51937 111749 -51929
rect 111805 -51937 111849 -51929
rect 111905 -51937 111949 -51929
rect 112005 -51937 112049 -51929
rect 112105 -51937 112149 -51929
rect 112205 -51937 112249 -51929
rect 112305 -51937 112349 -51929
rect 112405 -51937 112449 -51929
rect 112505 -51937 112549 -51929
rect 112605 -51937 112649 -51929
rect 112705 -51937 112749 -51929
rect 112805 -51937 112849 -51929
rect 113305 -51937 113349 -51929
rect 113405 -51937 113449 -51929
rect 113505 -51937 113549 -51929
rect 113605 -51937 113649 -51929
rect 113705 -51937 113749 -51929
rect 113805 -51937 113849 -51929
rect 113905 -51937 113949 -51929
rect 114005 -51937 114049 -51929
rect 114105 -51937 114149 -51929
rect 114205 -51937 114249 -51929
rect 114305 -51937 114349 -51929
rect 114405 -51937 114449 -51929
rect 114505 -51937 114549 -51929
rect 114605 -51937 114649 -51929
rect 114705 -51937 114749 -51929
rect 114805 -51937 114849 -51929
rect 115305 -51937 115349 -51929
rect 115405 -51937 115449 -51929
rect 115505 -51937 115549 -51929
rect 115605 -51937 115649 -51929
rect 115705 -51937 115749 -51929
rect 115805 -51937 115849 -51929
rect 115905 -51937 115949 -51929
rect 116005 -51937 116049 -51929
rect 116105 -51937 116149 -51929
rect 116205 -51937 116249 -51929
rect 116305 -51937 116349 -51929
rect 116405 -51937 116449 -51929
rect 116505 -51937 116549 -51929
rect 116605 -51937 116649 -51929
rect 116705 -51937 116749 -51929
rect 116805 -51937 116849 -51929
rect 109349 -51981 109357 -51937
rect 109449 -51981 109457 -51937
rect 109549 -51981 109557 -51937
rect 109649 -51981 109657 -51937
rect 109749 -51981 109757 -51937
rect 109849 -51981 109857 -51937
rect 109949 -51981 109957 -51937
rect 110049 -51981 110057 -51937
rect 110149 -51981 110157 -51937
rect 110249 -51981 110257 -51937
rect 110349 -51981 110357 -51937
rect 110449 -51981 110457 -51937
rect 110549 -51981 110557 -51937
rect 110649 -51981 110657 -51937
rect 110749 -51981 110757 -51937
rect 110849 -51981 110857 -51937
rect 111349 -51981 111357 -51937
rect 111449 -51981 111457 -51937
rect 111549 -51981 111557 -51937
rect 111649 -51981 111657 -51937
rect 111749 -51981 111757 -51937
rect 111849 -51981 111857 -51937
rect 111949 -51981 111957 -51937
rect 112049 -51981 112057 -51937
rect 112149 -51981 112157 -51937
rect 112249 -51981 112257 -51937
rect 112349 -51981 112357 -51937
rect 112449 -51981 112457 -51937
rect 112549 -51981 112557 -51937
rect 112649 -51981 112657 -51937
rect 112749 -51981 112757 -51937
rect 112849 -51981 112857 -51937
rect 113349 -51981 113357 -51937
rect 113449 -51981 113457 -51937
rect 113549 -51981 113557 -51937
rect 113649 -51981 113657 -51937
rect 113749 -51981 113757 -51937
rect 113849 -51981 113857 -51937
rect 113949 -51981 113957 -51937
rect 114049 -51981 114057 -51937
rect 114149 -51981 114157 -51937
rect 114249 -51981 114257 -51937
rect 114349 -51981 114357 -51937
rect 114449 -51981 114457 -51937
rect 114549 -51981 114557 -51937
rect 114649 -51981 114657 -51937
rect 114749 -51981 114757 -51937
rect 114849 -51981 114857 -51937
rect 115349 -51981 115357 -51937
rect 115449 -51981 115457 -51937
rect 115549 -51981 115557 -51937
rect 115649 -51981 115657 -51937
rect 115749 -51981 115757 -51937
rect 115849 -51981 115857 -51937
rect 115949 -51981 115957 -51937
rect 116049 -51981 116057 -51937
rect 116149 -51981 116157 -51937
rect 116249 -51981 116257 -51937
rect 116349 -51981 116357 -51937
rect 116449 -51981 116457 -51937
rect 116549 -51981 116557 -51937
rect 116649 -51981 116657 -51937
rect 116749 -51981 116757 -51937
rect 116849 -51981 116857 -51937
rect 109305 -52037 109349 -52029
rect 109405 -52037 109449 -52029
rect 109505 -52037 109549 -52029
rect 109605 -52037 109649 -52029
rect 109705 -52037 109749 -52029
rect 109805 -52037 109849 -52029
rect 109905 -52037 109949 -52029
rect 110005 -52037 110049 -52029
rect 110105 -52037 110149 -52029
rect 110205 -52037 110249 -52029
rect 110305 -52037 110349 -52029
rect 110405 -52037 110449 -52029
rect 110505 -52037 110549 -52029
rect 110605 -52037 110649 -52029
rect 110705 -52037 110749 -52029
rect 110805 -52037 110849 -52029
rect 111305 -52037 111349 -52029
rect 111405 -52037 111449 -52029
rect 111505 -52037 111549 -52029
rect 111605 -52037 111649 -52029
rect 111705 -52037 111749 -52029
rect 111805 -52037 111849 -52029
rect 111905 -52037 111949 -52029
rect 112005 -52037 112049 -52029
rect 112105 -52037 112149 -52029
rect 112205 -52037 112249 -52029
rect 112305 -52037 112349 -52029
rect 112405 -52037 112449 -52029
rect 112505 -52037 112549 -52029
rect 112605 -52037 112649 -52029
rect 112705 -52037 112749 -52029
rect 112805 -52037 112849 -52029
rect 113305 -52037 113349 -52029
rect 113405 -52037 113449 -52029
rect 113505 -52037 113549 -52029
rect 113605 -52037 113649 -52029
rect 113705 -52037 113749 -52029
rect 113805 -52037 113849 -52029
rect 113905 -52037 113949 -52029
rect 114005 -52037 114049 -52029
rect 114105 -52037 114149 -52029
rect 114205 -52037 114249 -52029
rect 114305 -52037 114349 -52029
rect 114405 -52037 114449 -52029
rect 114505 -52037 114549 -52029
rect 114605 -52037 114649 -52029
rect 114705 -52037 114749 -52029
rect 114805 -52037 114849 -52029
rect 115305 -52037 115349 -52029
rect 115405 -52037 115449 -52029
rect 115505 -52037 115549 -52029
rect 115605 -52037 115649 -52029
rect 115705 -52037 115749 -52029
rect 115805 -52037 115849 -52029
rect 115905 -52037 115949 -52029
rect 116005 -52037 116049 -52029
rect 116105 -52037 116149 -52029
rect 116205 -52037 116249 -52029
rect 116305 -52037 116349 -52029
rect 116405 -52037 116449 -52029
rect 116505 -52037 116549 -52029
rect 116605 -52037 116649 -52029
rect 116705 -52037 116749 -52029
rect 116805 -52037 116849 -52029
rect 109349 -52081 109357 -52037
rect 109449 -52081 109457 -52037
rect 109549 -52081 109557 -52037
rect 109649 -52081 109657 -52037
rect 109749 -52081 109757 -52037
rect 109849 -52081 109857 -52037
rect 109949 -52081 109957 -52037
rect 110049 -52081 110057 -52037
rect 110149 -52081 110157 -52037
rect 110249 -52081 110257 -52037
rect 110349 -52081 110357 -52037
rect 110449 -52081 110457 -52037
rect 110549 -52081 110557 -52037
rect 110649 -52081 110657 -52037
rect 110749 -52081 110757 -52037
rect 110849 -52081 110857 -52037
rect 111349 -52081 111357 -52037
rect 111449 -52081 111457 -52037
rect 111549 -52081 111557 -52037
rect 111649 -52081 111657 -52037
rect 111749 -52081 111757 -52037
rect 111849 -52081 111857 -52037
rect 111949 -52081 111957 -52037
rect 112049 -52081 112057 -52037
rect 112149 -52081 112157 -52037
rect 112249 -52081 112257 -52037
rect 112349 -52081 112357 -52037
rect 112449 -52081 112457 -52037
rect 112549 -52081 112557 -52037
rect 112649 -52081 112657 -52037
rect 112749 -52081 112757 -52037
rect 112849 -52081 112857 -52037
rect 113349 -52081 113357 -52037
rect 113449 -52081 113457 -52037
rect 113549 -52081 113557 -52037
rect 113649 -52081 113657 -52037
rect 113749 -52081 113757 -52037
rect 113849 -52081 113857 -52037
rect 113949 -52081 113957 -52037
rect 114049 -52081 114057 -52037
rect 114149 -52081 114157 -52037
rect 114249 -52081 114257 -52037
rect 114349 -52081 114357 -52037
rect 114449 -52081 114457 -52037
rect 114549 -52081 114557 -52037
rect 114649 -52081 114657 -52037
rect 114749 -52081 114757 -52037
rect 114849 -52081 114857 -52037
rect 115349 -52081 115357 -52037
rect 115449 -52081 115457 -52037
rect 115549 -52081 115557 -52037
rect 115649 -52081 115657 -52037
rect 115749 -52081 115757 -52037
rect 115849 -52081 115857 -52037
rect 115949 -52081 115957 -52037
rect 116049 -52081 116057 -52037
rect 116149 -52081 116157 -52037
rect 116249 -52081 116257 -52037
rect 116349 -52081 116357 -52037
rect 116449 -52081 116457 -52037
rect 116549 -52081 116557 -52037
rect 116649 -52081 116657 -52037
rect 116749 -52081 116757 -52037
rect 116849 -52081 116857 -52037
rect 109305 -52137 109349 -52129
rect 109405 -52137 109449 -52129
rect 109505 -52137 109549 -52129
rect 109605 -52137 109649 -52129
rect 109705 -52137 109749 -52129
rect 109805 -52137 109849 -52129
rect 109905 -52137 109949 -52129
rect 110005 -52137 110049 -52129
rect 110105 -52137 110149 -52129
rect 110205 -52137 110249 -52129
rect 110305 -52137 110349 -52129
rect 110405 -52137 110449 -52129
rect 110505 -52137 110549 -52129
rect 110605 -52137 110649 -52129
rect 110705 -52137 110749 -52129
rect 110805 -52137 110849 -52129
rect 111305 -52137 111349 -52129
rect 111405 -52137 111449 -52129
rect 111505 -52137 111549 -52129
rect 111605 -52137 111649 -52129
rect 111705 -52137 111749 -52129
rect 111805 -52137 111849 -52129
rect 111905 -52137 111949 -52129
rect 112005 -52137 112049 -52129
rect 112105 -52137 112149 -52129
rect 112205 -52137 112249 -52129
rect 112305 -52137 112349 -52129
rect 112405 -52137 112449 -52129
rect 112505 -52137 112549 -52129
rect 112605 -52137 112649 -52129
rect 112705 -52137 112749 -52129
rect 112805 -52137 112849 -52129
rect 113305 -52137 113349 -52129
rect 113405 -52137 113449 -52129
rect 113505 -52137 113549 -52129
rect 113605 -52137 113649 -52129
rect 113705 -52137 113749 -52129
rect 113805 -52137 113849 -52129
rect 113905 -52137 113949 -52129
rect 114005 -52137 114049 -52129
rect 114105 -52137 114149 -52129
rect 114205 -52137 114249 -52129
rect 114305 -52137 114349 -52129
rect 114405 -52137 114449 -52129
rect 114505 -52137 114549 -52129
rect 114605 -52137 114649 -52129
rect 114705 -52137 114749 -52129
rect 114805 -52137 114849 -52129
rect 115305 -52137 115349 -52129
rect 115405 -52137 115449 -52129
rect 115505 -52137 115549 -52129
rect 115605 -52137 115649 -52129
rect 115705 -52137 115749 -52129
rect 115805 -52137 115849 -52129
rect 115905 -52137 115949 -52129
rect 116005 -52137 116049 -52129
rect 116105 -52137 116149 -52129
rect 116205 -52137 116249 -52129
rect 116305 -52137 116349 -52129
rect 116405 -52137 116449 -52129
rect 116505 -52137 116549 -52129
rect 116605 -52137 116649 -52129
rect 116705 -52137 116749 -52129
rect 116805 -52137 116849 -52129
rect 109349 -52181 109357 -52137
rect 109449 -52181 109457 -52137
rect 109549 -52181 109557 -52137
rect 109649 -52181 109657 -52137
rect 109749 -52181 109757 -52137
rect 109849 -52181 109857 -52137
rect 109949 -52181 109957 -52137
rect 110049 -52181 110057 -52137
rect 110149 -52181 110157 -52137
rect 110249 -52181 110257 -52137
rect 110349 -52181 110357 -52137
rect 110449 -52181 110457 -52137
rect 110549 -52181 110557 -52137
rect 110649 -52181 110657 -52137
rect 110749 -52181 110757 -52137
rect 110849 -52181 110857 -52137
rect 111349 -52181 111357 -52137
rect 111449 -52181 111457 -52137
rect 111549 -52181 111557 -52137
rect 111649 -52181 111657 -52137
rect 111749 -52181 111757 -52137
rect 111849 -52181 111857 -52137
rect 111949 -52181 111957 -52137
rect 112049 -52181 112057 -52137
rect 112149 -52181 112157 -52137
rect 112249 -52181 112257 -52137
rect 112349 -52181 112357 -52137
rect 112449 -52181 112457 -52137
rect 112549 -52181 112557 -52137
rect 112649 -52181 112657 -52137
rect 112749 -52181 112757 -52137
rect 112849 -52181 112857 -52137
rect 113349 -52181 113357 -52137
rect 113449 -52181 113457 -52137
rect 113549 -52181 113557 -52137
rect 113649 -52181 113657 -52137
rect 113749 -52181 113757 -52137
rect 113849 -52181 113857 -52137
rect 113949 -52181 113957 -52137
rect 114049 -52181 114057 -52137
rect 114149 -52181 114157 -52137
rect 114249 -52181 114257 -52137
rect 114349 -52181 114357 -52137
rect 114449 -52181 114457 -52137
rect 114549 -52181 114557 -52137
rect 114649 -52181 114657 -52137
rect 114749 -52181 114757 -52137
rect 114849 -52181 114857 -52137
rect 115349 -52181 115357 -52137
rect 115449 -52181 115457 -52137
rect 115549 -52181 115557 -52137
rect 115649 -52181 115657 -52137
rect 115749 -52181 115757 -52137
rect 115849 -52181 115857 -52137
rect 115949 -52181 115957 -52137
rect 116049 -52181 116057 -52137
rect 116149 -52181 116157 -52137
rect 116249 -52181 116257 -52137
rect 116349 -52181 116357 -52137
rect 116449 -52181 116457 -52137
rect 116549 -52181 116557 -52137
rect 116649 -52181 116657 -52137
rect 116749 -52181 116757 -52137
rect 116849 -52181 116857 -52137
rect 109305 -52237 109349 -52229
rect 109405 -52237 109449 -52229
rect 109505 -52237 109549 -52229
rect 109605 -52237 109649 -52229
rect 109705 -52237 109749 -52229
rect 109805 -52237 109849 -52229
rect 109905 -52237 109949 -52229
rect 110005 -52237 110049 -52229
rect 110105 -52237 110149 -52229
rect 110205 -52237 110249 -52229
rect 110305 -52237 110349 -52229
rect 110405 -52237 110449 -52229
rect 110505 -52237 110549 -52229
rect 110605 -52237 110649 -52229
rect 110705 -52237 110749 -52229
rect 110805 -52237 110849 -52229
rect 111305 -52237 111349 -52229
rect 111405 -52237 111449 -52229
rect 111505 -52237 111549 -52229
rect 111605 -52237 111649 -52229
rect 111705 -52237 111749 -52229
rect 111805 -52237 111849 -52229
rect 111905 -52237 111949 -52229
rect 112005 -52237 112049 -52229
rect 112105 -52237 112149 -52229
rect 112205 -52237 112249 -52229
rect 112305 -52237 112349 -52229
rect 112405 -52237 112449 -52229
rect 112505 -52237 112549 -52229
rect 112605 -52237 112649 -52229
rect 112705 -52237 112749 -52229
rect 112805 -52237 112849 -52229
rect 113305 -52237 113349 -52229
rect 113405 -52237 113449 -52229
rect 113505 -52237 113549 -52229
rect 113605 -52237 113649 -52229
rect 113705 -52237 113749 -52229
rect 113805 -52237 113849 -52229
rect 113905 -52237 113949 -52229
rect 114005 -52237 114049 -52229
rect 114105 -52237 114149 -52229
rect 114205 -52237 114249 -52229
rect 114305 -52237 114349 -52229
rect 114405 -52237 114449 -52229
rect 114505 -52237 114549 -52229
rect 114605 -52237 114649 -52229
rect 114705 -52237 114749 -52229
rect 114805 -52237 114849 -52229
rect 115305 -52237 115349 -52229
rect 115405 -52237 115449 -52229
rect 115505 -52237 115549 -52229
rect 115605 -52237 115649 -52229
rect 115705 -52237 115749 -52229
rect 115805 -52237 115849 -52229
rect 115905 -52237 115949 -52229
rect 116005 -52237 116049 -52229
rect 116105 -52237 116149 -52229
rect 116205 -52237 116249 -52229
rect 116305 -52237 116349 -52229
rect 116405 -52237 116449 -52229
rect 116505 -52237 116549 -52229
rect 116605 -52237 116649 -52229
rect 116705 -52237 116749 -52229
rect 116805 -52237 116849 -52229
rect 109349 -52281 109357 -52237
rect 109449 -52281 109457 -52237
rect 109549 -52281 109557 -52237
rect 109649 -52281 109657 -52237
rect 109749 -52281 109757 -52237
rect 109849 -52281 109857 -52237
rect 109949 -52281 109957 -52237
rect 110049 -52281 110057 -52237
rect 110149 -52281 110157 -52237
rect 110249 -52281 110257 -52237
rect 110349 -52281 110357 -52237
rect 110449 -52281 110457 -52237
rect 110549 -52281 110557 -52237
rect 110649 -52281 110657 -52237
rect 110749 -52281 110757 -52237
rect 110849 -52281 110857 -52237
rect 111349 -52281 111357 -52237
rect 111449 -52281 111457 -52237
rect 111549 -52281 111557 -52237
rect 111649 -52281 111657 -52237
rect 111749 -52281 111757 -52237
rect 111849 -52281 111857 -52237
rect 111949 -52281 111957 -52237
rect 112049 -52281 112057 -52237
rect 112149 -52281 112157 -52237
rect 112249 -52281 112257 -52237
rect 112349 -52281 112357 -52237
rect 112449 -52281 112457 -52237
rect 112549 -52281 112557 -52237
rect 112649 -52281 112657 -52237
rect 112749 -52281 112757 -52237
rect 112849 -52281 112857 -52237
rect 113349 -52281 113357 -52237
rect 113449 -52281 113457 -52237
rect 113549 -52281 113557 -52237
rect 113649 -52281 113657 -52237
rect 113749 -52281 113757 -52237
rect 113849 -52281 113857 -52237
rect 113949 -52281 113957 -52237
rect 114049 -52281 114057 -52237
rect 114149 -52281 114157 -52237
rect 114249 -52281 114257 -52237
rect 114349 -52281 114357 -52237
rect 114449 -52281 114457 -52237
rect 114549 -52281 114557 -52237
rect 114649 -52281 114657 -52237
rect 114749 -52281 114757 -52237
rect 114849 -52281 114857 -52237
rect 115349 -52281 115357 -52237
rect 115449 -52281 115457 -52237
rect 115549 -52281 115557 -52237
rect 115649 -52281 115657 -52237
rect 115749 -52281 115757 -52237
rect 115849 -52281 115857 -52237
rect 115949 -52281 115957 -52237
rect 116049 -52281 116057 -52237
rect 116149 -52281 116157 -52237
rect 116249 -52281 116257 -52237
rect 116349 -52281 116357 -52237
rect 116449 -52281 116457 -52237
rect 116549 -52281 116557 -52237
rect 116649 -52281 116657 -52237
rect 116749 -52281 116757 -52237
rect 116849 -52281 116857 -52237
rect 109305 -52337 109349 -52329
rect 109405 -52337 109449 -52329
rect 109505 -52337 109549 -52329
rect 109605 -52337 109649 -52329
rect 109705 -52337 109749 -52329
rect 109805 -52337 109849 -52329
rect 109905 -52337 109949 -52329
rect 110005 -52337 110049 -52329
rect 110105 -52337 110149 -52329
rect 110205 -52337 110249 -52329
rect 110305 -52337 110349 -52329
rect 110405 -52337 110449 -52329
rect 110505 -52337 110549 -52329
rect 110605 -52337 110649 -52329
rect 110705 -52337 110749 -52329
rect 110805 -52337 110849 -52329
rect 111305 -52337 111349 -52329
rect 111405 -52337 111449 -52329
rect 111505 -52337 111549 -52329
rect 111605 -52337 111649 -52329
rect 111705 -52337 111749 -52329
rect 111805 -52337 111849 -52329
rect 111905 -52337 111949 -52329
rect 112005 -52337 112049 -52329
rect 112105 -52337 112149 -52329
rect 112205 -52337 112249 -52329
rect 112305 -52337 112349 -52329
rect 112405 -52337 112449 -52329
rect 112505 -52337 112549 -52329
rect 112605 -52337 112649 -52329
rect 112705 -52337 112749 -52329
rect 112805 -52337 112849 -52329
rect 113305 -52337 113349 -52329
rect 113405 -52337 113449 -52329
rect 113505 -52337 113549 -52329
rect 113605 -52337 113649 -52329
rect 113705 -52337 113749 -52329
rect 113805 -52337 113849 -52329
rect 113905 -52337 113949 -52329
rect 114005 -52337 114049 -52329
rect 114105 -52337 114149 -52329
rect 114205 -52337 114249 -52329
rect 114305 -52337 114349 -52329
rect 114405 -52337 114449 -52329
rect 114505 -52337 114549 -52329
rect 114605 -52337 114649 -52329
rect 114705 -52337 114749 -52329
rect 114805 -52337 114849 -52329
rect 115305 -52337 115349 -52329
rect 115405 -52337 115449 -52329
rect 115505 -52337 115549 -52329
rect 115605 -52337 115649 -52329
rect 115705 -52337 115749 -52329
rect 115805 -52337 115849 -52329
rect 115905 -52337 115949 -52329
rect 116005 -52337 116049 -52329
rect 116105 -52337 116149 -52329
rect 116205 -52337 116249 -52329
rect 116305 -52337 116349 -52329
rect 116405 -52337 116449 -52329
rect 116505 -52337 116549 -52329
rect 116605 -52337 116649 -52329
rect 116705 -52337 116749 -52329
rect 116805 -52337 116849 -52329
rect 109349 -52381 109357 -52337
rect 109449 -52381 109457 -52337
rect 109549 -52381 109557 -52337
rect 109649 -52381 109657 -52337
rect 109749 -52381 109757 -52337
rect 109849 -52381 109857 -52337
rect 109949 -52381 109957 -52337
rect 110049 -52381 110057 -52337
rect 110149 -52381 110157 -52337
rect 110249 -52381 110257 -52337
rect 110349 -52381 110357 -52337
rect 110449 -52381 110457 -52337
rect 110549 -52381 110557 -52337
rect 110649 -52381 110657 -52337
rect 110749 -52381 110757 -52337
rect 110849 -52381 110857 -52337
rect 111349 -52381 111357 -52337
rect 111449 -52381 111457 -52337
rect 111549 -52381 111557 -52337
rect 111649 -52381 111657 -52337
rect 111749 -52381 111757 -52337
rect 111849 -52381 111857 -52337
rect 111949 -52381 111957 -52337
rect 112049 -52381 112057 -52337
rect 112149 -52381 112157 -52337
rect 112249 -52381 112257 -52337
rect 112349 -52381 112357 -52337
rect 112449 -52381 112457 -52337
rect 112549 -52381 112557 -52337
rect 112649 -52381 112657 -52337
rect 112749 -52381 112757 -52337
rect 112849 -52381 112857 -52337
rect 113349 -52381 113357 -52337
rect 113449 -52381 113457 -52337
rect 113549 -52381 113557 -52337
rect 113649 -52381 113657 -52337
rect 113749 -52381 113757 -52337
rect 113849 -52381 113857 -52337
rect 113949 -52381 113957 -52337
rect 114049 -52381 114057 -52337
rect 114149 -52381 114157 -52337
rect 114249 -52381 114257 -52337
rect 114349 -52381 114357 -52337
rect 114449 -52381 114457 -52337
rect 114549 -52381 114557 -52337
rect 114649 -52381 114657 -52337
rect 114749 -52381 114757 -52337
rect 114849 -52381 114857 -52337
rect 115349 -52381 115357 -52337
rect 115449 -52381 115457 -52337
rect 115549 -52381 115557 -52337
rect 115649 -52381 115657 -52337
rect 115749 -52381 115757 -52337
rect 115849 -52381 115857 -52337
rect 115949 -52381 115957 -52337
rect 116049 -52381 116057 -52337
rect 116149 -52381 116157 -52337
rect 116249 -52381 116257 -52337
rect 116349 -52381 116357 -52337
rect 116449 -52381 116457 -52337
rect 116549 -52381 116557 -52337
rect 116649 -52381 116657 -52337
rect 116749 -52381 116757 -52337
rect 116849 -52381 116857 -52337
rect 109305 -52437 109349 -52429
rect 109405 -52437 109449 -52429
rect 109505 -52437 109549 -52429
rect 109605 -52437 109649 -52429
rect 109705 -52437 109749 -52429
rect 109805 -52437 109849 -52429
rect 109905 -52437 109949 -52429
rect 110005 -52437 110049 -52429
rect 110105 -52437 110149 -52429
rect 110205 -52437 110249 -52429
rect 110305 -52437 110349 -52429
rect 110405 -52437 110449 -52429
rect 110505 -52437 110549 -52429
rect 110605 -52437 110649 -52429
rect 110705 -52437 110749 -52429
rect 110805 -52437 110849 -52429
rect 111305 -52437 111349 -52429
rect 111405 -52437 111449 -52429
rect 111505 -52437 111549 -52429
rect 111605 -52437 111649 -52429
rect 111705 -52437 111749 -52429
rect 111805 -52437 111849 -52429
rect 111905 -52437 111949 -52429
rect 112005 -52437 112049 -52429
rect 112105 -52437 112149 -52429
rect 112205 -52437 112249 -52429
rect 112305 -52437 112349 -52429
rect 112405 -52437 112449 -52429
rect 112505 -52437 112549 -52429
rect 112605 -52437 112649 -52429
rect 112705 -52437 112749 -52429
rect 112805 -52437 112849 -52429
rect 113305 -52437 113349 -52429
rect 113405 -52437 113449 -52429
rect 113505 -52437 113549 -52429
rect 113605 -52437 113649 -52429
rect 113705 -52437 113749 -52429
rect 113805 -52437 113849 -52429
rect 113905 -52437 113949 -52429
rect 114005 -52437 114049 -52429
rect 114105 -52437 114149 -52429
rect 114205 -52437 114249 -52429
rect 114305 -52437 114349 -52429
rect 114405 -52437 114449 -52429
rect 114505 -52437 114549 -52429
rect 114605 -52437 114649 -52429
rect 114705 -52437 114749 -52429
rect 114805 -52437 114849 -52429
rect 115305 -52437 115349 -52429
rect 115405 -52437 115449 -52429
rect 115505 -52437 115549 -52429
rect 115605 -52437 115649 -52429
rect 115705 -52437 115749 -52429
rect 115805 -52437 115849 -52429
rect 115905 -52437 115949 -52429
rect 116005 -52437 116049 -52429
rect 116105 -52437 116149 -52429
rect 116205 -52437 116249 -52429
rect 116305 -52437 116349 -52429
rect 116405 -52437 116449 -52429
rect 116505 -52437 116549 -52429
rect 116605 -52437 116649 -52429
rect 116705 -52437 116749 -52429
rect 116805 -52437 116849 -52429
rect 109349 -52481 109357 -52437
rect 109449 -52481 109457 -52437
rect 109549 -52481 109557 -52437
rect 109649 -52481 109657 -52437
rect 109749 -52481 109757 -52437
rect 109849 -52481 109857 -52437
rect 109949 -52481 109957 -52437
rect 110049 -52481 110057 -52437
rect 110149 -52481 110157 -52437
rect 110249 -52481 110257 -52437
rect 110349 -52481 110357 -52437
rect 110449 -52481 110457 -52437
rect 110549 -52481 110557 -52437
rect 110649 -52481 110657 -52437
rect 110749 -52481 110757 -52437
rect 110849 -52481 110857 -52437
rect 111349 -52481 111357 -52437
rect 111449 -52481 111457 -52437
rect 111549 -52481 111557 -52437
rect 111649 -52481 111657 -52437
rect 111749 -52481 111757 -52437
rect 111849 -52481 111857 -52437
rect 111949 -52481 111957 -52437
rect 112049 -52481 112057 -52437
rect 112149 -52481 112157 -52437
rect 112249 -52481 112257 -52437
rect 112349 -52481 112357 -52437
rect 112449 -52481 112457 -52437
rect 112549 -52481 112557 -52437
rect 112649 -52481 112657 -52437
rect 112749 -52481 112757 -52437
rect 112849 -52481 112857 -52437
rect 113349 -52481 113357 -52437
rect 113449 -52481 113457 -52437
rect 113549 -52481 113557 -52437
rect 113649 -52481 113657 -52437
rect 113749 -52481 113757 -52437
rect 113849 -52481 113857 -52437
rect 113949 -52481 113957 -52437
rect 114049 -52481 114057 -52437
rect 114149 -52481 114157 -52437
rect 114249 -52481 114257 -52437
rect 114349 -52481 114357 -52437
rect 114449 -52481 114457 -52437
rect 114549 -52481 114557 -52437
rect 114649 -52481 114657 -52437
rect 114749 -52481 114757 -52437
rect 114849 -52481 114857 -52437
rect 115349 -52481 115357 -52437
rect 115449 -52481 115457 -52437
rect 115549 -52481 115557 -52437
rect 115649 -52481 115657 -52437
rect 115749 -52481 115757 -52437
rect 115849 -52481 115857 -52437
rect 115949 -52481 115957 -52437
rect 116049 -52481 116057 -52437
rect 116149 -52481 116157 -52437
rect 116249 -52481 116257 -52437
rect 116349 -52481 116357 -52437
rect 116449 -52481 116457 -52437
rect 116549 -52481 116557 -52437
rect 116649 -52481 116657 -52437
rect 116749 -52481 116757 -52437
rect 116849 -52481 116857 -52437
rect 109305 -52537 109349 -52529
rect 109405 -52537 109449 -52529
rect 109505 -52537 109549 -52529
rect 109605 -52537 109649 -52529
rect 109705 -52537 109749 -52529
rect 109805 -52537 109849 -52529
rect 109905 -52537 109949 -52529
rect 110005 -52537 110049 -52529
rect 110105 -52537 110149 -52529
rect 110205 -52537 110249 -52529
rect 110305 -52537 110349 -52529
rect 110405 -52537 110449 -52529
rect 110505 -52537 110549 -52529
rect 110605 -52537 110649 -52529
rect 110705 -52537 110749 -52529
rect 110805 -52537 110849 -52529
rect 111305 -52537 111349 -52529
rect 111405 -52537 111449 -52529
rect 111505 -52537 111549 -52529
rect 111605 -52537 111649 -52529
rect 111705 -52537 111749 -52529
rect 111805 -52537 111849 -52529
rect 111905 -52537 111949 -52529
rect 112005 -52537 112049 -52529
rect 112105 -52537 112149 -52529
rect 112205 -52537 112249 -52529
rect 112305 -52537 112349 -52529
rect 112405 -52537 112449 -52529
rect 112505 -52537 112549 -52529
rect 112605 -52537 112649 -52529
rect 112705 -52537 112749 -52529
rect 112805 -52537 112849 -52529
rect 113305 -52537 113349 -52529
rect 113405 -52537 113449 -52529
rect 113505 -52537 113549 -52529
rect 113605 -52537 113649 -52529
rect 113705 -52537 113749 -52529
rect 113805 -52537 113849 -52529
rect 113905 -52537 113949 -52529
rect 114005 -52537 114049 -52529
rect 114105 -52537 114149 -52529
rect 114205 -52537 114249 -52529
rect 114305 -52537 114349 -52529
rect 114405 -52537 114449 -52529
rect 114505 -52537 114549 -52529
rect 114605 -52537 114649 -52529
rect 114705 -52537 114749 -52529
rect 114805 -52537 114849 -52529
rect 115305 -52537 115349 -52529
rect 115405 -52537 115449 -52529
rect 115505 -52537 115549 -52529
rect 115605 -52537 115649 -52529
rect 115705 -52537 115749 -52529
rect 115805 -52537 115849 -52529
rect 115905 -52537 115949 -52529
rect 116005 -52537 116049 -52529
rect 116105 -52537 116149 -52529
rect 116205 -52537 116249 -52529
rect 116305 -52537 116349 -52529
rect 116405 -52537 116449 -52529
rect 116505 -52537 116549 -52529
rect 116605 -52537 116649 -52529
rect 116705 -52537 116749 -52529
rect 116805 -52537 116849 -52529
rect 109349 -52581 109357 -52537
rect 109449 -52581 109457 -52537
rect 109549 -52581 109557 -52537
rect 109649 -52581 109657 -52537
rect 109749 -52581 109757 -52537
rect 109849 -52581 109857 -52537
rect 109949 -52581 109957 -52537
rect 110049 -52581 110057 -52537
rect 110149 -52581 110157 -52537
rect 110249 -52581 110257 -52537
rect 110349 -52581 110357 -52537
rect 110449 -52581 110457 -52537
rect 110549 -52581 110557 -52537
rect 110649 -52581 110657 -52537
rect 110749 -52581 110757 -52537
rect 110849 -52581 110857 -52537
rect 111349 -52581 111357 -52537
rect 111449 -52581 111457 -52537
rect 111549 -52581 111557 -52537
rect 111649 -52581 111657 -52537
rect 111749 -52581 111757 -52537
rect 111849 -52581 111857 -52537
rect 111949 -52581 111957 -52537
rect 112049 -52581 112057 -52537
rect 112149 -52581 112157 -52537
rect 112249 -52581 112257 -52537
rect 112349 -52581 112357 -52537
rect 112449 -52581 112457 -52537
rect 112549 -52581 112557 -52537
rect 112649 -52581 112657 -52537
rect 112749 -52581 112757 -52537
rect 112849 -52581 112857 -52537
rect 113349 -52581 113357 -52537
rect 113449 -52581 113457 -52537
rect 113549 -52581 113557 -52537
rect 113649 -52581 113657 -52537
rect 113749 -52581 113757 -52537
rect 113849 -52581 113857 -52537
rect 113949 -52581 113957 -52537
rect 114049 -52581 114057 -52537
rect 114149 -52581 114157 -52537
rect 114249 -52581 114257 -52537
rect 114349 -52581 114357 -52537
rect 114449 -52581 114457 -52537
rect 114549 -52581 114557 -52537
rect 114649 -52581 114657 -52537
rect 114749 -52581 114757 -52537
rect 114849 -52581 114857 -52537
rect 115349 -52581 115357 -52537
rect 115449 -52581 115457 -52537
rect 115549 -52581 115557 -52537
rect 115649 -52581 115657 -52537
rect 115749 -52581 115757 -52537
rect 115849 -52581 115857 -52537
rect 115949 -52581 115957 -52537
rect 116049 -52581 116057 -52537
rect 116149 -52581 116157 -52537
rect 116249 -52581 116257 -52537
rect 116349 -52581 116357 -52537
rect 116449 -52581 116457 -52537
rect 116549 -52581 116557 -52537
rect 116649 -52581 116657 -52537
rect 116749 -52581 116757 -52537
rect 116849 -52581 116857 -52537
rect 109305 -52637 109349 -52629
rect 109405 -52637 109449 -52629
rect 109505 -52637 109549 -52629
rect 109605 -52637 109649 -52629
rect 109705 -52637 109749 -52629
rect 109805 -52637 109849 -52629
rect 109905 -52637 109949 -52629
rect 110005 -52637 110049 -52629
rect 110105 -52637 110149 -52629
rect 110205 -52637 110249 -52629
rect 110305 -52637 110349 -52629
rect 110405 -52637 110449 -52629
rect 110505 -52637 110549 -52629
rect 110605 -52637 110649 -52629
rect 110705 -52637 110749 -52629
rect 110805 -52637 110849 -52629
rect 111305 -52637 111349 -52629
rect 111405 -52637 111449 -52629
rect 111505 -52637 111549 -52629
rect 111605 -52637 111649 -52629
rect 111705 -52637 111749 -52629
rect 111805 -52637 111849 -52629
rect 111905 -52637 111949 -52629
rect 112005 -52637 112049 -52629
rect 112105 -52637 112149 -52629
rect 112205 -52637 112249 -52629
rect 112305 -52637 112349 -52629
rect 112405 -52637 112449 -52629
rect 112505 -52637 112549 -52629
rect 112605 -52637 112649 -52629
rect 112705 -52637 112749 -52629
rect 112805 -52637 112849 -52629
rect 113305 -52637 113349 -52629
rect 113405 -52637 113449 -52629
rect 113505 -52637 113549 -52629
rect 113605 -52637 113649 -52629
rect 113705 -52637 113749 -52629
rect 113805 -52637 113849 -52629
rect 113905 -52637 113949 -52629
rect 114005 -52637 114049 -52629
rect 114105 -52637 114149 -52629
rect 114205 -52637 114249 -52629
rect 114305 -52637 114349 -52629
rect 114405 -52637 114449 -52629
rect 114505 -52637 114549 -52629
rect 114605 -52637 114649 -52629
rect 114705 -52637 114749 -52629
rect 114805 -52637 114849 -52629
rect 115305 -52637 115349 -52629
rect 115405 -52637 115449 -52629
rect 115505 -52637 115549 -52629
rect 115605 -52637 115649 -52629
rect 115705 -52637 115749 -52629
rect 115805 -52637 115849 -52629
rect 115905 -52637 115949 -52629
rect 116005 -52637 116049 -52629
rect 116105 -52637 116149 -52629
rect 116205 -52637 116249 -52629
rect 116305 -52637 116349 -52629
rect 116405 -52637 116449 -52629
rect 116505 -52637 116549 -52629
rect 116605 -52637 116649 -52629
rect 116705 -52637 116749 -52629
rect 116805 -52637 116849 -52629
rect 109349 -52681 109357 -52637
rect 109449 -52681 109457 -52637
rect 109549 -52681 109557 -52637
rect 109649 -52681 109657 -52637
rect 109749 -52681 109757 -52637
rect 109849 -52681 109857 -52637
rect 109949 -52681 109957 -52637
rect 110049 -52681 110057 -52637
rect 110149 -52681 110157 -52637
rect 110249 -52681 110257 -52637
rect 110349 -52681 110357 -52637
rect 110449 -52681 110457 -52637
rect 110549 -52681 110557 -52637
rect 110649 -52681 110657 -52637
rect 110749 -52681 110757 -52637
rect 110849 -52681 110857 -52637
rect 111349 -52681 111357 -52637
rect 111449 -52681 111457 -52637
rect 111549 -52681 111557 -52637
rect 111649 -52681 111657 -52637
rect 111749 -52681 111757 -52637
rect 111849 -52681 111857 -52637
rect 111949 -52681 111957 -52637
rect 112049 -52681 112057 -52637
rect 112149 -52681 112157 -52637
rect 112249 -52681 112257 -52637
rect 112349 -52681 112357 -52637
rect 112449 -52681 112457 -52637
rect 112549 -52681 112557 -52637
rect 112649 -52681 112657 -52637
rect 112749 -52681 112757 -52637
rect 112849 -52681 112857 -52637
rect 113349 -52681 113357 -52637
rect 113449 -52681 113457 -52637
rect 113549 -52681 113557 -52637
rect 113649 -52681 113657 -52637
rect 113749 -52681 113757 -52637
rect 113849 -52681 113857 -52637
rect 113949 -52681 113957 -52637
rect 114049 -52681 114057 -52637
rect 114149 -52681 114157 -52637
rect 114249 -52681 114257 -52637
rect 114349 -52681 114357 -52637
rect 114449 -52681 114457 -52637
rect 114549 -52681 114557 -52637
rect 114649 -52681 114657 -52637
rect 114749 -52681 114757 -52637
rect 114849 -52681 114857 -52637
rect 115349 -52681 115357 -52637
rect 115449 -52681 115457 -52637
rect 115549 -52681 115557 -52637
rect 115649 -52681 115657 -52637
rect 115749 -52681 115757 -52637
rect 115849 -52681 115857 -52637
rect 115949 -52681 115957 -52637
rect 116049 -52681 116057 -52637
rect 116149 -52681 116157 -52637
rect 116249 -52681 116257 -52637
rect 116349 -52681 116357 -52637
rect 116449 -52681 116457 -52637
rect 116549 -52681 116557 -52637
rect 116649 -52681 116657 -52637
rect 116749 -52681 116757 -52637
rect 116849 -52681 116857 -52637
rect -109180 -74119 -109178 -54119
rect -109114 -74119 -109112 -54119
rect -77180 -74119 -77178 -54119
rect -77114 -74119 -77112 -54119
rect -45180 -74119 -45178 -54119
rect -45114 -74119 -45112 -54119
rect -13180 -74119 -13178 -54119
rect -13114 -74119 -13112 -54119
rect 18820 -74119 18822 -54119
rect 18886 -74119 18888 -54119
rect 50820 -74119 50822 -54119
rect 50886 -74119 50888 -54119
rect 82820 -74119 82822 -54119
rect 82886 -74119 82888 -54119
rect 114820 -74119 114822 -54119
rect 114886 -74119 114888 -54119
rect 146820 -74119 146822 -54119
rect 146886 -74119 146888 -54119
rect 9236 -75188 9280 -75180
rect 9336 -75188 9380 -75180
rect 9436 -75188 9480 -75180
rect 9536 -75188 9580 -75180
rect 9636 -75188 9680 -75180
rect 9736 -75188 9780 -75180
rect 9836 -75188 9880 -75180
rect 9936 -75188 9980 -75180
rect 10036 -75188 10080 -75180
rect 10136 -75188 10180 -75180
rect 10236 -75188 10280 -75180
rect 10336 -75188 10380 -75180
rect 10436 -75188 10480 -75180
rect 10536 -75188 10580 -75180
rect 10636 -75188 10680 -75180
rect 10736 -75188 10780 -75180
rect 11236 -75188 11280 -75180
rect 11336 -75188 11380 -75180
rect 11436 -75188 11480 -75180
rect 11536 -75188 11580 -75180
rect 11636 -75188 11680 -75180
rect 11736 -75188 11780 -75180
rect 11836 -75188 11880 -75180
rect 11936 -75188 11980 -75180
rect 12036 -75188 12080 -75180
rect 12136 -75188 12180 -75180
rect 12236 -75188 12280 -75180
rect 12336 -75188 12380 -75180
rect 12436 -75188 12480 -75180
rect 12536 -75188 12580 -75180
rect 12636 -75188 12680 -75180
rect 12736 -75188 12780 -75180
rect 13236 -75188 13280 -75180
rect 13336 -75188 13380 -75180
rect 13436 -75188 13480 -75180
rect 13536 -75188 13580 -75180
rect 13636 -75188 13680 -75180
rect 13736 -75188 13780 -75180
rect 13836 -75188 13880 -75180
rect 13936 -75188 13980 -75180
rect 14036 -75188 14080 -75180
rect 14136 -75188 14180 -75180
rect 14236 -75188 14280 -75180
rect 14336 -75188 14380 -75180
rect 14436 -75188 14480 -75180
rect 14536 -75188 14580 -75180
rect 14636 -75188 14680 -75180
rect 14736 -75188 14780 -75180
rect 15236 -75188 15280 -75180
rect 15336 -75188 15380 -75180
rect 15436 -75188 15480 -75180
rect 15536 -75188 15580 -75180
rect 15636 -75188 15680 -75180
rect 15736 -75188 15780 -75180
rect 15836 -75188 15880 -75180
rect 15936 -75188 15980 -75180
rect 16036 -75188 16080 -75180
rect 16136 -75188 16180 -75180
rect 16236 -75188 16280 -75180
rect 16336 -75188 16380 -75180
rect 16436 -75188 16480 -75180
rect 16536 -75188 16580 -75180
rect 16636 -75188 16680 -75180
rect 16736 -75188 16780 -75180
rect 9280 -75232 9288 -75188
rect 9380 -75232 9388 -75188
rect 9480 -75232 9488 -75188
rect 9580 -75232 9588 -75188
rect 9680 -75232 9688 -75188
rect 9780 -75232 9788 -75188
rect 9880 -75232 9888 -75188
rect 9980 -75232 9988 -75188
rect 10080 -75232 10088 -75188
rect 10180 -75232 10188 -75188
rect 10280 -75232 10288 -75188
rect 10380 -75232 10388 -75188
rect 10480 -75232 10488 -75188
rect 10580 -75232 10588 -75188
rect 10680 -75232 10688 -75188
rect 10780 -75232 10788 -75188
rect 11280 -75232 11288 -75188
rect 11380 -75232 11388 -75188
rect 11480 -75232 11488 -75188
rect 11580 -75232 11588 -75188
rect 11680 -75232 11688 -75188
rect 11780 -75232 11788 -75188
rect 11880 -75232 11888 -75188
rect 11980 -75232 11988 -75188
rect 12080 -75232 12088 -75188
rect 12180 -75232 12188 -75188
rect 12280 -75232 12288 -75188
rect 12380 -75232 12388 -75188
rect 12480 -75232 12488 -75188
rect 12580 -75232 12588 -75188
rect 12680 -75232 12688 -75188
rect 12780 -75232 12788 -75188
rect 13280 -75232 13288 -75188
rect 13380 -75232 13388 -75188
rect 13480 -75232 13488 -75188
rect 13580 -75232 13588 -75188
rect 13680 -75232 13688 -75188
rect 13780 -75232 13788 -75188
rect 13880 -75232 13888 -75188
rect 13980 -75232 13988 -75188
rect 14080 -75232 14088 -75188
rect 14180 -75232 14188 -75188
rect 14280 -75232 14288 -75188
rect 14380 -75232 14388 -75188
rect 14480 -75232 14488 -75188
rect 14580 -75232 14588 -75188
rect 14680 -75232 14688 -75188
rect 14780 -75232 14788 -75188
rect 15280 -75232 15288 -75188
rect 15380 -75232 15388 -75188
rect 15480 -75232 15488 -75188
rect 15580 -75232 15588 -75188
rect 15680 -75232 15688 -75188
rect 15780 -75232 15788 -75188
rect 15880 -75232 15888 -75188
rect 15980 -75232 15988 -75188
rect 16080 -75232 16088 -75188
rect 16180 -75232 16188 -75188
rect 16280 -75232 16288 -75188
rect 16380 -75232 16388 -75188
rect 16480 -75232 16488 -75188
rect 16580 -75232 16588 -75188
rect 16680 -75232 16688 -75188
rect 16780 -75232 16788 -75188
rect 9236 -75288 9280 -75280
rect 9336 -75288 9380 -75280
rect 9436 -75288 9480 -75280
rect 9536 -75288 9580 -75280
rect 9636 -75288 9680 -75280
rect 9736 -75288 9780 -75280
rect 9836 -75288 9880 -75280
rect 9936 -75288 9980 -75280
rect 10036 -75288 10080 -75280
rect 10136 -75288 10180 -75280
rect 10236 -75288 10280 -75280
rect 10336 -75288 10380 -75280
rect 10436 -75288 10480 -75280
rect 10536 -75288 10580 -75280
rect 10636 -75288 10680 -75280
rect 10736 -75288 10780 -75280
rect 11236 -75288 11280 -75280
rect 11336 -75288 11380 -75280
rect 11436 -75288 11480 -75280
rect 11536 -75288 11580 -75280
rect 11636 -75288 11680 -75280
rect 11736 -75288 11780 -75280
rect 11836 -75288 11880 -75280
rect 11936 -75288 11980 -75280
rect 12036 -75288 12080 -75280
rect 12136 -75288 12180 -75280
rect 12236 -75288 12280 -75280
rect 12336 -75288 12380 -75280
rect 12436 -75288 12480 -75280
rect 12536 -75288 12580 -75280
rect 12636 -75288 12680 -75280
rect 12736 -75288 12780 -75280
rect 13236 -75288 13280 -75280
rect 13336 -75288 13380 -75280
rect 13436 -75288 13480 -75280
rect 13536 -75288 13580 -75280
rect 13636 -75288 13680 -75280
rect 13736 -75288 13780 -75280
rect 13836 -75288 13880 -75280
rect 13936 -75288 13980 -75280
rect 14036 -75288 14080 -75280
rect 14136 -75288 14180 -75280
rect 14236 -75288 14280 -75280
rect 14336 -75288 14380 -75280
rect 14436 -75288 14480 -75280
rect 14536 -75288 14580 -75280
rect 14636 -75288 14680 -75280
rect 14736 -75288 14780 -75280
rect 15236 -75288 15280 -75280
rect 15336 -75288 15380 -75280
rect 15436 -75288 15480 -75280
rect 15536 -75288 15580 -75280
rect 15636 -75288 15680 -75280
rect 15736 -75288 15780 -75280
rect 15836 -75288 15880 -75280
rect 15936 -75288 15980 -75280
rect 16036 -75288 16080 -75280
rect 16136 -75288 16180 -75280
rect 16236 -75288 16280 -75280
rect 16336 -75288 16380 -75280
rect 16436 -75288 16480 -75280
rect 16536 -75288 16580 -75280
rect 16636 -75288 16680 -75280
rect 16736 -75288 16780 -75280
rect 9280 -75332 9288 -75288
rect 9380 -75332 9388 -75288
rect 9480 -75332 9488 -75288
rect 9580 -75332 9588 -75288
rect 9680 -75332 9688 -75288
rect 9780 -75332 9788 -75288
rect 9880 -75332 9888 -75288
rect 9980 -75332 9988 -75288
rect 10080 -75332 10088 -75288
rect 10180 -75332 10188 -75288
rect 10280 -75332 10288 -75288
rect 10380 -75332 10388 -75288
rect 10480 -75332 10488 -75288
rect 10580 -75332 10588 -75288
rect 10680 -75332 10688 -75288
rect 10780 -75332 10788 -75288
rect 11280 -75332 11288 -75288
rect 11380 -75332 11388 -75288
rect 11480 -75332 11488 -75288
rect 11580 -75332 11588 -75288
rect 11680 -75332 11688 -75288
rect 11780 -75332 11788 -75288
rect 11880 -75332 11888 -75288
rect 11980 -75332 11988 -75288
rect 12080 -75332 12088 -75288
rect 12180 -75332 12188 -75288
rect 12280 -75332 12288 -75288
rect 12380 -75332 12388 -75288
rect 12480 -75332 12488 -75288
rect 12580 -75332 12588 -75288
rect 12680 -75332 12688 -75288
rect 12780 -75332 12788 -75288
rect 13280 -75332 13288 -75288
rect 13380 -75332 13388 -75288
rect 13480 -75332 13488 -75288
rect 13580 -75332 13588 -75288
rect 13680 -75332 13688 -75288
rect 13780 -75332 13788 -75288
rect 13880 -75332 13888 -75288
rect 13980 -75332 13988 -75288
rect 14080 -75332 14088 -75288
rect 14180 -75332 14188 -75288
rect 14280 -75332 14288 -75288
rect 14380 -75332 14388 -75288
rect 14480 -75332 14488 -75288
rect 14580 -75332 14588 -75288
rect 14680 -75332 14688 -75288
rect 14780 -75332 14788 -75288
rect 15280 -75332 15288 -75288
rect 15380 -75332 15388 -75288
rect 15480 -75332 15488 -75288
rect 15580 -75332 15588 -75288
rect 15680 -75332 15688 -75288
rect 15780 -75332 15788 -75288
rect 15880 -75332 15888 -75288
rect 15980 -75332 15988 -75288
rect 16080 -75332 16088 -75288
rect 16180 -75332 16188 -75288
rect 16280 -75332 16288 -75288
rect 16380 -75332 16388 -75288
rect 16480 -75332 16488 -75288
rect 16580 -75332 16588 -75288
rect 16680 -75332 16688 -75288
rect 16780 -75332 16788 -75288
rect 9236 -75388 9280 -75380
rect 9336 -75388 9380 -75380
rect 9436 -75388 9480 -75380
rect 9536 -75388 9580 -75380
rect 9636 -75388 9680 -75380
rect 9736 -75388 9780 -75380
rect 9836 -75388 9880 -75380
rect 9936 -75388 9980 -75380
rect 10036 -75388 10080 -75380
rect 10136 -75388 10180 -75380
rect 10236 -75388 10280 -75380
rect 10336 -75388 10380 -75380
rect 10436 -75388 10480 -75380
rect 10536 -75388 10580 -75380
rect 10636 -75388 10680 -75380
rect 10736 -75388 10780 -75380
rect 11236 -75388 11280 -75380
rect 11336 -75388 11380 -75380
rect 11436 -75388 11480 -75380
rect 11536 -75388 11580 -75380
rect 11636 -75388 11680 -75380
rect 11736 -75388 11780 -75380
rect 11836 -75388 11880 -75380
rect 11936 -75388 11980 -75380
rect 12036 -75388 12080 -75380
rect 12136 -75388 12180 -75380
rect 12236 -75388 12280 -75380
rect 12336 -75388 12380 -75380
rect 12436 -75388 12480 -75380
rect 12536 -75388 12580 -75380
rect 12636 -75388 12680 -75380
rect 12736 -75388 12780 -75380
rect 13236 -75388 13280 -75380
rect 13336 -75388 13380 -75380
rect 13436 -75388 13480 -75380
rect 13536 -75388 13580 -75380
rect 13636 -75388 13680 -75380
rect 13736 -75388 13780 -75380
rect 13836 -75388 13880 -75380
rect 13936 -75388 13980 -75380
rect 14036 -75388 14080 -75380
rect 14136 -75388 14180 -75380
rect 14236 -75388 14280 -75380
rect 14336 -75388 14380 -75380
rect 14436 -75388 14480 -75380
rect 14536 -75388 14580 -75380
rect 14636 -75388 14680 -75380
rect 14736 -75388 14780 -75380
rect 15236 -75388 15280 -75380
rect 15336 -75388 15380 -75380
rect 15436 -75388 15480 -75380
rect 15536 -75388 15580 -75380
rect 15636 -75388 15680 -75380
rect 15736 -75388 15780 -75380
rect 15836 -75388 15880 -75380
rect 15936 -75388 15980 -75380
rect 16036 -75388 16080 -75380
rect 16136 -75388 16180 -75380
rect 16236 -75388 16280 -75380
rect 16336 -75388 16380 -75380
rect 16436 -75388 16480 -75380
rect 16536 -75388 16580 -75380
rect 16636 -75388 16680 -75380
rect 16736 -75388 16780 -75380
rect 9280 -75432 9288 -75388
rect 9380 -75432 9388 -75388
rect 9480 -75432 9488 -75388
rect 9580 -75432 9588 -75388
rect 9680 -75432 9688 -75388
rect 9780 -75432 9788 -75388
rect 9880 -75432 9888 -75388
rect 9980 -75432 9988 -75388
rect 10080 -75432 10088 -75388
rect 10180 -75432 10188 -75388
rect 10280 -75432 10288 -75388
rect 10380 -75432 10388 -75388
rect 10480 -75432 10488 -75388
rect 10580 -75432 10588 -75388
rect 10680 -75432 10688 -75388
rect 10780 -75432 10788 -75388
rect 11280 -75432 11288 -75388
rect 11380 -75432 11388 -75388
rect 11480 -75432 11488 -75388
rect 11580 -75432 11588 -75388
rect 11680 -75432 11688 -75388
rect 11780 -75432 11788 -75388
rect 11880 -75432 11888 -75388
rect 11980 -75432 11988 -75388
rect 12080 -75432 12088 -75388
rect 12180 -75432 12188 -75388
rect 12280 -75432 12288 -75388
rect 12380 -75432 12388 -75388
rect 12480 -75432 12488 -75388
rect 12580 -75432 12588 -75388
rect 12680 -75432 12688 -75388
rect 12780 -75432 12788 -75388
rect 13280 -75432 13288 -75388
rect 13380 -75432 13388 -75388
rect 13480 -75432 13488 -75388
rect 13580 -75432 13588 -75388
rect 13680 -75432 13688 -75388
rect 13780 -75432 13788 -75388
rect 13880 -75432 13888 -75388
rect 13980 -75432 13988 -75388
rect 14080 -75432 14088 -75388
rect 14180 -75432 14188 -75388
rect 14280 -75432 14288 -75388
rect 14380 -75432 14388 -75388
rect 14480 -75432 14488 -75388
rect 14580 -75432 14588 -75388
rect 14680 -75432 14688 -75388
rect 14780 -75432 14788 -75388
rect 15280 -75432 15288 -75388
rect 15380 -75432 15388 -75388
rect 15480 -75432 15488 -75388
rect 15580 -75432 15588 -75388
rect 15680 -75432 15688 -75388
rect 15780 -75432 15788 -75388
rect 15880 -75432 15888 -75388
rect 15980 -75432 15988 -75388
rect 16080 -75432 16088 -75388
rect 16180 -75432 16188 -75388
rect 16280 -75432 16288 -75388
rect 16380 -75432 16388 -75388
rect 16480 -75432 16488 -75388
rect 16580 -75432 16588 -75388
rect 16680 -75432 16688 -75388
rect 16780 -75432 16788 -75388
rect 9236 -75488 9280 -75480
rect 9336 -75488 9380 -75480
rect 9436 -75488 9480 -75480
rect 9536 -75488 9580 -75480
rect 9636 -75488 9680 -75480
rect 9736 -75488 9780 -75480
rect 9836 -75488 9880 -75480
rect 9936 -75488 9980 -75480
rect 10036 -75488 10080 -75480
rect 10136 -75488 10180 -75480
rect 10236 -75488 10280 -75480
rect 10336 -75488 10380 -75480
rect 10436 -75488 10480 -75480
rect 10536 -75488 10580 -75480
rect 10636 -75488 10680 -75480
rect 10736 -75488 10780 -75480
rect 11236 -75488 11280 -75480
rect 11336 -75488 11380 -75480
rect 11436 -75488 11480 -75480
rect 11536 -75488 11580 -75480
rect 11636 -75488 11680 -75480
rect 11736 -75488 11780 -75480
rect 11836 -75488 11880 -75480
rect 11936 -75488 11980 -75480
rect 12036 -75488 12080 -75480
rect 12136 -75488 12180 -75480
rect 12236 -75488 12280 -75480
rect 12336 -75488 12380 -75480
rect 12436 -75488 12480 -75480
rect 12536 -75488 12580 -75480
rect 12636 -75488 12680 -75480
rect 12736 -75488 12780 -75480
rect 13236 -75488 13280 -75480
rect 13336 -75488 13380 -75480
rect 13436 -75488 13480 -75480
rect 13536 -75488 13580 -75480
rect 13636 -75488 13680 -75480
rect 13736 -75488 13780 -75480
rect 13836 -75488 13880 -75480
rect 13936 -75488 13980 -75480
rect 14036 -75488 14080 -75480
rect 14136 -75488 14180 -75480
rect 14236 -75488 14280 -75480
rect 14336 -75488 14380 -75480
rect 14436 -75488 14480 -75480
rect 14536 -75488 14580 -75480
rect 14636 -75488 14680 -75480
rect 14736 -75488 14780 -75480
rect 15236 -75488 15280 -75480
rect 15336 -75488 15380 -75480
rect 15436 -75488 15480 -75480
rect 15536 -75488 15580 -75480
rect 15636 -75488 15680 -75480
rect 15736 -75488 15780 -75480
rect 15836 -75488 15880 -75480
rect 15936 -75488 15980 -75480
rect 16036 -75488 16080 -75480
rect 16136 -75488 16180 -75480
rect 16236 -75488 16280 -75480
rect 16336 -75488 16380 -75480
rect 16436 -75488 16480 -75480
rect 16536 -75488 16580 -75480
rect 16636 -75488 16680 -75480
rect 16736 -75488 16780 -75480
rect 9280 -75532 9288 -75488
rect 9380 -75532 9388 -75488
rect 9480 -75532 9488 -75488
rect 9580 -75532 9588 -75488
rect 9680 -75532 9688 -75488
rect 9780 -75532 9788 -75488
rect 9880 -75532 9888 -75488
rect 9980 -75532 9988 -75488
rect 10080 -75532 10088 -75488
rect 10180 -75532 10188 -75488
rect 10280 -75532 10288 -75488
rect 10380 -75532 10388 -75488
rect 10480 -75532 10488 -75488
rect 10580 -75532 10588 -75488
rect 10680 -75532 10688 -75488
rect 10780 -75532 10788 -75488
rect 11280 -75532 11288 -75488
rect 11380 -75532 11388 -75488
rect 11480 -75532 11488 -75488
rect 11580 -75532 11588 -75488
rect 11680 -75532 11688 -75488
rect 11780 -75532 11788 -75488
rect 11880 -75532 11888 -75488
rect 11980 -75532 11988 -75488
rect 12080 -75532 12088 -75488
rect 12180 -75532 12188 -75488
rect 12280 -75532 12288 -75488
rect 12380 -75532 12388 -75488
rect 12480 -75532 12488 -75488
rect 12580 -75532 12588 -75488
rect 12680 -75532 12688 -75488
rect 12780 -75532 12788 -75488
rect 13280 -75532 13288 -75488
rect 13380 -75532 13388 -75488
rect 13480 -75532 13488 -75488
rect 13580 -75532 13588 -75488
rect 13680 -75532 13688 -75488
rect 13780 -75532 13788 -75488
rect 13880 -75532 13888 -75488
rect 13980 -75532 13988 -75488
rect 14080 -75532 14088 -75488
rect 14180 -75532 14188 -75488
rect 14280 -75532 14288 -75488
rect 14380 -75532 14388 -75488
rect 14480 -75532 14488 -75488
rect 14580 -75532 14588 -75488
rect 14680 -75532 14688 -75488
rect 14780 -75532 14788 -75488
rect 15280 -75532 15288 -75488
rect 15380 -75532 15388 -75488
rect 15480 -75532 15488 -75488
rect 15580 -75532 15588 -75488
rect 15680 -75532 15688 -75488
rect 15780 -75532 15788 -75488
rect 15880 -75532 15888 -75488
rect 15980 -75532 15988 -75488
rect 16080 -75532 16088 -75488
rect 16180 -75532 16188 -75488
rect 16280 -75532 16288 -75488
rect 16380 -75532 16388 -75488
rect 16480 -75532 16488 -75488
rect 16580 -75532 16588 -75488
rect 16680 -75532 16688 -75488
rect 16780 -75532 16788 -75488
rect 9236 -75588 9280 -75580
rect 9336 -75588 9380 -75580
rect 9436 -75588 9480 -75580
rect 9536 -75588 9580 -75580
rect 9636 -75588 9680 -75580
rect 9736 -75588 9780 -75580
rect 9836 -75588 9880 -75580
rect 9936 -75588 9980 -75580
rect 10036 -75588 10080 -75580
rect 10136 -75588 10180 -75580
rect 10236 -75588 10280 -75580
rect 10336 -75588 10380 -75580
rect 10436 -75588 10480 -75580
rect 10536 -75588 10580 -75580
rect 10636 -75588 10680 -75580
rect 10736 -75588 10780 -75580
rect 11236 -75588 11280 -75580
rect 11336 -75588 11380 -75580
rect 11436 -75588 11480 -75580
rect 11536 -75588 11580 -75580
rect 11636 -75588 11680 -75580
rect 11736 -75588 11780 -75580
rect 11836 -75588 11880 -75580
rect 11936 -75588 11980 -75580
rect 12036 -75588 12080 -75580
rect 12136 -75588 12180 -75580
rect 12236 -75588 12280 -75580
rect 12336 -75588 12380 -75580
rect 12436 -75588 12480 -75580
rect 12536 -75588 12580 -75580
rect 12636 -75588 12680 -75580
rect 12736 -75588 12780 -75580
rect 13236 -75588 13280 -75580
rect 13336 -75588 13380 -75580
rect 13436 -75588 13480 -75580
rect 13536 -75588 13580 -75580
rect 13636 -75588 13680 -75580
rect 13736 -75588 13780 -75580
rect 13836 -75588 13880 -75580
rect 13936 -75588 13980 -75580
rect 14036 -75588 14080 -75580
rect 14136 -75588 14180 -75580
rect 14236 -75588 14280 -75580
rect 14336 -75588 14380 -75580
rect 14436 -75588 14480 -75580
rect 14536 -75588 14580 -75580
rect 14636 -75588 14680 -75580
rect 14736 -75588 14780 -75580
rect 15236 -75588 15280 -75580
rect 15336 -75588 15380 -75580
rect 15436 -75588 15480 -75580
rect 15536 -75588 15580 -75580
rect 15636 -75588 15680 -75580
rect 15736 -75588 15780 -75580
rect 15836 -75588 15880 -75580
rect 15936 -75588 15980 -75580
rect 16036 -75588 16080 -75580
rect 16136 -75588 16180 -75580
rect 16236 -75588 16280 -75580
rect 16336 -75588 16380 -75580
rect 16436 -75588 16480 -75580
rect 16536 -75588 16580 -75580
rect 16636 -75588 16680 -75580
rect 16736 -75588 16780 -75580
rect 9280 -75632 9288 -75588
rect 9380 -75632 9388 -75588
rect 9480 -75632 9488 -75588
rect 9580 -75632 9588 -75588
rect 9680 -75632 9688 -75588
rect 9780 -75632 9788 -75588
rect 9880 -75632 9888 -75588
rect 9980 -75632 9988 -75588
rect 10080 -75632 10088 -75588
rect 10180 -75632 10188 -75588
rect 10280 -75632 10288 -75588
rect 10380 -75632 10388 -75588
rect 10480 -75632 10488 -75588
rect 10580 -75632 10588 -75588
rect 10680 -75632 10688 -75588
rect 10780 -75632 10788 -75588
rect 11280 -75632 11288 -75588
rect 11380 -75632 11388 -75588
rect 11480 -75632 11488 -75588
rect 11580 -75632 11588 -75588
rect 11680 -75632 11688 -75588
rect 11780 -75632 11788 -75588
rect 11880 -75632 11888 -75588
rect 11980 -75632 11988 -75588
rect 12080 -75632 12088 -75588
rect 12180 -75632 12188 -75588
rect 12280 -75632 12288 -75588
rect 12380 -75632 12388 -75588
rect 12480 -75632 12488 -75588
rect 12580 -75632 12588 -75588
rect 12680 -75632 12688 -75588
rect 12780 -75632 12788 -75588
rect 13280 -75632 13288 -75588
rect 13380 -75632 13388 -75588
rect 13480 -75632 13488 -75588
rect 13580 -75632 13588 -75588
rect 13680 -75632 13688 -75588
rect 13780 -75632 13788 -75588
rect 13880 -75632 13888 -75588
rect 13980 -75632 13988 -75588
rect 14080 -75632 14088 -75588
rect 14180 -75632 14188 -75588
rect 14280 -75632 14288 -75588
rect 14380 -75632 14388 -75588
rect 14480 -75632 14488 -75588
rect 14580 -75632 14588 -75588
rect 14680 -75632 14688 -75588
rect 14780 -75632 14788 -75588
rect 15280 -75632 15288 -75588
rect 15380 -75632 15388 -75588
rect 15480 -75632 15488 -75588
rect 15580 -75632 15588 -75588
rect 15680 -75632 15688 -75588
rect 15780 -75632 15788 -75588
rect 15880 -75632 15888 -75588
rect 15980 -75632 15988 -75588
rect 16080 -75632 16088 -75588
rect 16180 -75632 16188 -75588
rect 16280 -75632 16288 -75588
rect 16380 -75632 16388 -75588
rect 16480 -75632 16488 -75588
rect 16580 -75632 16588 -75588
rect 16680 -75632 16688 -75588
rect 16780 -75632 16788 -75588
rect 9236 -75688 9280 -75680
rect 9336 -75688 9380 -75680
rect 9436 -75688 9480 -75680
rect 9536 -75688 9580 -75680
rect 9636 -75688 9680 -75680
rect 9736 -75688 9780 -75680
rect 9836 -75688 9880 -75680
rect 9936 -75688 9980 -75680
rect 10036 -75688 10080 -75680
rect 10136 -75688 10180 -75680
rect 10236 -75688 10280 -75680
rect 10336 -75688 10380 -75680
rect 10436 -75688 10480 -75680
rect 10536 -75688 10580 -75680
rect 10636 -75688 10680 -75680
rect 10736 -75688 10780 -75680
rect 11236 -75688 11280 -75680
rect 11336 -75688 11380 -75680
rect 11436 -75688 11480 -75680
rect 11536 -75688 11580 -75680
rect 11636 -75688 11680 -75680
rect 11736 -75688 11780 -75680
rect 11836 -75688 11880 -75680
rect 11936 -75688 11980 -75680
rect 12036 -75688 12080 -75680
rect 12136 -75688 12180 -75680
rect 12236 -75688 12280 -75680
rect 12336 -75688 12380 -75680
rect 12436 -75688 12480 -75680
rect 12536 -75688 12580 -75680
rect 12636 -75688 12680 -75680
rect 12736 -75688 12780 -75680
rect 13236 -75688 13280 -75680
rect 13336 -75688 13380 -75680
rect 13436 -75688 13480 -75680
rect 13536 -75688 13580 -75680
rect 13636 -75688 13680 -75680
rect 13736 -75688 13780 -75680
rect 13836 -75688 13880 -75680
rect 13936 -75688 13980 -75680
rect 14036 -75688 14080 -75680
rect 14136 -75688 14180 -75680
rect 14236 -75688 14280 -75680
rect 14336 -75688 14380 -75680
rect 14436 -75688 14480 -75680
rect 14536 -75688 14580 -75680
rect 14636 -75688 14680 -75680
rect 14736 -75688 14780 -75680
rect 15236 -75688 15280 -75680
rect 15336 -75688 15380 -75680
rect 15436 -75688 15480 -75680
rect 15536 -75688 15580 -75680
rect 15636 -75688 15680 -75680
rect 15736 -75688 15780 -75680
rect 15836 -75688 15880 -75680
rect 15936 -75688 15980 -75680
rect 16036 -75688 16080 -75680
rect 16136 -75688 16180 -75680
rect 16236 -75688 16280 -75680
rect 16336 -75688 16380 -75680
rect 16436 -75688 16480 -75680
rect 16536 -75688 16580 -75680
rect 16636 -75688 16680 -75680
rect 16736 -75688 16780 -75680
rect 9280 -75732 9288 -75688
rect 9380 -75732 9388 -75688
rect 9480 -75732 9488 -75688
rect 9580 -75732 9588 -75688
rect 9680 -75732 9688 -75688
rect 9780 -75732 9788 -75688
rect 9880 -75732 9888 -75688
rect 9980 -75732 9988 -75688
rect 10080 -75732 10088 -75688
rect 10180 -75732 10188 -75688
rect 10280 -75732 10288 -75688
rect 10380 -75732 10388 -75688
rect 10480 -75732 10488 -75688
rect 10580 -75732 10588 -75688
rect 10680 -75732 10688 -75688
rect 10780 -75732 10788 -75688
rect 11280 -75732 11288 -75688
rect 11380 -75732 11388 -75688
rect 11480 -75732 11488 -75688
rect 11580 -75732 11588 -75688
rect 11680 -75732 11688 -75688
rect 11780 -75732 11788 -75688
rect 11880 -75732 11888 -75688
rect 11980 -75732 11988 -75688
rect 12080 -75732 12088 -75688
rect 12180 -75732 12188 -75688
rect 12280 -75732 12288 -75688
rect 12380 -75732 12388 -75688
rect 12480 -75732 12488 -75688
rect 12580 -75732 12588 -75688
rect 12680 -75732 12688 -75688
rect 12780 -75732 12788 -75688
rect 13280 -75732 13288 -75688
rect 13380 -75732 13388 -75688
rect 13480 -75732 13488 -75688
rect 13580 -75732 13588 -75688
rect 13680 -75732 13688 -75688
rect 13780 -75732 13788 -75688
rect 13880 -75732 13888 -75688
rect 13980 -75732 13988 -75688
rect 14080 -75732 14088 -75688
rect 14180 -75732 14188 -75688
rect 14280 -75732 14288 -75688
rect 14380 -75732 14388 -75688
rect 14480 -75732 14488 -75688
rect 14580 -75732 14588 -75688
rect 14680 -75732 14688 -75688
rect 14780 -75732 14788 -75688
rect 15280 -75732 15288 -75688
rect 15380 -75732 15388 -75688
rect 15480 -75732 15488 -75688
rect 15580 -75732 15588 -75688
rect 15680 -75732 15688 -75688
rect 15780 -75732 15788 -75688
rect 15880 -75732 15888 -75688
rect 15980 -75732 15988 -75688
rect 16080 -75732 16088 -75688
rect 16180 -75732 16188 -75688
rect 16280 -75732 16288 -75688
rect 16380 -75732 16388 -75688
rect 16480 -75732 16488 -75688
rect 16580 -75732 16588 -75688
rect 16680 -75732 16688 -75688
rect 16780 -75732 16788 -75688
rect 9236 -75788 9280 -75780
rect 9336 -75788 9380 -75780
rect 9436 -75788 9480 -75780
rect 9536 -75788 9580 -75780
rect 9636 -75788 9680 -75780
rect 9736 -75788 9780 -75780
rect 9836 -75788 9880 -75780
rect 9936 -75788 9980 -75780
rect 10036 -75788 10080 -75780
rect 10136 -75788 10180 -75780
rect 10236 -75788 10280 -75780
rect 10336 -75788 10380 -75780
rect 10436 -75788 10480 -75780
rect 10536 -75788 10580 -75780
rect 10636 -75788 10680 -75780
rect 10736 -75788 10780 -75780
rect 11236 -75788 11280 -75780
rect 11336 -75788 11380 -75780
rect 11436 -75788 11480 -75780
rect 11536 -75788 11580 -75780
rect 11636 -75788 11680 -75780
rect 11736 -75788 11780 -75780
rect 11836 -75788 11880 -75780
rect 11936 -75788 11980 -75780
rect 12036 -75788 12080 -75780
rect 12136 -75788 12180 -75780
rect 12236 -75788 12280 -75780
rect 12336 -75788 12380 -75780
rect 12436 -75788 12480 -75780
rect 12536 -75788 12580 -75780
rect 12636 -75788 12680 -75780
rect 12736 -75788 12780 -75780
rect 13236 -75788 13280 -75780
rect 13336 -75788 13380 -75780
rect 13436 -75788 13480 -75780
rect 13536 -75788 13580 -75780
rect 13636 -75788 13680 -75780
rect 13736 -75788 13780 -75780
rect 13836 -75788 13880 -75780
rect 13936 -75788 13980 -75780
rect 14036 -75788 14080 -75780
rect 14136 -75788 14180 -75780
rect 14236 -75788 14280 -75780
rect 14336 -75788 14380 -75780
rect 14436 -75788 14480 -75780
rect 14536 -75788 14580 -75780
rect 14636 -75788 14680 -75780
rect 14736 -75788 14780 -75780
rect 15236 -75788 15280 -75780
rect 15336 -75788 15380 -75780
rect 15436 -75788 15480 -75780
rect 15536 -75788 15580 -75780
rect 15636 -75788 15680 -75780
rect 15736 -75788 15780 -75780
rect 15836 -75788 15880 -75780
rect 15936 -75788 15980 -75780
rect 16036 -75788 16080 -75780
rect 16136 -75788 16180 -75780
rect 16236 -75788 16280 -75780
rect 16336 -75788 16380 -75780
rect 16436 -75788 16480 -75780
rect 16536 -75788 16580 -75780
rect 16636 -75788 16680 -75780
rect 16736 -75788 16780 -75780
rect 9280 -75832 9288 -75788
rect 9380 -75832 9388 -75788
rect 9480 -75832 9488 -75788
rect 9580 -75832 9588 -75788
rect 9680 -75832 9688 -75788
rect 9780 -75832 9788 -75788
rect 9880 -75832 9888 -75788
rect 9980 -75832 9988 -75788
rect 10080 -75832 10088 -75788
rect 10180 -75832 10188 -75788
rect 10280 -75832 10288 -75788
rect 10380 -75832 10388 -75788
rect 10480 -75832 10488 -75788
rect 10580 -75832 10588 -75788
rect 10680 -75832 10688 -75788
rect 10780 -75832 10788 -75788
rect 11280 -75832 11288 -75788
rect 11380 -75832 11388 -75788
rect 11480 -75832 11488 -75788
rect 11580 -75832 11588 -75788
rect 11680 -75832 11688 -75788
rect 11780 -75832 11788 -75788
rect 11880 -75832 11888 -75788
rect 11980 -75832 11988 -75788
rect 12080 -75832 12088 -75788
rect 12180 -75832 12188 -75788
rect 12280 -75832 12288 -75788
rect 12380 -75832 12388 -75788
rect 12480 -75832 12488 -75788
rect 12580 -75832 12588 -75788
rect 12680 -75832 12688 -75788
rect 12780 -75832 12788 -75788
rect 13280 -75832 13288 -75788
rect 13380 -75832 13388 -75788
rect 13480 -75832 13488 -75788
rect 13580 -75832 13588 -75788
rect 13680 -75832 13688 -75788
rect 13780 -75832 13788 -75788
rect 13880 -75832 13888 -75788
rect 13980 -75832 13988 -75788
rect 14080 -75832 14088 -75788
rect 14180 -75832 14188 -75788
rect 14280 -75832 14288 -75788
rect 14380 -75832 14388 -75788
rect 14480 -75832 14488 -75788
rect 14580 -75832 14588 -75788
rect 14680 -75832 14688 -75788
rect 14780 -75832 14788 -75788
rect 15280 -75832 15288 -75788
rect 15380 -75832 15388 -75788
rect 15480 -75832 15488 -75788
rect 15580 -75832 15588 -75788
rect 15680 -75832 15688 -75788
rect 15780 -75832 15788 -75788
rect 15880 -75832 15888 -75788
rect 15980 -75832 15988 -75788
rect 16080 -75832 16088 -75788
rect 16180 -75832 16188 -75788
rect 16280 -75832 16288 -75788
rect 16380 -75832 16388 -75788
rect 16480 -75832 16488 -75788
rect 16580 -75832 16588 -75788
rect 16680 -75832 16688 -75788
rect 16780 -75832 16788 -75788
rect 9236 -75888 9280 -75880
rect 9336 -75888 9380 -75880
rect 9436 -75888 9480 -75880
rect 9536 -75888 9580 -75880
rect 9636 -75888 9680 -75880
rect 9736 -75888 9780 -75880
rect 9836 -75888 9880 -75880
rect 9936 -75888 9980 -75880
rect 10036 -75888 10080 -75880
rect 10136 -75888 10180 -75880
rect 10236 -75888 10280 -75880
rect 10336 -75888 10380 -75880
rect 10436 -75888 10480 -75880
rect 10536 -75888 10580 -75880
rect 10636 -75888 10680 -75880
rect 10736 -75888 10780 -75880
rect 11236 -75888 11280 -75880
rect 11336 -75888 11380 -75880
rect 11436 -75888 11480 -75880
rect 11536 -75888 11580 -75880
rect 11636 -75888 11680 -75880
rect 11736 -75888 11780 -75880
rect 11836 -75888 11880 -75880
rect 11936 -75888 11980 -75880
rect 12036 -75888 12080 -75880
rect 12136 -75888 12180 -75880
rect 12236 -75888 12280 -75880
rect 12336 -75888 12380 -75880
rect 12436 -75888 12480 -75880
rect 12536 -75888 12580 -75880
rect 12636 -75888 12680 -75880
rect 12736 -75888 12780 -75880
rect 13236 -75888 13280 -75880
rect 13336 -75888 13380 -75880
rect 13436 -75888 13480 -75880
rect 13536 -75888 13580 -75880
rect 13636 -75888 13680 -75880
rect 13736 -75888 13780 -75880
rect 13836 -75888 13880 -75880
rect 13936 -75888 13980 -75880
rect 14036 -75888 14080 -75880
rect 14136 -75888 14180 -75880
rect 14236 -75888 14280 -75880
rect 14336 -75888 14380 -75880
rect 14436 -75888 14480 -75880
rect 14536 -75888 14580 -75880
rect 14636 -75888 14680 -75880
rect 14736 -75888 14780 -75880
rect 15236 -75888 15280 -75880
rect 15336 -75888 15380 -75880
rect 15436 -75888 15480 -75880
rect 15536 -75888 15580 -75880
rect 15636 -75888 15680 -75880
rect 15736 -75888 15780 -75880
rect 15836 -75888 15880 -75880
rect 15936 -75888 15980 -75880
rect 16036 -75888 16080 -75880
rect 16136 -75888 16180 -75880
rect 16236 -75888 16280 -75880
rect 16336 -75888 16380 -75880
rect 16436 -75888 16480 -75880
rect 16536 -75888 16580 -75880
rect 16636 -75888 16680 -75880
rect 16736 -75888 16780 -75880
rect 9280 -75932 9288 -75888
rect 9380 -75932 9388 -75888
rect 9480 -75932 9488 -75888
rect 9580 -75932 9588 -75888
rect 9680 -75932 9688 -75888
rect 9780 -75932 9788 -75888
rect 9880 -75932 9888 -75888
rect 9980 -75932 9988 -75888
rect 10080 -75932 10088 -75888
rect 10180 -75932 10188 -75888
rect 10280 -75932 10288 -75888
rect 10380 -75932 10388 -75888
rect 10480 -75932 10488 -75888
rect 10580 -75932 10588 -75888
rect 10680 -75932 10688 -75888
rect 10780 -75932 10788 -75888
rect 11280 -75932 11288 -75888
rect 11380 -75932 11388 -75888
rect 11480 -75932 11488 -75888
rect 11580 -75932 11588 -75888
rect 11680 -75932 11688 -75888
rect 11780 -75932 11788 -75888
rect 11880 -75932 11888 -75888
rect 11980 -75932 11988 -75888
rect 12080 -75932 12088 -75888
rect 12180 -75932 12188 -75888
rect 12280 -75932 12288 -75888
rect 12380 -75932 12388 -75888
rect 12480 -75932 12488 -75888
rect 12580 -75932 12588 -75888
rect 12680 -75932 12688 -75888
rect 12780 -75932 12788 -75888
rect 13280 -75932 13288 -75888
rect 13380 -75932 13388 -75888
rect 13480 -75932 13488 -75888
rect 13580 -75932 13588 -75888
rect 13680 -75932 13688 -75888
rect 13780 -75932 13788 -75888
rect 13880 -75932 13888 -75888
rect 13980 -75932 13988 -75888
rect 14080 -75932 14088 -75888
rect 14180 -75932 14188 -75888
rect 14280 -75932 14288 -75888
rect 14380 -75932 14388 -75888
rect 14480 -75932 14488 -75888
rect 14580 -75932 14588 -75888
rect 14680 -75932 14688 -75888
rect 14780 -75932 14788 -75888
rect 15280 -75932 15288 -75888
rect 15380 -75932 15388 -75888
rect 15480 -75932 15488 -75888
rect 15580 -75932 15588 -75888
rect 15680 -75932 15688 -75888
rect 15780 -75932 15788 -75888
rect 15880 -75932 15888 -75888
rect 15980 -75932 15988 -75888
rect 16080 -75932 16088 -75888
rect 16180 -75932 16188 -75888
rect 16280 -75932 16288 -75888
rect 16380 -75932 16388 -75888
rect 16480 -75932 16488 -75888
rect 16580 -75932 16588 -75888
rect 16680 -75932 16688 -75888
rect 16780 -75932 16788 -75888
rect 9236 -75988 9280 -75980
rect 9336 -75988 9380 -75980
rect 9436 -75988 9480 -75980
rect 9536 -75988 9580 -75980
rect 9636 -75988 9680 -75980
rect 9736 -75988 9780 -75980
rect 9836 -75988 9880 -75980
rect 9936 -75988 9980 -75980
rect 10036 -75988 10080 -75980
rect 10136 -75988 10180 -75980
rect 10236 -75988 10280 -75980
rect 10336 -75988 10380 -75980
rect 10436 -75988 10480 -75980
rect 10536 -75988 10580 -75980
rect 10636 -75988 10680 -75980
rect 10736 -75988 10780 -75980
rect 11236 -75988 11280 -75980
rect 11336 -75988 11380 -75980
rect 11436 -75988 11480 -75980
rect 11536 -75988 11580 -75980
rect 11636 -75988 11680 -75980
rect 11736 -75988 11780 -75980
rect 11836 -75988 11880 -75980
rect 11936 -75988 11980 -75980
rect 12036 -75988 12080 -75980
rect 12136 -75988 12180 -75980
rect 12236 -75988 12280 -75980
rect 12336 -75988 12380 -75980
rect 12436 -75988 12480 -75980
rect 12536 -75988 12580 -75980
rect 12636 -75988 12680 -75980
rect 12736 -75988 12780 -75980
rect 13236 -75988 13280 -75980
rect 13336 -75988 13380 -75980
rect 13436 -75988 13480 -75980
rect 13536 -75988 13580 -75980
rect 13636 -75988 13680 -75980
rect 13736 -75988 13780 -75980
rect 13836 -75988 13880 -75980
rect 13936 -75988 13980 -75980
rect 14036 -75988 14080 -75980
rect 14136 -75988 14180 -75980
rect 14236 -75988 14280 -75980
rect 14336 -75988 14380 -75980
rect 14436 -75988 14480 -75980
rect 14536 -75988 14580 -75980
rect 14636 -75988 14680 -75980
rect 14736 -75988 14780 -75980
rect 15236 -75988 15280 -75980
rect 15336 -75988 15380 -75980
rect 15436 -75988 15480 -75980
rect 15536 -75988 15580 -75980
rect 15636 -75988 15680 -75980
rect 15736 -75988 15780 -75980
rect 15836 -75988 15880 -75980
rect 15936 -75988 15980 -75980
rect 16036 -75988 16080 -75980
rect 16136 -75988 16180 -75980
rect 16236 -75988 16280 -75980
rect 16336 -75988 16380 -75980
rect 16436 -75988 16480 -75980
rect 16536 -75988 16580 -75980
rect 16636 -75988 16680 -75980
rect 16736 -75988 16780 -75980
rect 9280 -76032 9288 -75988
rect 9380 -76032 9388 -75988
rect 9480 -76032 9488 -75988
rect 9580 -76032 9588 -75988
rect 9680 -76032 9688 -75988
rect 9780 -76032 9788 -75988
rect 9880 -76032 9888 -75988
rect 9980 -76032 9988 -75988
rect 10080 -76032 10088 -75988
rect 10180 -76032 10188 -75988
rect 10280 -76032 10288 -75988
rect 10380 -76032 10388 -75988
rect 10480 -76032 10488 -75988
rect 10580 -76032 10588 -75988
rect 10680 -76032 10688 -75988
rect 10780 -76032 10788 -75988
rect 11280 -76032 11288 -75988
rect 11380 -76032 11388 -75988
rect 11480 -76032 11488 -75988
rect 11580 -76032 11588 -75988
rect 11680 -76032 11688 -75988
rect 11780 -76032 11788 -75988
rect 11880 -76032 11888 -75988
rect 11980 -76032 11988 -75988
rect 12080 -76032 12088 -75988
rect 12180 -76032 12188 -75988
rect 12280 -76032 12288 -75988
rect 12380 -76032 12388 -75988
rect 12480 -76032 12488 -75988
rect 12580 -76032 12588 -75988
rect 12680 -76032 12688 -75988
rect 12780 -76032 12788 -75988
rect 13280 -76032 13288 -75988
rect 13380 -76032 13388 -75988
rect 13480 -76032 13488 -75988
rect 13580 -76032 13588 -75988
rect 13680 -76032 13688 -75988
rect 13780 -76032 13788 -75988
rect 13880 -76032 13888 -75988
rect 13980 -76032 13988 -75988
rect 14080 -76032 14088 -75988
rect 14180 -76032 14188 -75988
rect 14280 -76032 14288 -75988
rect 14380 -76032 14388 -75988
rect 14480 -76032 14488 -75988
rect 14580 -76032 14588 -75988
rect 14680 -76032 14688 -75988
rect 14780 -76032 14788 -75988
rect 15280 -76032 15288 -75988
rect 15380 -76032 15388 -75988
rect 15480 -76032 15488 -75988
rect 15580 -76032 15588 -75988
rect 15680 -76032 15688 -75988
rect 15780 -76032 15788 -75988
rect 15880 -76032 15888 -75988
rect 15980 -76032 15988 -75988
rect 16080 -76032 16088 -75988
rect 16180 -76032 16188 -75988
rect 16280 -76032 16288 -75988
rect 16380 -76032 16388 -75988
rect 16480 -76032 16488 -75988
rect 16580 -76032 16588 -75988
rect 16680 -76032 16688 -75988
rect 16780 -76032 16788 -75988
rect 9236 -76088 9280 -76080
rect 9336 -76088 9380 -76080
rect 9436 -76088 9480 -76080
rect 9536 -76088 9580 -76080
rect 9636 -76088 9680 -76080
rect 9736 -76088 9780 -76080
rect 9836 -76088 9880 -76080
rect 9936 -76088 9980 -76080
rect 10036 -76088 10080 -76080
rect 10136 -76088 10180 -76080
rect 10236 -76088 10280 -76080
rect 10336 -76088 10380 -76080
rect 10436 -76088 10480 -76080
rect 10536 -76088 10580 -76080
rect 10636 -76088 10680 -76080
rect 10736 -76088 10780 -76080
rect 11236 -76088 11280 -76080
rect 11336 -76088 11380 -76080
rect 11436 -76088 11480 -76080
rect 11536 -76088 11580 -76080
rect 11636 -76088 11680 -76080
rect 11736 -76088 11780 -76080
rect 11836 -76088 11880 -76080
rect 11936 -76088 11980 -76080
rect 12036 -76088 12080 -76080
rect 12136 -76088 12180 -76080
rect 12236 -76088 12280 -76080
rect 12336 -76088 12380 -76080
rect 12436 -76088 12480 -76080
rect 12536 -76088 12580 -76080
rect 12636 -76088 12680 -76080
rect 12736 -76088 12780 -76080
rect 13236 -76088 13280 -76080
rect 13336 -76088 13380 -76080
rect 13436 -76088 13480 -76080
rect 13536 -76088 13580 -76080
rect 13636 -76088 13680 -76080
rect 13736 -76088 13780 -76080
rect 13836 -76088 13880 -76080
rect 13936 -76088 13980 -76080
rect 14036 -76088 14080 -76080
rect 14136 -76088 14180 -76080
rect 14236 -76088 14280 -76080
rect 14336 -76088 14380 -76080
rect 14436 -76088 14480 -76080
rect 14536 -76088 14580 -76080
rect 14636 -76088 14680 -76080
rect 14736 -76088 14780 -76080
rect 15236 -76088 15280 -76080
rect 15336 -76088 15380 -76080
rect 15436 -76088 15480 -76080
rect 15536 -76088 15580 -76080
rect 15636 -76088 15680 -76080
rect 15736 -76088 15780 -76080
rect 15836 -76088 15880 -76080
rect 15936 -76088 15980 -76080
rect 16036 -76088 16080 -76080
rect 16136 -76088 16180 -76080
rect 16236 -76088 16280 -76080
rect 16336 -76088 16380 -76080
rect 16436 -76088 16480 -76080
rect 16536 -76088 16580 -76080
rect 16636 -76088 16680 -76080
rect 16736 -76088 16780 -76080
rect 9280 -76132 9288 -76088
rect 9380 -76132 9388 -76088
rect 9480 -76132 9488 -76088
rect 9580 -76132 9588 -76088
rect 9680 -76132 9688 -76088
rect 9780 -76132 9788 -76088
rect 9880 -76132 9888 -76088
rect 9980 -76132 9988 -76088
rect 10080 -76132 10088 -76088
rect 10180 -76132 10188 -76088
rect 10280 -76132 10288 -76088
rect 10380 -76132 10388 -76088
rect 10480 -76132 10488 -76088
rect 10580 -76132 10588 -76088
rect 10680 -76132 10688 -76088
rect 10780 -76132 10788 -76088
rect 11280 -76132 11288 -76088
rect 11380 -76132 11388 -76088
rect 11480 -76132 11488 -76088
rect 11580 -76132 11588 -76088
rect 11680 -76132 11688 -76088
rect 11780 -76132 11788 -76088
rect 11880 -76132 11888 -76088
rect 11980 -76132 11988 -76088
rect 12080 -76132 12088 -76088
rect 12180 -76132 12188 -76088
rect 12280 -76132 12288 -76088
rect 12380 -76132 12388 -76088
rect 12480 -76132 12488 -76088
rect 12580 -76132 12588 -76088
rect 12680 -76132 12688 -76088
rect 12780 -76132 12788 -76088
rect 13280 -76132 13288 -76088
rect 13380 -76132 13388 -76088
rect 13480 -76132 13488 -76088
rect 13580 -76132 13588 -76088
rect 13680 -76132 13688 -76088
rect 13780 -76132 13788 -76088
rect 13880 -76132 13888 -76088
rect 13980 -76132 13988 -76088
rect 14080 -76132 14088 -76088
rect 14180 -76132 14188 -76088
rect 14280 -76132 14288 -76088
rect 14380 -76132 14388 -76088
rect 14480 -76132 14488 -76088
rect 14580 -76132 14588 -76088
rect 14680 -76132 14688 -76088
rect 14780 -76132 14788 -76088
rect 15280 -76132 15288 -76088
rect 15380 -76132 15388 -76088
rect 15480 -76132 15488 -76088
rect 15580 -76132 15588 -76088
rect 15680 -76132 15688 -76088
rect 15780 -76132 15788 -76088
rect 15880 -76132 15888 -76088
rect 15980 -76132 15988 -76088
rect 16080 -76132 16088 -76088
rect 16180 -76132 16188 -76088
rect 16280 -76132 16288 -76088
rect 16380 -76132 16388 -76088
rect 16480 -76132 16488 -76088
rect 16580 -76132 16588 -76088
rect 16680 -76132 16688 -76088
rect 16780 -76132 16788 -76088
rect 9236 -76188 9280 -76180
rect 9336 -76188 9380 -76180
rect 9436 -76188 9480 -76180
rect 9536 -76188 9580 -76180
rect 9636 -76188 9680 -76180
rect 9736 -76188 9780 -76180
rect 9836 -76188 9880 -76180
rect 9936 -76188 9980 -76180
rect 10036 -76188 10080 -76180
rect 10136 -76188 10180 -76180
rect 10236 -76188 10280 -76180
rect 10336 -76188 10380 -76180
rect 10436 -76188 10480 -76180
rect 10536 -76188 10580 -76180
rect 10636 -76188 10680 -76180
rect 10736 -76188 10780 -76180
rect 11236 -76188 11280 -76180
rect 11336 -76188 11380 -76180
rect 11436 -76188 11480 -76180
rect 11536 -76188 11580 -76180
rect 11636 -76188 11680 -76180
rect 11736 -76188 11780 -76180
rect 11836 -76188 11880 -76180
rect 11936 -76188 11980 -76180
rect 12036 -76188 12080 -76180
rect 12136 -76188 12180 -76180
rect 12236 -76188 12280 -76180
rect 12336 -76188 12380 -76180
rect 12436 -76188 12480 -76180
rect 12536 -76188 12580 -76180
rect 12636 -76188 12680 -76180
rect 12736 -76188 12780 -76180
rect 13236 -76188 13280 -76180
rect 13336 -76188 13380 -76180
rect 13436 -76188 13480 -76180
rect 13536 -76188 13580 -76180
rect 13636 -76188 13680 -76180
rect 13736 -76188 13780 -76180
rect 13836 -76188 13880 -76180
rect 13936 -76188 13980 -76180
rect 14036 -76188 14080 -76180
rect 14136 -76188 14180 -76180
rect 14236 -76188 14280 -76180
rect 14336 -76188 14380 -76180
rect 14436 -76188 14480 -76180
rect 14536 -76188 14580 -76180
rect 14636 -76188 14680 -76180
rect 14736 -76188 14780 -76180
rect 15236 -76188 15280 -76180
rect 15336 -76188 15380 -76180
rect 15436 -76188 15480 -76180
rect 15536 -76188 15580 -76180
rect 15636 -76188 15680 -76180
rect 15736 -76188 15780 -76180
rect 15836 -76188 15880 -76180
rect 15936 -76188 15980 -76180
rect 16036 -76188 16080 -76180
rect 16136 -76188 16180 -76180
rect 16236 -76188 16280 -76180
rect 16336 -76188 16380 -76180
rect 16436 -76188 16480 -76180
rect 16536 -76188 16580 -76180
rect 16636 -76188 16680 -76180
rect 16736 -76188 16780 -76180
rect 9280 -76232 9288 -76188
rect 9380 -76232 9388 -76188
rect 9480 -76232 9488 -76188
rect 9580 -76232 9588 -76188
rect 9680 -76232 9688 -76188
rect 9780 -76232 9788 -76188
rect 9880 -76232 9888 -76188
rect 9980 -76232 9988 -76188
rect 10080 -76232 10088 -76188
rect 10180 -76232 10188 -76188
rect 10280 -76232 10288 -76188
rect 10380 -76232 10388 -76188
rect 10480 -76232 10488 -76188
rect 10580 -76232 10588 -76188
rect 10680 -76232 10688 -76188
rect 10780 -76232 10788 -76188
rect 11280 -76232 11288 -76188
rect 11380 -76232 11388 -76188
rect 11480 -76232 11488 -76188
rect 11580 -76232 11588 -76188
rect 11680 -76232 11688 -76188
rect 11780 -76232 11788 -76188
rect 11880 -76232 11888 -76188
rect 11980 -76232 11988 -76188
rect 12080 -76232 12088 -76188
rect 12180 -76232 12188 -76188
rect 12280 -76232 12288 -76188
rect 12380 -76232 12388 -76188
rect 12480 -76232 12488 -76188
rect 12580 -76232 12588 -76188
rect 12680 -76232 12688 -76188
rect 12780 -76232 12788 -76188
rect 13280 -76232 13288 -76188
rect 13380 -76232 13388 -76188
rect 13480 -76232 13488 -76188
rect 13580 -76232 13588 -76188
rect 13680 -76232 13688 -76188
rect 13780 -76232 13788 -76188
rect 13880 -76232 13888 -76188
rect 13980 -76232 13988 -76188
rect 14080 -76232 14088 -76188
rect 14180 -76232 14188 -76188
rect 14280 -76232 14288 -76188
rect 14380 -76232 14388 -76188
rect 14480 -76232 14488 -76188
rect 14580 -76232 14588 -76188
rect 14680 -76232 14688 -76188
rect 14780 -76232 14788 -76188
rect 15280 -76232 15288 -76188
rect 15380 -76232 15388 -76188
rect 15480 -76232 15488 -76188
rect 15580 -76232 15588 -76188
rect 15680 -76232 15688 -76188
rect 15780 -76232 15788 -76188
rect 15880 -76232 15888 -76188
rect 15980 -76232 15988 -76188
rect 16080 -76232 16088 -76188
rect 16180 -76232 16188 -76188
rect 16280 -76232 16288 -76188
rect 16380 -76232 16388 -76188
rect 16480 -76232 16488 -76188
rect 16580 -76232 16588 -76188
rect 16680 -76232 16688 -76188
rect 16780 -76232 16788 -76188
rect 9236 -76288 9280 -76280
rect 9336 -76288 9380 -76280
rect 9436 -76288 9480 -76280
rect 9536 -76288 9580 -76280
rect 9636 -76288 9680 -76280
rect 9736 -76288 9780 -76280
rect 9836 -76288 9880 -76280
rect 9936 -76288 9980 -76280
rect 10036 -76288 10080 -76280
rect 10136 -76288 10180 -76280
rect 10236 -76288 10280 -76280
rect 10336 -76288 10380 -76280
rect 10436 -76288 10480 -76280
rect 10536 -76288 10580 -76280
rect 10636 -76288 10680 -76280
rect 10736 -76288 10780 -76280
rect 11236 -76288 11280 -76280
rect 11336 -76288 11380 -76280
rect 11436 -76288 11480 -76280
rect 11536 -76288 11580 -76280
rect 11636 -76288 11680 -76280
rect 11736 -76288 11780 -76280
rect 11836 -76288 11880 -76280
rect 11936 -76288 11980 -76280
rect 12036 -76288 12080 -76280
rect 12136 -76288 12180 -76280
rect 12236 -76288 12280 -76280
rect 12336 -76288 12380 -76280
rect 12436 -76288 12480 -76280
rect 12536 -76288 12580 -76280
rect 12636 -76288 12680 -76280
rect 12736 -76288 12780 -76280
rect 13236 -76288 13280 -76280
rect 13336 -76288 13380 -76280
rect 13436 -76288 13480 -76280
rect 13536 -76288 13580 -76280
rect 13636 -76288 13680 -76280
rect 13736 -76288 13780 -76280
rect 13836 -76288 13880 -76280
rect 13936 -76288 13980 -76280
rect 14036 -76288 14080 -76280
rect 14136 -76288 14180 -76280
rect 14236 -76288 14280 -76280
rect 14336 -76288 14380 -76280
rect 14436 -76288 14480 -76280
rect 14536 -76288 14580 -76280
rect 14636 -76288 14680 -76280
rect 14736 -76288 14780 -76280
rect 15236 -76288 15280 -76280
rect 15336 -76288 15380 -76280
rect 15436 -76288 15480 -76280
rect 15536 -76288 15580 -76280
rect 15636 -76288 15680 -76280
rect 15736 -76288 15780 -76280
rect 15836 -76288 15880 -76280
rect 15936 -76288 15980 -76280
rect 16036 -76288 16080 -76280
rect 16136 -76288 16180 -76280
rect 16236 -76288 16280 -76280
rect 16336 -76288 16380 -76280
rect 16436 -76288 16480 -76280
rect 16536 -76288 16580 -76280
rect 16636 -76288 16680 -76280
rect 16736 -76288 16780 -76280
rect 9280 -76332 9288 -76288
rect 9380 -76332 9388 -76288
rect 9480 -76332 9488 -76288
rect 9580 -76332 9588 -76288
rect 9680 -76332 9688 -76288
rect 9780 -76332 9788 -76288
rect 9880 -76332 9888 -76288
rect 9980 -76332 9988 -76288
rect 10080 -76332 10088 -76288
rect 10180 -76332 10188 -76288
rect 10280 -76332 10288 -76288
rect 10380 -76332 10388 -76288
rect 10480 -76332 10488 -76288
rect 10580 -76332 10588 -76288
rect 10680 -76332 10688 -76288
rect 10780 -76332 10788 -76288
rect 11280 -76332 11288 -76288
rect 11380 -76332 11388 -76288
rect 11480 -76332 11488 -76288
rect 11580 -76332 11588 -76288
rect 11680 -76332 11688 -76288
rect 11780 -76332 11788 -76288
rect 11880 -76332 11888 -76288
rect 11980 -76332 11988 -76288
rect 12080 -76332 12088 -76288
rect 12180 -76332 12188 -76288
rect 12280 -76332 12288 -76288
rect 12380 -76332 12388 -76288
rect 12480 -76332 12488 -76288
rect 12580 -76332 12588 -76288
rect 12680 -76332 12688 -76288
rect 12780 -76332 12788 -76288
rect 13280 -76332 13288 -76288
rect 13380 -76332 13388 -76288
rect 13480 -76332 13488 -76288
rect 13580 -76332 13588 -76288
rect 13680 -76332 13688 -76288
rect 13780 -76332 13788 -76288
rect 13880 -76332 13888 -76288
rect 13980 -76332 13988 -76288
rect 14080 -76332 14088 -76288
rect 14180 -76332 14188 -76288
rect 14280 -76332 14288 -76288
rect 14380 -76332 14388 -76288
rect 14480 -76332 14488 -76288
rect 14580 -76332 14588 -76288
rect 14680 -76332 14688 -76288
rect 14780 -76332 14788 -76288
rect 15280 -76332 15288 -76288
rect 15380 -76332 15388 -76288
rect 15480 -76332 15488 -76288
rect 15580 -76332 15588 -76288
rect 15680 -76332 15688 -76288
rect 15780 -76332 15788 -76288
rect 15880 -76332 15888 -76288
rect 15980 -76332 15988 -76288
rect 16080 -76332 16088 -76288
rect 16180 -76332 16188 -76288
rect 16280 -76332 16288 -76288
rect 16380 -76332 16388 -76288
rect 16480 -76332 16488 -76288
rect 16580 -76332 16588 -76288
rect 16680 -76332 16688 -76288
rect 16780 -76332 16788 -76288
rect 9236 -76388 9280 -76380
rect 9336 -76388 9380 -76380
rect 9436 -76388 9480 -76380
rect 9536 -76388 9580 -76380
rect 9636 -76388 9680 -76380
rect 9736 -76388 9780 -76380
rect 9836 -76388 9880 -76380
rect 9936 -76388 9980 -76380
rect 10036 -76388 10080 -76380
rect 10136 -76388 10180 -76380
rect 10236 -76388 10280 -76380
rect 10336 -76388 10380 -76380
rect 10436 -76388 10480 -76380
rect 10536 -76388 10580 -76380
rect 10636 -76388 10680 -76380
rect 10736 -76388 10780 -76380
rect 11236 -76388 11280 -76380
rect 11336 -76388 11380 -76380
rect 11436 -76388 11480 -76380
rect 11536 -76388 11580 -76380
rect 11636 -76388 11680 -76380
rect 11736 -76388 11780 -76380
rect 11836 -76388 11880 -76380
rect 11936 -76388 11980 -76380
rect 12036 -76388 12080 -76380
rect 12136 -76388 12180 -76380
rect 12236 -76388 12280 -76380
rect 12336 -76388 12380 -76380
rect 12436 -76388 12480 -76380
rect 12536 -76388 12580 -76380
rect 12636 -76388 12680 -76380
rect 12736 -76388 12780 -76380
rect 13236 -76388 13280 -76380
rect 13336 -76388 13380 -76380
rect 13436 -76388 13480 -76380
rect 13536 -76388 13580 -76380
rect 13636 -76388 13680 -76380
rect 13736 -76388 13780 -76380
rect 13836 -76388 13880 -76380
rect 13936 -76388 13980 -76380
rect 14036 -76388 14080 -76380
rect 14136 -76388 14180 -76380
rect 14236 -76388 14280 -76380
rect 14336 -76388 14380 -76380
rect 14436 -76388 14480 -76380
rect 14536 -76388 14580 -76380
rect 14636 -76388 14680 -76380
rect 14736 -76388 14780 -76380
rect 15236 -76388 15280 -76380
rect 15336 -76388 15380 -76380
rect 15436 -76388 15480 -76380
rect 15536 -76388 15580 -76380
rect 15636 -76388 15680 -76380
rect 15736 -76388 15780 -76380
rect 15836 -76388 15880 -76380
rect 15936 -76388 15980 -76380
rect 16036 -76388 16080 -76380
rect 16136 -76388 16180 -76380
rect 16236 -76388 16280 -76380
rect 16336 -76388 16380 -76380
rect 16436 -76388 16480 -76380
rect 16536 -76388 16580 -76380
rect 16636 -76388 16680 -76380
rect 16736 -76388 16780 -76380
rect 9280 -76432 9288 -76388
rect 9380 -76432 9388 -76388
rect 9480 -76432 9488 -76388
rect 9580 -76432 9588 -76388
rect 9680 -76432 9688 -76388
rect 9780 -76432 9788 -76388
rect 9880 -76432 9888 -76388
rect 9980 -76432 9988 -76388
rect 10080 -76432 10088 -76388
rect 10180 -76432 10188 -76388
rect 10280 -76432 10288 -76388
rect 10380 -76432 10388 -76388
rect 10480 -76432 10488 -76388
rect 10580 -76432 10588 -76388
rect 10680 -76432 10688 -76388
rect 10780 -76432 10788 -76388
rect 11280 -76432 11288 -76388
rect 11380 -76432 11388 -76388
rect 11480 -76432 11488 -76388
rect 11580 -76432 11588 -76388
rect 11680 -76432 11688 -76388
rect 11780 -76432 11788 -76388
rect 11880 -76432 11888 -76388
rect 11980 -76432 11988 -76388
rect 12080 -76432 12088 -76388
rect 12180 -76432 12188 -76388
rect 12280 -76432 12288 -76388
rect 12380 -76432 12388 -76388
rect 12480 -76432 12488 -76388
rect 12580 -76432 12588 -76388
rect 12680 -76432 12688 -76388
rect 12780 -76432 12788 -76388
rect 13280 -76432 13288 -76388
rect 13380 -76432 13388 -76388
rect 13480 -76432 13488 -76388
rect 13580 -76432 13588 -76388
rect 13680 -76432 13688 -76388
rect 13780 -76432 13788 -76388
rect 13880 -76432 13888 -76388
rect 13980 -76432 13988 -76388
rect 14080 -76432 14088 -76388
rect 14180 -76432 14188 -76388
rect 14280 -76432 14288 -76388
rect 14380 -76432 14388 -76388
rect 14480 -76432 14488 -76388
rect 14580 -76432 14588 -76388
rect 14680 -76432 14688 -76388
rect 14780 -76432 14788 -76388
rect 15280 -76432 15288 -76388
rect 15380 -76432 15388 -76388
rect 15480 -76432 15488 -76388
rect 15580 -76432 15588 -76388
rect 15680 -76432 15688 -76388
rect 15780 -76432 15788 -76388
rect 15880 -76432 15888 -76388
rect 15980 -76432 15988 -76388
rect 16080 -76432 16088 -76388
rect 16180 -76432 16188 -76388
rect 16280 -76432 16288 -76388
rect 16380 -76432 16388 -76388
rect 16480 -76432 16488 -76388
rect 16580 -76432 16588 -76388
rect 16680 -76432 16688 -76388
rect 16780 -76432 16788 -76388
rect 9236 -76488 9280 -76480
rect 9336 -76488 9380 -76480
rect 9436 -76488 9480 -76480
rect 9536 -76488 9580 -76480
rect 9636 -76488 9680 -76480
rect 9736 -76488 9780 -76480
rect 9836 -76488 9880 -76480
rect 9936 -76488 9980 -76480
rect 10036 -76488 10080 -76480
rect 10136 -76488 10180 -76480
rect 10236 -76488 10280 -76480
rect 10336 -76488 10380 -76480
rect 10436 -76488 10480 -76480
rect 10536 -76488 10580 -76480
rect 10636 -76488 10680 -76480
rect 10736 -76488 10780 -76480
rect 11236 -76488 11280 -76480
rect 11336 -76488 11380 -76480
rect 11436 -76488 11480 -76480
rect 11536 -76488 11580 -76480
rect 11636 -76488 11680 -76480
rect 11736 -76488 11780 -76480
rect 11836 -76488 11880 -76480
rect 11936 -76488 11980 -76480
rect 12036 -76488 12080 -76480
rect 12136 -76488 12180 -76480
rect 12236 -76488 12280 -76480
rect 12336 -76488 12380 -76480
rect 12436 -76488 12480 -76480
rect 12536 -76488 12580 -76480
rect 12636 -76488 12680 -76480
rect 12736 -76488 12780 -76480
rect 13236 -76488 13280 -76480
rect 13336 -76488 13380 -76480
rect 13436 -76488 13480 -76480
rect 13536 -76488 13580 -76480
rect 13636 -76488 13680 -76480
rect 13736 -76488 13780 -76480
rect 13836 -76488 13880 -76480
rect 13936 -76488 13980 -76480
rect 14036 -76488 14080 -76480
rect 14136 -76488 14180 -76480
rect 14236 -76488 14280 -76480
rect 14336 -76488 14380 -76480
rect 14436 -76488 14480 -76480
rect 14536 -76488 14580 -76480
rect 14636 -76488 14680 -76480
rect 14736 -76488 14780 -76480
rect 15236 -76488 15280 -76480
rect 15336 -76488 15380 -76480
rect 15436 -76488 15480 -76480
rect 15536 -76488 15580 -76480
rect 15636 -76488 15680 -76480
rect 15736 -76488 15780 -76480
rect 15836 -76488 15880 -76480
rect 15936 -76488 15980 -76480
rect 16036 -76488 16080 -76480
rect 16136 -76488 16180 -76480
rect 16236 -76488 16280 -76480
rect 16336 -76488 16380 -76480
rect 16436 -76488 16480 -76480
rect 16536 -76488 16580 -76480
rect 16636 -76488 16680 -76480
rect 16736 -76488 16780 -76480
rect 9280 -76532 9288 -76488
rect 9380 -76532 9388 -76488
rect 9480 -76532 9488 -76488
rect 9580 -76532 9588 -76488
rect 9680 -76532 9688 -76488
rect 9780 -76532 9788 -76488
rect 9880 -76532 9888 -76488
rect 9980 -76532 9988 -76488
rect 10080 -76532 10088 -76488
rect 10180 -76532 10188 -76488
rect 10280 -76532 10288 -76488
rect 10380 -76532 10388 -76488
rect 10480 -76532 10488 -76488
rect 10580 -76532 10588 -76488
rect 10680 -76532 10688 -76488
rect 10780 -76532 10788 -76488
rect 11280 -76532 11288 -76488
rect 11380 -76532 11388 -76488
rect 11480 -76532 11488 -76488
rect 11580 -76532 11588 -76488
rect 11680 -76532 11688 -76488
rect 11780 -76532 11788 -76488
rect 11880 -76532 11888 -76488
rect 11980 -76532 11988 -76488
rect 12080 -76532 12088 -76488
rect 12180 -76532 12188 -76488
rect 12280 -76532 12288 -76488
rect 12380 -76532 12388 -76488
rect 12480 -76532 12488 -76488
rect 12580 -76532 12588 -76488
rect 12680 -76532 12688 -76488
rect 12780 -76532 12788 -76488
rect 13280 -76532 13288 -76488
rect 13380 -76532 13388 -76488
rect 13480 -76532 13488 -76488
rect 13580 -76532 13588 -76488
rect 13680 -76532 13688 -76488
rect 13780 -76532 13788 -76488
rect 13880 -76532 13888 -76488
rect 13980 -76532 13988 -76488
rect 14080 -76532 14088 -76488
rect 14180 -76532 14188 -76488
rect 14280 -76532 14288 -76488
rect 14380 -76532 14388 -76488
rect 14480 -76532 14488 -76488
rect 14580 -76532 14588 -76488
rect 14680 -76532 14688 -76488
rect 14780 -76532 14788 -76488
rect 15280 -76532 15288 -76488
rect 15380 -76532 15388 -76488
rect 15480 -76532 15488 -76488
rect 15580 -76532 15588 -76488
rect 15680 -76532 15688 -76488
rect 15780 -76532 15788 -76488
rect 15880 -76532 15888 -76488
rect 15980 -76532 15988 -76488
rect 16080 -76532 16088 -76488
rect 16180 -76532 16188 -76488
rect 16280 -76532 16288 -76488
rect 16380 -76532 16388 -76488
rect 16480 -76532 16488 -76488
rect 16580 -76532 16588 -76488
rect 16680 -76532 16688 -76488
rect 16780 -76532 16788 -76488
rect 9236 -76588 9280 -76580
rect 9336 -76588 9380 -76580
rect 9436 -76588 9480 -76580
rect 9536 -76588 9580 -76580
rect 9636 -76588 9680 -76580
rect 9736 -76588 9780 -76580
rect 9836 -76588 9880 -76580
rect 9936 -76588 9980 -76580
rect 10036 -76588 10080 -76580
rect 10136 -76588 10180 -76580
rect 10236 -76588 10280 -76580
rect 10336 -76588 10380 -76580
rect 10436 -76588 10480 -76580
rect 10536 -76588 10580 -76580
rect 10636 -76588 10680 -76580
rect 10736 -76588 10780 -76580
rect 11236 -76588 11280 -76580
rect 11336 -76588 11380 -76580
rect 11436 -76588 11480 -76580
rect 11536 -76588 11580 -76580
rect 11636 -76588 11680 -76580
rect 11736 -76588 11780 -76580
rect 11836 -76588 11880 -76580
rect 11936 -76588 11980 -76580
rect 12036 -76588 12080 -76580
rect 12136 -76588 12180 -76580
rect 12236 -76588 12280 -76580
rect 12336 -76588 12380 -76580
rect 12436 -76588 12480 -76580
rect 12536 -76588 12580 -76580
rect 12636 -76588 12680 -76580
rect 12736 -76588 12780 -76580
rect 13236 -76588 13280 -76580
rect 13336 -76588 13380 -76580
rect 13436 -76588 13480 -76580
rect 13536 -76588 13580 -76580
rect 13636 -76588 13680 -76580
rect 13736 -76588 13780 -76580
rect 13836 -76588 13880 -76580
rect 13936 -76588 13980 -76580
rect 14036 -76588 14080 -76580
rect 14136 -76588 14180 -76580
rect 14236 -76588 14280 -76580
rect 14336 -76588 14380 -76580
rect 14436 -76588 14480 -76580
rect 14536 -76588 14580 -76580
rect 14636 -76588 14680 -76580
rect 14736 -76588 14780 -76580
rect 15236 -76588 15280 -76580
rect 15336 -76588 15380 -76580
rect 15436 -76588 15480 -76580
rect 15536 -76588 15580 -76580
rect 15636 -76588 15680 -76580
rect 15736 -76588 15780 -76580
rect 15836 -76588 15880 -76580
rect 15936 -76588 15980 -76580
rect 16036 -76588 16080 -76580
rect 16136 -76588 16180 -76580
rect 16236 -76588 16280 -76580
rect 16336 -76588 16380 -76580
rect 16436 -76588 16480 -76580
rect 16536 -76588 16580 -76580
rect 16636 -76588 16680 -76580
rect 16736 -76588 16780 -76580
rect 9280 -76632 9288 -76588
rect 9380 -76632 9388 -76588
rect 9480 -76632 9488 -76588
rect 9580 -76632 9588 -76588
rect 9680 -76632 9688 -76588
rect 9780 -76632 9788 -76588
rect 9880 -76632 9888 -76588
rect 9980 -76632 9988 -76588
rect 10080 -76632 10088 -76588
rect 10180 -76632 10188 -76588
rect 10280 -76632 10288 -76588
rect 10380 -76632 10388 -76588
rect 10480 -76632 10488 -76588
rect 10580 -76632 10588 -76588
rect 10680 -76632 10688 -76588
rect 10780 -76632 10788 -76588
rect 11280 -76632 11288 -76588
rect 11380 -76632 11388 -76588
rect 11480 -76632 11488 -76588
rect 11580 -76632 11588 -76588
rect 11680 -76632 11688 -76588
rect 11780 -76632 11788 -76588
rect 11880 -76632 11888 -76588
rect 11980 -76632 11988 -76588
rect 12080 -76632 12088 -76588
rect 12180 -76632 12188 -76588
rect 12280 -76632 12288 -76588
rect 12380 -76632 12388 -76588
rect 12480 -76632 12488 -76588
rect 12580 -76632 12588 -76588
rect 12680 -76632 12688 -76588
rect 12780 -76632 12788 -76588
rect 13280 -76632 13288 -76588
rect 13380 -76632 13388 -76588
rect 13480 -76632 13488 -76588
rect 13580 -76632 13588 -76588
rect 13680 -76632 13688 -76588
rect 13780 -76632 13788 -76588
rect 13880 -76632 13888 -76588
rect 13980 -76632 13988 -76588
rect 14080 -76632 14088 -76588
rect 14180 -76632 14188 -76588
rect 14280 -76632 14288 -76588
rect 14380 -76632 14388 -76588
rect 14480 -76632 14488 -76588
rect 14580 -76632 14588 -76588
rect 14680 -76632 14688 -76588
rect 14780 -76632 14788 -76588
rect 15280 -76632 15288 -76588
rect 15380 -76632 15388 -76588
rect 15480 -76632 15488 -76588
rect 15580 -76632 15588 -76588
rect 15680 -76632 15688 -76588
rect 15780 -76632 15788 -76588
rect 15880 -76632 15888 -76588
rect 15980 -76632 15988 -76588
rect 16080 -76632 16088 -76588
rect 16180 -76632 16188 -76588
rect 16280 -76632 16288 -76588
rect 16380 -76632 16388 -76588
rect 16480 -76632 16488 -76588
rect 16580 -76632 16588 -76588
rect 16680 -76632 16688 -76588
rect 16780 -76632 16788 -76588
rect 9236 -76688 9280 -76680
rect 9336 -76688 9380 -76680
rect 9436 -76688 9480 -76680
rect 9536 -76688 9580 -76680
rect 9636 -76688 9680 -76680
rect 9736 -76688 9780 -76680
rect 9836 -76688 9880 -76680
rect 9936 -76688 9980 -76680
rect 10036 -76688 10080 -76680
rect 10136 -76688 10180 -76680
rect 10236 -76688 10280 -76680
rect 10336 -76688 10380 -76680
rect 10436 -76688 10480 -76680
rect 10536 -76688 10580 -76680
rect 10636 -76688 10680 -76680
rect 10736 -76688 10780 -76680
rect 11236 -76688 11280 -76680
rect 11336 -76688 11380 -76680
rect 11436 -76688 11480 -76680
rect 11536 -76688 11580 -76680
rect 11636 -76688 11680 -76680
rect 11736 -76688 11780 -76680
rect 11836 -76688 11880 -76680
rect 11936 -76688 11980 -76680
rect 12036 -76688 12080 -76680
rect 12136 -76688 12180 -76680
rect 12236 -76688 12280 -76680
rect 12336 -76688 12380 -76680
rect 12436 -76688 12480 -76680
rect 12536 -76688 12580 -76680
rect 12636 -76688 12680 -76680
rect 12736 -76688 12780 -76680
rect 13236 -76688 13280 -76680
rect 13336 -76688 13380 -76680
rect 13436 -76688 13480 -76680
rect 13536 -76688 13580 -76680
rect 13636 -76688 13680 -76680
rect 13736 -76688 13780 -76680
rect 13836 -76688 13880 -76680
rect 13936 -76688 13980 -76680
rect 14036 -76688 14080 -76680
rect 14136 -76688 14180 -76680
rect 14236 -76688 14280 -76680
rect 14336 -76688 14380 -76680
rect 14436 -76688 14480 -76680
rect 14536 -76688 14580 -76680
rect 14636 -76688 14680 -76680
rect 14736 -76688 14780 -76680
rect 15236 -76688 15280 -76680
rect 15336 -76688 15380 -76680
rect 15436 -76688 15480 -76680
rect 15536 -76688 15580 -76680
rect 15636 -76688 15680 -76680
rect 15736 -76688 15780 -76680
rect 15836 -76688 15880 -76680
rect 15936 -76688 15980 -76680
rect 16036 -76688 16080 -76680
rect 16136 -76688 16180 -76680
rect 16236 -76688 16280 -76680
rect 16336 -76688 16380 -76680
rect 16436 -76688 16480 -76680
rect 16536 -76688 16580 -76680
rect 16636 -76688 16680 -76680
rect 16736 -76688 16780 -76680
rect 9280 -76732 9288 -76688
rect 9380 -76732 9388 -76688
rect 9480 -76732 9488 -76688
rect 9580 -76732 9588 -76688
rect 9680 -76732 9688 -76688
rect 9780 -76732 9788 -76688
rect 9880 -76732 9888 -76688
rect 9980 -76732 9988 -76688
rect 10080 -76732 10088 -76688
rect 10180 -76732 10188 -76688
rect 10280 -76732 10288 -76688
rect 10380 -76732 10388 -76688
rect 10480 -76732 10488 -76688
rect 10580 -76732 10588 -76688
rect 10680 -76732 10688 -76688
rect 10780 -76732 10788 -76688
rect 11280 -76732 11288 -76688
rect 11380 -76732 11388 -76688
rect 11480 -76732 11488 -76688
rect 11580 -76732 11588 -76688
rect 11680 -76732 11688 -76688
rect 11780 -76732 11788 -76688
rect 11880 -76732 11888 -76688
rect 11980 -76732 11988 -76688
rect 12080 -76732 12088 -76688
rect 12180 -76732 12188 -76688
rect 12280 -76732 12288 -76688
rect 12380 -76732 12388 -76688
rect 12480 -76732 12488 -76688
rect 12580 -76732 12588 -76688
rect 12680 -76732 12688 -76688
rect 12780 -76732 12788 -76688
rect 13280 -76732 13288 -76688
rect 13380 -76732 13388 -76688
rect 13480 -76732 13488 -76688
rect 13580 -76732 13588 -76688
rect 13680 -76732 13688 -76688
rect 13780 -76732 13788 -76688
rect 13880 -76732 13888 -76688
rect 13980 -76732 13988 -76688
rect 14080 -76732 14088 -76688
rect 14180 -76732 14188 -76688
rect 14280 -76732 14288 -76688
rect 14380 -76732 14388 -76688
rect 14480 -76732 14488 -76688
rect 14580 -76732 14588 -76688
rect 14680 -76732 14688 -76688
rect 14780 -76732 14788 -76688
rect 15280 -76732 15288 -76688
rect 15380 -76732 15388 -76688
rect 15480 -76732 15488 -76688
rect 15580 -76732 15588 -76688
rect 15680 -76732 15688 -76688
rect 15780 -76732 15788 -76688
rect 15880 -76732 15888 -76688
rect 15980 -76732 15988 -76688
rect 16080 -76732 16088 -76688
rect 16180 -76732 16188 -76688
rect 16280 -76732 16288 -76688
rect 16380 -76732 16388 -76688
rect 16480 -76732 16488 -76688
rect 16580 -76732 16588 -76688
rect 16680 -76732 16688 -76688
rect 16780 -76732 16788 -76688
rect -82968 -80459 -82924 -80451
rect -82868 -80459 -82824 -80451
rect -82768 -80459 -82724 -80451
rect -82668 -80459 -82624 -80451
rect -82568 -80459 -82524 -80451
rect -82468 -80459 -82424 -80451
rect -82368 -80459 -82324 -80451
rect -82268 -80459 -82224 -80451
rect -82168 -80459 -82124 -80451
rect -82068 -80459 -82024 -80451
rect -81968 -80459 -81924 -80451
rect -81868 -80459 -81824 -80451
rect -81768 -80459 -81724 -80451
rect -81668 -80459 -81624 -80451
rect -81568 -80459 -81524 -80451
rect -81468 -80459 -81424 -80451
rect -80968 -80459 -80924 -80451
rect -80868 -80459 -80824 -80451
rect -80768 -80459 -80724 -80451
rect -80668 -80459 -80624 -80451
rect -80568 -80459 -80524 -80451
rect -80468 -80459 -80424 -80451
rect -80368 -80459 -80324 -80451
rect -80268 -80459 -80224 -80451
rect -80168 -80459 -80124 -80451
rect -80068 -80459 -80024 -80451
rect -79968 -80459 -79924 -80451
rect -79868 -80459 -79824 -80451
rect -79768 -80459 -79724 -80451
rect -79668 -80459 -79624 -80451
rect -79568 -80459 -79524 -80451
rect -79468 -80459 -79424 -80451
rect -78968 -80459 -78924 -80451
rect -78868 -80459 -78824 -80451
rect -78768 -80459 -78724 -80451
rect -78668 -80459 -78624 -80451
rect -78568 -80459 -78524 -80451
rect -78468 -80459 -78424 -80451
rect -78368 -80459 -78324 -80451
rect -78268 -80459 -78224 -80451
rect -78168 -80459 -78124 -80451
rect -78068 -80459 -78024 -80451
rect -77968 -80459 -77924 -80451
rect -77868 -80459 -77824 -80451
rect -77768 -80459 -77724 -80451
rect -77668 -80459 -77624 -80451
rect -77568 -80459 -77524 -80451
rect -77468 -80459 -77424 -80451
rect -76968 -80459 -76924 -80451
rect -76868 -80459 -76824 -80451
rect -76768 -80459 -76724 -80451
rect -76668 -80459 -76624 -80451
rect -76568 -80459 -76524 -80451
rect -76468 -80459 -76424 -80451
rect -76368 -80459 -76324 -80451
rect -76268 -80459 -76224 -80451
rect -76168 -80459 -76124 -80451
rect -76068 -80459 -76024 -80451
rect -75968 -80459 -75924 -80451
rect -75868 -80459 -75824 -80451
rect -75768 -80459 -75724 -80451
rect -75668 -80459 -75624 -80451
rect -75568 -80459 -75524 -80451
rect -75468 -80459 -75424 -80451
rect -82924 -80503 -82916 -80459
rect -82824 -80503 -82816 -80459
rect -82724 -80503 -82716 -80459
rect -82624 -80503 -82616 -80459
rect -82524 -80503 -82516 -80459
rect -82424 -80503 -82416 -80459
rect -82324 -80503 -82316 -80459
rect -82224 -80503 -82216 -80459
rect -82124 -80503 -82116 -80459
rect -82024 -80503 -82016 -80459
rect -81924 -80503 -81916 -80459
rect -81824 -80503 -81816 -80459
rect -81724 -80503 -81716 -80459
rect -81624 -80503 -81616 -80459
rect -81524 -80503 -81516 -80459
rect -81424 -80503 -81416 -80459
rect -80924 -80503 -80916 -80459
rect -80824 -80503 -80816 -80459
rect -80724 -80503 -80716 -80459
rect -80624 -80503 -80616 -80459
rect -80524 -80503 -80516 -80459
rect -80424 -80503 -80416 -80459
rect -80324 -80503 -80316 -80459
rect -80224 -80503 -80216 -80459
rect -80124 -80503 -80116 -80459
rect -80024 -80503 -80016 -80459
rect -79924 -80503 -79916 -80459
rect -79824 -80503 -79816 -80459
rect -79724 -80503 -79716 -80459
rect -79624 -80503 -79616 -80459
rect -79524 -80503 -79516 -80459
rect -79424 -80503 -79416 -80459
rect -78924 -80503 -78916 -80459
rect -78824 -80503 -78816 -80459
rect -78724 -80503 -78716 -80459
rect -78624 -80503 -78616 -80459
rect -78524 -80503 -78516 -80459
rect -78424 -80503 -78416 -80459
rect -78324 -80503 -78316 -80459
rect -78224 -80503 -78216 -80459
rect -78124 -80503 -78116 -80459
rect -78024 -80503 -78016 -80459
rect -77924 -80503 -77916 -80459
rect -77824 -80503 -77816 -80459
rect -77724 -80503 -77716 -80459
rect -77624 -80503 -77616 -80459
rect -77524 -80503 -77516 -80459
rect -77424 -80503 -77416 -80459
rect -76924 -80503 -76916 -80459
rect -76824 -80503 -76816 -80459
rect -76724 -80503 -76716 -80459
rect -76624 -80503 -76616 -80459
rect -76524 -80503 -76516 -80459
rect -76424 -80503 -76416 -80459
rect -76324 -80503 -76316 -80459
rect -76224 -80503 -76216 -80459
rect -76124 -80503 -76116 -80459
rect -76024 -80503 -76016 -80459
rect -75924 -80503 -75916 -80459
rect -75824 -80503 -75816 -80459
rect -75724 -80503 -75716 -80459
rect -75624 -80503 -75616 -80459
rect -75524 -80503 -75516 -80459
rect -75424 -80503 -75416 -80459
rect -50017 -80461 -49973 -80453
rect -49917 -80461 -49873 -80453
rect -49817 -80461 -49773 -80453
rect -49717 -80461 -49673 -80453
rect -49617 -80461 -49573 -80453
rect -49517 -80461 -49473 -80453
rect -49417 -80461 -49373 -80453
rect -49317 -80461 -49273 -80453
rect -49217 -80461 -49173 -80453
rect -49117 -80461 -49073 -80453
rect -49017 -80461 -48973 -80453
rect -48917 -80461 -48873 -80453
rect -48817 -80461 -48773 -80453
rect -48717 -80461 -48673 -80453
rect -48617 -80461 -48573 -80453
rect -48517 -80461 -48473 -80453
rect -48017 -80461 -47973 -80453
rect -47917 -80461 -47873 -80453
rect -47817 -80461 -47773 -80453
rect -47717 -80461 -47673 -80453
rect -47617 -80461 -47573 -80453
rect -47517 -80461 -47473 -80453
rect -47417 -80461 -47373 -80453
rect -47317 -80461 -47273 -80453
rect -47217 -80461 -47173 -80453
rect -47117 -80461 -47073 -80453
rect -47017 -80461 -46973 -80453
rect -46917 -80461 -46873 -80453
rect -46817 -80461 -46773 -80453
rect -46717 -80461 -46673 -80453
rect -46617 -80461 -46573 -80453
rect -46517 -80461 -46473 -80453
rect -46017 -80461 -45973 -80453
rect -45917 -80461 -45873 -80453
rect -45817 -80461 -45773 -80453
rect -45717 -80461 -45673 -80453
rect -45617 -80461 -45573 -80453
rect -45517 -80461 -45473 -80453
rect -45417 -80461 -45373 -80453
rect -45317 -80461 -45273 -80453
rect -45217 -80461 -45173 -80453
rect -45117 -80461 -45073 -80453
rect -45017 -80461 -44973 -80453
rect -44917 -80461 -44873 -80453
rect -44817 -80461 -44773 -80453
rect -44717 -80461 -44673 -80453
rect -44617 -80461 -44573 -80453
rect -44517 -80461 -44473 -80453
rect -44017 -80461 -43973 -80453
rect -43917 -80461 -43873 -80453
rect -43817 -80461 -43773 -80453
rect -43717 -80461 -43673 -80453
rect -43617 -80461 -43573 -80453
rect -43517 -80461 -43473 -80453
rect -43417 -80461 -43373 -80453
rect -43317 -80461 -43273 -80453
rect -43217 -80461 -43173 -80453
rect -43117 -80461 -43073 -80453
rect -43017 -80461 -42973 -80453
rect -42917 -80461 -42873 -80453
rect -42817 -80461 -42773 -80453
rect -42717 -80461 -42673 -80453
rect -42617 -80461 -42573 -80453
rect -42517 -80461 -42473 -80453
rect 80737 -80455 80781 -80447
rect 80837 -80455 80881 -80447
rect 80937 -80455 80981 -80447
rect 81037 -80455 81081 -80447
rect 81137 -80455 81181 -80447
rect 81237 -80455 81281 -80447
rect 81337 -80455 81381 -80447
rect 81437 -80455 81481 -80447
rect 81537 -80455 81581 -80447
rect 81637 -80455 81681 -80447
rect 81737 -80455 81781 -80447
rect 81837 -80455 81881 -80447
rect 81937 -80455 81981 -80447
rect 82037 -80455 82081 -80447
rect 82137 -80455 82181 -80447
rect 82237 -80455 82281 -80447
rect 82737 -80455 82781 -80447
rect 82837 -80455 82881 -80447
rect 82937 -80455 82981 -80447
rect 83037 -80455 83081 -80447
rect 83137 -80455 83181 -80447
rect 83237 -80455 83281 -80447
rect 83337 -80455 83381 -80447
rect 83437 -80455 83481 -80447
rect 83537 -80455 83581 -80447
rect 83637 -80455 83681 -80447
rect 83737 -80455 83781 -80447
rect 83837 -80455 83881 -80447
rect 83937 -80455 83981 -80447
rect 84037 -80455 84081 -80447
rect 84137 -80455 84181 -80447
rect 84237 -80455 84281 -80447
rect 84737 -80455 84781 -80447
rect 84837 -80455 84881 -80447
rect 84937 -80455 84981 -80447
rect 85037 -80455 85081 -80447
rect 85137 -80455 85181 -80447
rect 85237 -80455 85281 -80447
rect 85337 -80455 85381 -80447
rect 85437 -80455 85481 -80447
rect 85537 -80455 85581 -80447
rect 85637 -80455 85681 -80447
rect 85737 -80455 85781 -80447
rect 85837 -80455 85881 -80447
rect 85937 -80455 85981 -80447
rect 86037 -80455 86081 -80447
rect 86137 -80455 86181 -80447
rect 86237 -80455 86281 -80447
rect 86737 -80455 86781 -80447
rect 86837 -80455 86881 -80447
rect 86937 -80455 86981 -80447
rect 87037 -80455 87081 -80447
rect 87137 -80455 87181 -80447
rect 87237 -80455 87281 -80447
rect 87337 -80455 87381 -80447
rect 87437 -80455 87481 -80447
rect 87537 -80455 87581 -80447
rect 87637 -80455 87681 -80447
rect 87737 -80455 87781 -80447
rect 87837 -80455 87881 -80447
rect 87937 -80455 87981 -80447
rect 88037 -80455 88081 -80447
rect 88137 -80455 88181 -80447
rect 88237 -80455 88281 -80447
rect -49973 -80505 -49965 -80461
rect -49873 -80505 -49865 -80461
rect -49773 -80505 -49765 -80461
rect -49673 -80505 -49665 -80461
rect -49573 -80505 -49565 -80461
rect -49473 -80505 -49465 -80461
rect -49373 -80505 -49365 -80461
rect -49273 -80505 -49265 -80461
rect -49173 -80505 -49165 -80461
rect -49073 -80505 -49065 -80461
rect -48973 -80505 -48965 -80461
rect -48873 -80505 -48865 -80461
rect -48773 -80505 -48765 -80461
rect -48673 -80505 -48665 -80461
rect -48573 -80505 -48565 -80461
rect -48473 -80505 -48465 -80461
rect -47973 -80505 -47965 -80461
rect -47873 -80505 -47865 -80461
rect -47773 -80505 -47765 -80461
rect -47673 -80505 -47665 -80461
rect -47573 -80505 -47565 -80461
rect -47473 -80505 -47465 -80461
rect -47373 -80505 -47365 -80461
rect -47273 -80505 -47265 -80461
rect -47173 -80505 -47165 -80461
rect -47073 -80505 -47065 -80461
rect -46973 -80505 -46965 -80461
rect -46873 -80505 -46865 -80461
rect -46773 -80505 -46765 -80461
rect -46673 -80505 -46665 -80461
rect -46573 -80505 -46565 -80461
rect -46473 -80505 -46465 -80461
rect -45973 -80505 -45965 -80461
rect -45873 -80505 -45865 -80461
rect -45773 -80505 -45765 -80461
rect -45673 -80505 -45665 -80461
rect -45573 -80505 -45565 -80461
rect -45473 -80505 -45465 -80461
rect -45373 -80505 -45365 -80461
rect -45273 -80505 -45265 -80461
rect -45173 -80505 -45165 -80461
rect -45073 -80505 -45065 -80461
rect -44973 -80505 -44965 -80461
rect -44873 -80505 -44865 -80461
rect -44773 -80505 -44765 -80461
rect -44673 -80505 -44665 -80461
rect -44573 -80505 -44565 -80461
rect -44473 -80505 -44465 -80461
rect -43973 -80505 -43965 -80461
rect -43873 -80505 -43865 -80461
rect -43773 -80505 -43765 -80461
rect -43673 -80505 -43665 -80461
rect -43573 -80505 -43565 -80461
rect -43473 -80505 -43465 -80461
rect -43373 -80505 -43365 -80461
rect -43273 -80505 -43265 -80461
rect -43173 -80505 -43165 -80461
rect -43073 -80505 -43065 -80461
rect -42973 -80505 -42965 -80461
rect -42873 -80505 -42865 -80461
rect -42773 -80505 -42765 -80461
rect -42673 -80505 -42665 -80461
rect -42573 -80505 -42565 -80461
rect -42473 -80505 -42465 -80461
rect 80781 -80499 80789 -80455
rect 80881 -80499 80889 -80455
rect 80981 -80499 80989 -80455
rect 81081 -80499 81089 -80455
rect 81181 -80499 81189 -80455
rect 81281 -80499 81289 -80455
rect 81381 -80499 81389 -80455
rect 81481 -80499 81489 -80455
rect 81581 -80499 81589 -80455
rect 81681 -80499 81689 -80455
rect 81781 -80499 81789 -80455
rect 81881 -80499 81889 -80455
rect 81981 -80499 81989 -80455
rect 82081 -80499 82089 -80455
rect 82181 -80499 82189 -80455
rect 82281 -80499 82289 -80455
rect 82781 -80499 82789 -80455
rect 82881 -80499 82889 -80455
rect 82981 -80499 82989 -80455
rect 83081 -80499 83089 -80455
rect 83181 -80499 83189 -80455
rect 83281 -80499 83289 -80455
rect 83381 -80499 83389 -80455
rect 83481 -80499 83489 -80455
rect 83581 -80499 83589 -80455
rect 83681 -80499 83689 -80455
rect 83781 -80499 83789 -80455
rect 83881 -80499 83889 -80455
rect 83981 -80499 83989 -80455
rect 84081 -80499 84089 -80455
rect 84181 -80499 84189 -80455
rect 84281 -80499 84289 -80455
rect 84781 -80499 84789 -80455
rect 84881 -80499 84889 -80455
rect 84981 -80499 84989 -80455
rect 85081 -80499 85089 -80455
rect 85181 -80499 85189 -80455
rect 85281 -80499 85289 -80455
rect 85381 -80499 85389 -80455
rect 85481 -80499 85489 -80455
rect 85581 -80499 85589 -80455
rect 85681 -80499 85689 -80455
rect 85781 -80499 85789 -80455
rect 85881 -80499 85889 -80455
rect 85981 -80499 85989 -80455
rect 86081 -80499 86089 -80455
rect 86181 -80499 86189 -80455
rect 86281 -80499 86289 -80455
rect 86781 -80499 86789 -80455
rect 86881 -80499 86889 -80455
rect 86981 -80499 86989 -80455
rect 87081 -80499 87089 -80455
rect 87181 -80499 87189 -80455
rect 87281 -80499 87289 -80455
rect 87381 -80499 87389 -80455
rect 87481 -80499 87489 -80455
rect 87581 -80499 87589 -80455
rect 87681 -80499 87689 -80455
rect 87781 -80499 87789 -80455
rect 87881 -80499 87889 -80455
rect 87981 -80499 87989 -80455
rect 88081 -80499 88089 -80455
rect 88181 -80499 88189 -80455
rect 88281 -80499 88289 -80455
rect -82968 -80559 -82924 -80551
rect -82868 -80559 -82824 -80551
rect -82768 -80559 -82724 -80551
rect -82668 -80559 -82624 -80551
rect -82568 -80559 -82524 -80551
rect -82468 -80559 -82424 -80551
rect -82368 -80559 -82324 -80551
rect -82268 -80559 -82224 -80551
rect -82168 -80559 -82124 -80551
rect -82068 -80559 -82024 -80551
rect -81968 -80559 -81924 -80551
rect -81868 -80559 -81824 -80551
rect -81768 -80559 -81724 -80551
rect -81668 -80559 -81624 -80551
rect -81568 -80559 -81524 -80551
rect -81468 -80559 -81424 -80551
rect -80968 -80559 -80924 -80551
rect -80868 -80559 -80824 -80551
rect -80768 -80559 -80724 -80551
rect -80668 -80559 -80624 -80551
rect -80568 -80559 -80524 -80551
rect -80468 -80559 -80424 -80551
rect -80368 -80559 -80324 -80551
rect -80268 -80559 -80224 -80551
rect -80168 -80559 -80124 -80551
rect -80068 -80559 -80024 -80551
rect -79968 -80559 -79924 -80551
rect -79868 -80559 -79824 -80551
rect -79768 -80559 -79724 -80551
rect -79668 -80559 -79624 -80551
rect -79568 -80559 -79524 -80551
rect -79468 -80559 -79424 -80551
rect -78968 -80559 -78924 -80551
rect -78868 -80559 -78824 -80551
rect -78768 -80559 -78724 -80551
rect -78668 -80559 -78624 -80551
rect -78568 -80559 -78524 -80551
rect -78468 -80559 -78424 -80551
rect -78368 -80559 -78324 -80551
rect -78268 -80559 -78224 -80551
rect -78168 -80559 -78124 -80551
rect -78068 -80559 -78024 -80551
rect -77968 -80559 -77924 -80551
rect -77868 -80559 -77824 -80551
rect -77768 -80559 -77724 -80551
rect -77668 -80559 -77624 -80551
rect -77568 -80559 -77524 -80551
rect -77468 -80559 -77424 -80551
rect -76968 -80559 -76924 -80551
rect -76868 -80559 -76824 -80551
rect -76768 -80559 -76724 -80551
rect -76668 -80559 -76624 -80551
rect -76568 -80559 -76524 -80551
rect -76468 -80559 -76424 -80551
rect -76368 -80559 -76324 -80551
rect -76268 -80559 -76224 -80551
rect -76168 -80559 -76124 -80551
rect -76068 -80559 -76024 -80551
rect -75968 -80559 -75924 -80551
rect -75868 -80559 -75824 -80551
rect -75768 -80559 -75724 -80551
rect -75668 -80559 -75624 -80551
rect -75568 -80559 -75524 -80551
rect -75468 -80559 -75424 -80551
rect -82924 -80603 -82916 -80559
rect -82824 -80603 -82816 -80559
rect -82724 -80603 -82716 -80559
rect -82624 -80603 -82616 -80559
rect -82524 -80603 -82516 -80559
rect -82424 -80603 -82416 -80559
rect -82324 -80603 -82316 -80559
rect -82224 -80603 -82216 -80559
rect -82124 -80603 -82116 -80559
rect -82024 -80603 -82016 -80559
rect -81924 -80603 -81916 -80559
rect -81824 -80603 -81816 -80559
rect -81724 -80603 -81716 -80559
rect -81624 -80603 -81616 -80559
rect -81524 -80603 -81516 -80559
rect -81424 -80603 -81416 -80559
rect -80924 -80603 -80916 -80559
rect -80824 -80603 -80816 -80559
rect -80724 -80603 -80716 -80559
rect -80624 -80603 -80616 -80559
rect -80524 -80603 -80516 -80559
rect -80424 -80603 -80416 -80559
rect -80324 -80603 -80316 -80559
rect -80224 -80603 -80216 -80559
rect -80124 -80603 -80116 -80559
rect -80024 -80603 -80016 -80559
rect -79924 -80603 -79916 -80559
rect -79824 -80603 -79816 -80559
rect -79724 -80603 -79716 -80559
rect -79624 -80603 -79616 -80559
rect -79524 -80603 -79516 -80559
rect -79424 -80603 -79416 -80559
rect -78924 -80603 -78916 -80559
rect -78824 -80603 -78816 -80559
rect -78724 -80603 -78716 -80559
rect -78624 -80603 -78616 -80559
rect -78524 -80603 -78516 -80559
rect -78424 -80603 -78416 -80559
rect -78324 -80603 -78316 -80559
rect -78224 -80603 -78216 -80559
rect -78124 -80603 -78116 -80559
rect -78024 -80603 -78016 -80559
rect -77924 -80603 -77916 -80559
rect -77824 -80603 -77816 -80559
rect -77724 -80603 -77716 -80559
rect -77624 -80603 -77616 -80559
rect -77524 -80603 -77516 -80559
rect -77424 -80603 -77416 -80559
rect -76924 -80603 -76916 -80559
rect -76824 -80603 -76816 -80559
rect -76724 -80603 -76716 -80559
rect -76624 -80603 -76616 -80559
rect -76524 -80603 -76516 -80559
rect -76424 -80603 -76416 -80559
rect -76324 -80603 -76316 -80559
rect -76224 -80603 -76216 -80559
rect -76124 -80603 -76116 -80559
rect -76024 -80603 -76016 -80559
rect -75924 -80603 -75916 -80559
rect -75824 -80603 -75816 -80559
rect -75724 -80603 -75716 -80559
rect -75624 -80603 -75616 -80559
rect -75524 -80603 -75516 -80559
rect -75424 -80603 -75416 -80559
rect -50017 -80561 -49973 -80553
rect -49917 -80561 -49873 -80553
rect -49817 -80561 -49773 -80553
rect -49717 -80561 -49673 -80553
rect -49617 -80561 -49573 -80553
rect -49517 -80561 -49473 -80553
rect -49417 -80561 -49373 -80553
rect -49317 -80561 -49273 -80553
rect -49217 -80561 -49173 -80553
rect -49117 -80561 -49073 -80553
rect -49017 -80561 -48973 -80553
rect -48917 -80561 -48873 -80553
rect -48817 -80561 -48773 -80553
rect -48717 -80561 -48673 -80553
rect -48617 -80561 -48573 -80553
rect -48517 -80561 -48473 -80553
rect -48017 -80561 -47973 -80553
rect -47917 -80561 -47873 -80553
rect -47817 -80561 -47773 -80553
rect -47717 -80561 -47673 -80553
rect -47617 -80561 -47573 -80553
rect -47517 -80561 -47473 -80553
rect -47417 -80561 -47373 -80553
rect -47317 -80561 -47273 -80553
rect -47217 -80561 -47173 -80553
rect -47117 -80561 -47073 -80553
rect -47017 -80561 -46973 -80553
rect -46917 -80561 -46873 -80553
rect -46817 -80561 -46773 -80553
rect -46717 -80561 -46673 -80553
rect -46617 -80561 -46573 -80553
rect -46517 -80561 -46473 -80553
rect -46017 -80561 -45973 -80553
rect -45917 -80561 -45873 -80553
rect -45817 -80561 -45773 -80553
rect -45717 -80561 -45673 -80553
rect -45617 -80561 -45573 -80553
rect -45517 -80561 -45473 -80553
rect -45417 -80561 -45373 -80553
rect -45317 -80561 -45273 -80553
rect -45217 -80561 -45173 -80553
rect -45117 -80561 -45073 -80553
rect -45017 -80561 -44973 -80553
rect -44917 -80561 -44873 -80553
rect -44817 -80561 -44773 -80553
rect -44717 -80561 -44673 -80553
rect -44617 -80561 -44573 -80553
rect -44517 -80561 -44473 -80553
rect -44017 -80561 -43973 -80553
rect -43917 -80561 -43873 -80553
rect -43817 -80561 -43773 -80553
rect -43717 -80561 -43673 -80553
rect -43617 -80561 -43573 -80553
rect -43517 -80561 -43473 -80553
rect -43417 -80561 -43373 -80553
rect -43317 -80561 -43273 -80553
rect -43217 -80561 -43173 -80553
rect -43117 -80561 -43073 -80553
rect -43017 -80561 -42973 -80553
rect -42917 -80561 -42873 -80553
rect -42817 -80561 -42773 -80553
rect -42717 -80561 -42673 -80553
rect -42617 -80561 -42573 -80553
rect -42517 -80561 -42473 -80553
rect 80737 -80555 80781 -80547
rect 80837 -80555 80881 -80547
rect 80937 -80555 80981 -80547
rect 81037 -80555 81081 -80547
rect 81137 -80555 81181 -80547
rect 81237 -80555 81281 -80547
rect 81337 -80555 81381 -80547
rect 81437 -80555 81481 -80547
rect 81537 -80555 81581 -80547
rect 81637 -80555 81681 -80547
rect 81737 -80555 81781 -80547
rect 81837 -80555 81881 -80547
rect 81937 -80555 81981 -80547
rect 82037 -80555 82081 -80547
rect 82137 -80555 82181 -80547
rect 82237 -80555 82281 -80547
rect 82737 -80555 82781 -80547
rect 82837 -80555 82881 -80547
rect 82937 -80555 82981 -80547
rect 83037 -80555 83081 -80547
rect 83137 -80555 83181 -80547
rect 83237 -80555 83281 -80547
rect 83337 -80555 83381 -80547
rect 83437 -80555 83481 -80547
rect 83537 -80555 83581 -80547
rect 83637 -80555 83681 -80547
rect 83737 -80555 83781 -80547
rect 83837 -80555 83881 -80547
rect 83937 -80555 83981 -80547
rect 84037 -80555 84081 -80547
rect 84137 -80555 84181 -80547
rect 84237 -80555 84281 -80547
rect 84737 -80555 84781 -80547
rect 84837 -80555 84881 -80547
rect 84937 -80555 84981 -80547
rect 85037 -80555 85081 -80547
rect 85137 -80555 85181 -80547
rect 85237 -80555 85281 -80547
rect 85337 -80555 85381 -80547
rect 85437 -80555 85481 -80547
rect 85537 -80555 85581 -80547
rect 85637 -80555 85681 -80547
rect 85737 -80555 85781 -80547
rect 85837 -80555 85881 -80547
rect 85937 -80555 85981 -80547
rect 86037 -80555 86081 -80547
rect 86137 -80555 86181 -80547
rect 86237 -80555 86281 -80547
rect 86737 -80555 86781 -80547
rect 86837 -80555 86881 -80547
rect 86937 -80555 86981 -80547
rect 87037 -80555 87081 -80547
rect 87137 -80555 87181 -80547
rect 87237 -80555 87281 -80547
rect 87337 -80555 87381 -80547
rect 87437 -80555 87481 -80547
rect 87537 -80555 87581 -80547
rect 87637 -80555 87681 -80547
rect 87737 -80555 87781 -80547
rect 87837 -80555 87881 -80547
rect 87937 -80555 87981 -80547
rect 88037 -80555 88081 -80547
rect 88137 -80555 88181 -80547
rect 88237 -80555 88281 -80547
rect -49973 -80605 -49965 -80561
rect -49873 -80605 -49865 -80561
rect -49773 -80605 -49765 -80561
rect -49673 -80605 -49665 -80561
rect -49573 -80605 -49565 -80561
rect -49473 -80605 -49465 -80561
rect -49373 -80605 -49365 -80561
rect -49273 -80605 -49265 -80561
rect -49173 -80605 -49165 -80561
rect -49073 -80605 -49065 -80561
rect -48973 -80605 -48965 -80561
rect -48873 -80605 -48865 -80561
rect -48773 -80605 -48765 -80561
rect -48673 -80605 -48665 -80561
rect -48573 -80605 -48565 -80561
rect -48473 -80605 -48465 -80561
rect -47973 -80605 -47965 -80561
rect -47873 -80605 -47865 -80561
rect -47773 -80605 -47765 -80561
rect -47673 -80605 -47665 -80561
rect -47573 -80605 -47565 -80561
rect -47473 -80605 -47465 -80561
rect -47373 -80605 -47365 -80561
rect -47273 -80605 -47265 -80561
rect -47173 -80605 -47165 -80561
rect -47073 -80605 -47065 -80561
rect -46973 -80605 -46965 -80561
rect -46873 -80605 -46865 -80561
rect -46773 -80605 -46765 -80561
rect -46673 -80605 -46665 -80561
rect -46573 -80605 -46565 -80561
rect -46473 -80605 -46465 -80561
rect -45973 -80605 -45965 -80561
rect -45873 -80605 -45865 -80561
rect -45773 -80605 -45765 -80561
rect -45673 -80605 -45665 -80561
rect -45573 -80605 -45565 -80561
rect -45473 -80605 -45465 -80561
rect -45373 -80605 -45365 -80561
rect -45273 -80605 -45265 -80561
rect -45173 -80605 -45165 -80561
rect -45073 -80605 -45065 -80561
rect -44973 -80605 -44965 -80561
rect -44873 -80605 -44865 -80561
rect -44773 -80605 -44765 -80561
rect -44673 -80605 -44665 -80561
rect -44573 -80605 -44565 -80561
rect -44473 -80605 -44465 -80561
rect -43973 -80605 -43965 -80561
rect -43873 -80605 -43865 -80561
rect -43773 -80605 -43765 -80561
rect -43673 -80605 -43665 -80561
rect -43573 -80605 -43565 -80561
rect -43473 -80605 -43465 -80561
rect -43373 -80605 -43365 -80561
rect -43273 -80605 -43265 -80561
rect -43173 -80605 -43165 -80561
rect -43073 -80605 -43065 -80561
rect -42973 -80605 -42965 -80561
rect -42873 -80605 -42865 -80561
rect -42773 -80605 -42765 -80561
rect -42673 -80605 -42665 -80561
rect -42573 -80605 -42565 -80561
rect -42473 -80605 -42465 -80561
rect 80781 -80599 80789 -80555
rect 80881 -80599 80889 -80555
rect 80981 -80599 80989 -80555
rect 81081 -80599 81089 -80555
rect 81181 -80599 81189 -80555
rect 81281 -80599 81289 -80555
rect 81381 -80599 81389 -80555
rect 81481 -80599 81489 -80555
rect 81581 -80599 81589 -80555
rect 81681 -80599 81689 -80555
rect 81781 -80599 81789 -80555
rect 81881 -80599 81889 -80555
rect 81981 -80599 81989 -80555
rect 82081 -80599 82089 -80555
rect 82181 -80599 82189 -80555
rect 82281 -80599 82289 -80555
rect 82781 -80599 82789 -80555
rect 82881 -80599 82889 -80555
rect 82981 -80599 82989 -80555
rect 83081 -80599 83089 -80555
rect 83181 -80599 83189 -80555
rect 83281 -80599 83289 -80555
rect 83381 -80599 83389 -80555
rect 83481 -80599 83489 -80555
rect 83581 -80599 83589 -80555
rect 83681 -80599 83689 -80555
rect 83781 -80599 83789 -80555
rect 83881 -80599 83889 -80555
rect 83981 -80599 83989 -80555
rect 84081 -80599 84089 -80555
rect 84181 -80599 84189 -80555
rect 84281 -80599 84289 -80555
rect 84781 -80599 84789 -80555
rect 84881 -80599 84889 -80555
rect 84981 -80599 84989 -80555
rect 85081 -80599 85089 -80555
rect 85181 -80599 85189 -80555
rect 85281 -80599 85289 -80555
rect 85381 -80599 85389 -80555
rect 85481 -80599 85489 -80555
rect 85581 -80599 85589 -80555
rect 85681 -80599 85689 -80555
rect 85781 -80599 85789 -80555
rect 85881 -80599 85889 -80555
rect 85981 -80599 85989 -80555
rect 86081 -80599 86089 -80555
rect 86181 -80599 86189 -80555
rect 86281 -80599 86289 -80555
rect 86781 -80599 86789 -80555
rect 86881 -80599 86889 -80555
rect 86981 -80599 86989 -80555
rect 87081 -80599 87089 -80555
rect 87181 -80599 87189 -80555
rect 87281 -80599 87289 -80555
rect 87381 -80599 87389 -80555
rect 87481 -80599 87489 -80555
rect 87581 -80599 87589 -80555
rect 87681 -80599 87689 -80555
rect 87781 -80599 87789 -80555
rect 87881 -80599 87889 -80555
rect 87981 -80599 87989 -80555
rect 88081 -80599 88089 -80555
rect 88181 -80599 88189 -80555
rect 88281 -80599 88289 -80555
rect -82968 -80659 -82924 -80651
rect -82868 -80659 -82824 -80651
rect -82768 -80659 -82724 -80651
rect -82668 -80659 -82624 -80651
rect -82568 -80659 -82524 -80651
rect -82468 -80659 -82424 -80651
rect -82368 -80659 -82324 -80651
rect -82268 -80659 -82224 -80651
rect -82168 -80659 -82124 -80651
rect -82068 -80659 -82024 -80651
rect -81968 -80659 -81924 -80651
rect -81868 -80659 -81824 -80651
rect -81768 -80659 -81724 -80651
rect -81668 -80659 -81624 -80651
rect -81568 -80659 -81524 -80651
rect -81468 -80659 -81424 -80651
rect -80968 -80659 -80924 -80651
rect -80868 -80659 -80824 -80651
rect -80768 -80659 -80724 -80651
rect -80668 -80659 -80624 -80651
rect -80568 -80659 -80524 -80651
rect -80468 -80659 -80424 -80651
rect -80368 -80659 -80324 -80651
rect -80268 -80659 -80224 -80651
rect -80168 -80659 -80124 -80651
rect -80068 -80659 -80024 -80651
rect -79968 -80659 -79924 -80651
rect -79868 -80659 -79824 -80651
rect -79768 -80659 -79724 -80651
rect -79668 -80659 -79624 -80651
rect -79568 -80659 -79524 -80651
rect -79468 -80659 -79424 -80651
rect -78968 -80659 -78924 -80651
rect -78868 -80659 -78824 -80651
rect -78768 -80659 -78724 -80651
rect -78668 -80659 -78624 -80651
rect -78568 -80659 -78524 -80651
rect -78468 -80659 -78424 -80651
rect -78368 -80659 -78324 -80651
rect -78268 -80659 -78224 -80651
rect -78168 -80659 -78124 -80651
rect -78068 -80659 -78024 -80651
rect -77968 -80659 -77924 -80651
rect -77868 -80659 -77824 -80651
rect -77768 -80659 -77724 -80651
rect -77668 -80659 -77624 -80651
rect -77568 -80659 -77524 -80651
rect -77468 -80659 -77424 -80651
rect -76968 -80659 -76924 -80651
rect -76868 -80659 -76824 -80651
rect -76768 -80659 -76724 -80651
rect -76668 -80659 -76624 -80651
rect -76568 -80659 -76524 -80651
rect -76468 -80659 -76424 -80651
rect -76368 -80659 -76324 -80651
rect -76268 -80659 -76224 -80651
rect -76168 -80659 -76124 -80651
rect -76068 -80659 -76024 -80651
rect -75968 -80659 -75924 -80651
rect -75868 -80659 -75824 -80651
rect -75768 -80659 -75724 -80651
rect -75668 -80659 -75624 -80651
rect -75568 -80659 -75524 -80651
rect -75468 -80659 -75424 -80651
rect -82924 -80703 -82916 -80659
rect -82824 -80703 -82816 -80659
rect -82724 -80703 -82716 -80659
rect -82624 -80703 -82616 -80659
rect -82524 -80703 -82516 -80659
rect -82424 -80703 -82416 -80659
rect -82324 -80703 -82316 -80659
rect -82224 -80703 -82216 -80659
rect -82124 -80703 -82116 -80659
rect -82024 -80703 -82016 -80659
rect -81924 -80703 -81916 -80659
rect -81824 -80703 -81816 -80659
rect -81724 -80703 -81716 -80659
rect -81624 -80703 -81616 -80659
rect -81524 -80703 -81516 -80659
rect -81424 -80703 -81416 -80659
rect -80924 -80703 -80916 -80659
rect -80824 -80703 -80816 -80659
rect -80724 -80703 -80716 -80659
rect -80624 -80703 -80616 -80659
rect -80524 -80703 -80516 -80659
rect -80424 -80703 -80416 -80659
rect -80324 -80703 -80316 -80659
rect -80224 -80703 -80216 -80659
rect -80124 -80703 -80116 -80659
rect -80024 -80703 -80016 -80659
rect -79924 -80703 -79916 -80659
rect -79824 -80703 -79816 -80659
rect -79724 -80703 -79716 -80659
rect -79624 -80703 -79616 -80659
rect -79524 -80703 -79516 -80659
rect -79424 -80703 -79416 -80659
rect -78924 -80703 -78916 -80659
rect -78824 -80703 -78816 -80659
rect -78724 -80703 -78716 -80659
rect -78624 -80703 -78616 -80659
rect -78524 -80703 -78516 -80659
rect -78424 -80703 -78416 -80659
rect -78324 -80703 -78316 -80659
rect -78224 -80703 -78216 -80659
rect -78124 -80703 -78116 -80659
rect -78024 -80703 -78016 -80659
rect -77924 -80703 -77916 -80659
rect -77824 -80703 -77816 -80659
rect -77724 -80703 -77716 -80659
rect -77624 -80703 -77616 -80659
rect -77524 -80703 -77516 -80659
rect -77424 -80703 -77416 -80659
rect -76924 -80703 -76916 -80659
rect -76824 -80703 -76816 -80659
rect -76724 -80703 -76716 -80659
rect -76624 -80703 -76616 -80659
rect -76524 -80703 -76516 -80659
rect -76424 -80703 -76416 -80659
rect -76324 -80703 -76316 -80659
rect -76224 -80703 -76216 -80659
rect -76124 -80703 -76116 -80659
rect -76024 -80703 -76016 -80659
rect -75924 -80703 -75916 -80659
rect -75824 -80703 -75816 -80659
rect -75724 -80703 -75716 -80659
rect -75624 -80703 -75616 -80659
rect -75524 -80703 -75516 -80659
rect -75424 -80703 -75416 -80659
rect -50017 -80661 -49973 -80653
rect -49917 -80661 -49873 -80653
rect -49817 -80661 -49773 -80653
rect -49717 -80661 -49673 -80653
rect -49617 -80661 -49573 -80653
rect -49517 -80661 -49473 -80653
rect -49417 -80661 -49373 -80653
rect -49317 -80661 -49273 -80653
rect -49217 -80661 -49173 -80653
rect -49117 -80661 -49073 -80653
rect -49017 -80661 -48973 -80653
rect -48917 -80661 -48873 -80653
rect -48817 -80661 -48773 -80653
rect -48717 -80661 -48673 -80653
rect -48617 -80661 -48573 -80653
rect -48517 -80661 -48473 -80653
rect -48017 -80661 -47973 -80653
rect -47917 -80661 -47873 -80653
rect -47817 -80661 -47773 -80653
rect -47717 -80661 -47673 -80653
rect -47617 -80661 -47573 -80653
rect -47517 -80661 -47473 -80653
rect -47417 -80661 -47373 -80653
rect -47317 -80661 -47273 -80653
rect -47217 -80661 -47173 -80653
rect -47117 -80661 -47073 -80653
rect -47017 -80661 -46973 -80653
rect -46917 -80661 -46873 -80653
rect -46817 -80661 -46773 -80653
rect -46717 -80661 -46673 -80653
rect -46617 -80661 -46573 -80653
rect -46517 -80661 -46473 -80653
rect -46017 -80661 -45973 -80653
rect -45917 -80661 -45873 -80653
rect -45817 -80661 -45773 -80653
rect -45717 -80661 -45673 -80653
rect -45617 -80661 -45573 -80653
rect -45517 -80661 -45473 -80653
rect -45417 -80661 -45373 -80653
rect -45317 -80661 -45273 -80653
rect -45217 -80661 -45173 -80653
rect -45117 -80661 -45073 -80653
rect -45017 -80661 -44973 -80653
rect -44917 -80661 -44873 -80653
rect -44817 -80661 -44773 -80653
rect -44717 -80661 -44673 -80653
rect -44617 -80661 -44573 -80653
rect -44517 -80661 -44473 -80653
rect -44017 -80661 -43973 -80653
rect -43917 -80661 -43873 -80653
rect -43817 -80661 -43773 -80653
rect -43717 -80661 -43673 -80653
rect -43617 -80661 -43573 -80653
rect -43517 -80661 -43473 -80653
rect -43417 -80661 -43373 -80653
rect -43317 -80661 -43273 -80653
rect -43217 -80661 -43173 -80653
rect -43117 -80661 -43073 -80653
rect -43017 -80661 -42973 -80653
rect -42917 -80661 -42873 -80653
rect -42817 -80661 -42773 -80653
rect -42717 -80661 -42673 -80653
rect -42617 -80661 -42573 -80653
rect -42517 -80661 -42473 -80653
rect 80737 -80655 80781 -80647
rect 80837 -80655 80881 -80647
rect 80937 -80655 80981 -80647
rect 81037 -80655 81081 -80647
rect 81137 -80655 81181 -80647
rect 81237 -80655 81281 -80647
rect 81337 -80655 81381 -80647
rect 81437 -80655 81481 -80647
rect 81537 -80655 81581 -80647
rect 81637 -80655 81681 -80647
rect 81737 -80655 81781 -80647
rect 81837 -80655 81881 -80647
rect 81937 -80655 81981 -80647
rect 82037 -80655 82081 -80647
rect 82137 -80655 82181 -80647
rect 82237 -80655 82281 -80647
rect 82737 -80655 82781 -80647
rect 82837 -80655 82881 -80647
rect 82937 -80655 82981 -80647
rect 83037 -80655 83081 -80647
rect 83137 -80655 83181 -80647
rect 83237 -80655 83281 -80647
rect 83337 -80655 83381 -80647
rect 83437 -80655 83481 -80647
rect 83537 -80655 83581 -80647
rect 83637 -80655 83681 -80647
rect 83737 -80655 83781 -80647
rect 83837 -80655 83881 -80647
rect 83937 -80655 83981 -80647
rect 84037 -80655 84081 -80647
rect 84137 -80655 84181 -80647
rect 84237 -80655 84281 -80647
rect 84737 -80655 84781 -80647
rect 84837 -80655 84881 -80647
rect 84937 -80655 84981 -80647
rect 85037 -80655 85081 -80647
rect 85137 -80655 85181 -80647
rect 85237 -80655 85281 -80647
rect 85337 -80655 85381 -80647
rect 85437 -80655 85481 -80647
rect 85537 -80655 85581 -80647
rect 85637 -80655 85681 -80647
rect 85737 -80655 85781 -80647
rect 85837 -80655 85881 -80647
rect 85937 -80655 85981 -80647
rect 86037 -80655 86081 -80647
rect 86137 -80655 86181 -80647
rect 86237 -80655 86281 -80647
rect 86737 -80655 86781 -80647
rect 86837 -80655 86881 -80647
rect 86937 -80655 86981 -80647
rect 87037 -80655 87081 -80647
rect 87137 -80655 87181 -80647
rect 87237 -80655 87281 -80647
rect 87337 -80655 87381 -80647
rect 87437 -80655 87481 -80647
rect 87537 -80655 87581 -80647
rect 87637 -80655 87681 -80647
rect 87737 -80655 87781 -80647
rect 87837 -80655 87881 -80647
rect 87937 -80655 87981 -80647
rect 88037 -80655 88081 -80647
rect 88137 -80655 88181 -80647
rect 88237 -80655 88281 -80647
rect -49973 -80705 -49965 -80661
rect -49873 -80705 -49865 -80661
rect -49773 -80705 -49765 -80661
rect -49673 -80705 -49665 -80661
rect -49573 -80705 -49565 -80661
rect -49473 -80705 -49465 -80661
rect -49373 -80705 -49365 -80661
rect -49273 -80705 -49265 -80661
rect -49173 -80705 -49165 -80661
rect -49073 -80705 -49065 -80661
rect -48973 -80705 -48965 -80661
rect -48873 -80705 -48865 -80661
rect -48773 -80705 -48765 -80661
rect -48673 -80705 -48665 -80661
rect -48573 -80705 -48565 -80661
rect -48473 -80705 -48465 -80661
rect -47973 -80705 -47965 -80661
rect -47873 -80705 -47865 -80661
rect -47773 -80705 -47765 -80661
rect -47673 -80705 -47665 -80661
rect -47573 -80705 -47565 -80661
rect -47473 -80705 -47465 -80661
rect -47373 -80705 -47365 -80661
rect -47273 -80705 -47265 -80661
rect -47173 -80705 -47165 -80661
rect -47073 -80705 -47065 -80661
rect -46973 -80705 -46965 -80661
rect -46873 -80705 -46865 -80661
rect -46773 -80705 -46765 -80661
rect -46673 -80705 -46665 -80661
rect -46573 -80705 -46565 -80661
rect -46473 -80705 -46465 -80661
rect -45973 -80705 -45965 -80661
rect -45873 -80705 -45865 -80661
rect -45773 -80705 -45765 -80661
rect -45673 -80705 -45665 -80661
rect -45573 -80705 -45565 -80661
rect -45473 -80705 -45465 -80661
rect -45373 -80705 -45365 -80661
rect -45273 -80705 -45265 -80661
rect -45173 -80705 -45165 -80661
rect -45073 -80705 -45065 -80661
rect -44973 -80705 -44965 -80661
rect -44873 -80705 -44865 -80661
rect -44773 -80705 -44765 -80661
rect -44673 -80705 -44665 -80661
rect -44573 -80705 -44565 -80661
rect -44473 -80705 -44465 -80661
rect -43973 -80705 -43965 -80661
rect -43873 -80705 -43865 -80661
rect -43773 -80705 -43765 -80661
rect -43673 -80705 -43665 -80661
rect -43573 -80705 -43565 -80661
rect -43473 -80705 -43465 -80661
rect -43373 -80705 -43365 -80661
rect -43273 -80705 -43265 -80661
rect -43173 -80705 -43165 -80661
rect -43073 -80705 -43065 -80661
rect -42973 -80705 -42965 -80661
rect -42873 -80705 -42865 -80661
rect -42773 -80705 -42765 -80661
rect -42673 -80705 -42665 -80661
rect -42573 -80705 -42565 -80661
rect -42473 -80705 -42465 -80661
rect 80781 -80699 80789 -80655
rect 80881 -80699 80889 -80655
rect 80981 -80699 80989 -80655
rect 81081 -80699 81089 -80655
rect 81181 -80699 81189 -80655
rect 81281 -80699 81289 -80655
rect 81381 -80699 81389 -80655
rect 81481 -80699 81489 -80655
rect 81581 -80699 81589 -80655
rect 81681 -80699 81689 -80655
rect 81781 -80699 81789 -80655
rect 81881 -80699 81889 -80655
rect 81981 -80699 81989 -80655
rect 82081 -80699 82089 -80655
rect 82181 -80699 82189 -80655
rect 82281 -80699 82289 -80655
rect 82781 -80699 82789 -80655
rect 82881 -80699 82889 -80655
rect 82981 -80699 82989 -80655
rect 83081 -80699 83089 -80655
rect 83181 -80699 83189 -80655
rect 83281 -80699 83289 -80655
rect 83381 -80699 83389 -80655
rect 83481 -80699 83489 -80655
rect 83581 -80699 83589 -80655
rect 83681 -80699 83689 -80655
rect 83781 -80699 83789 -80655
rect 83881 -80699 83889 -80655
rect 83981 -80699 83989 -80655
rect 84081 -80699 84089 -80655
rect 84181 -80699 84189 -80655
rect 84281 -80699 84289 -80655
rect 84781 -80699 84789 -80655
rect 84881 -80699 84889 -80655
rect 84981 -80699 84989 -80655
rect 85081 -80699 85089 -80655
rect 85181 -80699 85189 -80655
rect 85281 -80699 85289 -80655
rect 85381 -80699 85389 -80655
rect 85481 -80699 85489 -80655
rect 85581 -80699 85589 -80655
rect 85681 -80699 85689 -80655
rect 85781 -80699 85789 -80655
rect 85881 -80699 85889 -80655
rect 85981 -80699 85989 -80655
rect 86081 -80699 86089 -80655
rect 86181 -80699 86189 -80655
rect 86281 -80699 86289 -80655
rect 86781 -80699 86789 -80655
rect 86881 -80699 86889 -80655
rect 86981 -80699 86989 -80655
rect 87081 -80699 87089 -80655
rect 87181 -80699 87189 -80655
rect 87281 -80699 87289 -80655
rect 87381 -80699 87389 -80655
rect 87481 -80699 87489 -80655
rect 87581 -80699 87589 -80655
rect 87681 -80699 87689 -80655
rect 87781 -80699 87789 -80655
rect 87881 -80699 87889 -80655
rect 87981 -80699 87989 -80655
rect 88081 -80699 88089 -80655
rect 88181 -80699 88189 -80655
rect 88281 -80699 88289 -80655
rect -82968 -80759 -82924 -80751
rect -82868 -80759 -82824 -80751
rect -82768 -80759 -82724 -80751
rect -82668 -80759 -82624 -80751
rect -82568 -80759 -82524 -80751
rect -82468 -80759 -82424 -80751
rect -82368 -80759 -82324 -80751
rect -82268 -80759 -82224 -80751
rect -82168 -80759 -82124 -80751
rect -82068 -80759 -82024 -80751
rect -81968 -80759 -81924 -80751
rect -81868 -80759 -81824 -80751
rect -81768 -80759 -81724 -80751
rect -81668 -80759 -81624 -80751
rect -81568 -80759 -81524 -80751
rect -81468 -80759 -81424 -80751
rect -80968 -80759 -80924 -80751
rect -80868 -80759 -80824 -80751
rect -80768 -80759 -80724 -80751
rect -80668 -80759 -80624 -80751
rect -80568 -80759 -80524 -80751
rect -80468 -80759 -80424 -80751
rect -80368 -80759 -80324 -80751
rect -80268 -80759 -80224 -80751
rect -80168 -80759 -80124 -80751
rect -80068 -80759 -80024 -80751
rect -79968 -80759 -79924 -80751
rect -79868 -80759 -79824 -80751
rect -79768 -80759 -79724 -80751
rect -79668 -80759 -79624 -80751
rect -79568 -80759 -79524 -80751
rect -79468 -80759 -79424 -80751
rect -78968 -80759 -78924 -80751
rect -78868 -80759 -78824 -80751
rect -78768 -80759 -78724 -80751
rect -78668 -80759 -78624 -80751
rect -78568 -80759 -78524 -80751
rect -78468 -80759 -78424 -80751
rect -78368 -80759 -78324 -80751
rect -78268 -80759 -78224 -80751
rect -78168 -80759 -78124 -80751
rect -78068 -80759 -78024 -80751
rect -77968 -80759 -77924 -80751
rect -77868 -80759 -77824 -80751
rect -77768 -80759 -77724 -80751
rect -77668 -80759 -77624 -80751
rect -77568 -80759 -77524 -80751
rect -77468 -80759 -77424 -80751
rect -76968 -80759 -76924 -80751
rect -76868 -80759 -76824 -80751
rect -76768 -80759 -76724 -80751
rect -76668 -80759 -76624 -80751
rect -76568 -80759 -76524 -80751
rect -76468 -80759 -76424 -80751
rect -76368 -80759 -76324 -80751
rect -76268 -80759 -76224 -80751
rect -76168 -80759 -76124 -80751
rect -76068 -80759 -76024 -80751
rect -75968 -80759 -75924 -80751
rect -75868 -80759 -75824 -80751
rect -75768 -80759 -75724 -80751
rect -75668 -80759 -75624 -80751
rect -75568 -80759 -75524 -80751
rect -75468 -80759 -75424 -80751
rect -82924 -80803 -82916 -80759
rect -82824 -80803 -82816 -80759
rect -82724 -80803 -82716 -80759
rect -82624 -80803 -82616 -80759
rect -82524 -80803 -82516 -80759
rect -82424 -80803 -82416 -80759
rect -82324 -80803 -82316 -80759
rect -82224 -80803 -82216 -80759
rect -82124 -80803 -82116 -80759
rect -82024 -80803 -82016 -80759
rect -81924 -80803 -81916 -80759
rect -81824 -80803 -81816 -80759
rect -81724 -80803 -81716 -80759
rect -81624 -80803 -81616 -80759
rect -81524 -80803 -81516 -80759
rect -81424 -80803 -81416 -80759
rect -80924 -80803 -80916 -80759
rect -80824 -80803 -80816 -80759
rect -80724 -80803 -80716 -80759
rect -80624 -80803 -80616 -80759
rect -80524 -80803 -80516 -80759
rect -80424 -80803 -80416 -80759
rect -80324 -80803 -80316 -80759
rect -80224 -80803 -80216 -80759
rect -80124 -80803 -80116 -80759
rect -80024 -80803 -80016 -80759
rect -79924 -80803 -79916 -80759
rect -79824 -80803 -79816 -80759
rect -79724 -80803 -79716 -80759
rect -79624 -80803 -79616 -80759
rect -79524 -80803 -79516 -80759
rect -79424 -80803 -79416 -80759
rect -78924 -80803 -78916 -80759
rect -78824 -80803 -78816 -80759
rect -78724 -80803 -78716 -80759
rect -78624 -80803 -78616 -80759
rect -78524 -80803 -78516 -80759
rect -78424 -80803 -78416 -80759
rect -78324 -80803 -78316 -80759
rect -78224 -80803 -78216 -80759
rect -78124 -80803 -78116 -80759
rect -78024 -80803 -78016 -80759
rect -77924 -80803 -77916 -80759
rect -77824 -80803 -77816 -80759
rect -77724 -80803 -77716 -80759
rect -77624 -80803 -77616 -80759
rect -77524 -80803 -77516 -80759
rect -77424 -80803 -77416 -80759
rect -76924 -80803 -76916 -80759
rect -76824 -80803 -76816 -80759
rect -76724 -80803 -76716 -80759
rect -76624 -80803 -76616 -80759
rect -76524 -80803 -76516 -80759
rect -76424 -80803 -76416 -80759
rect -76324 -80803 -76316 -80759
rect -76224 -80803 -76216 -80759
rect -76124 -80803 -76116 -80759
rect -76024 -80803 -76016 -80759
rect -75924 -80803 -75916 -80759
rect -75824 -80803 -75816 -80759
rect -75724 -80803 -75716 -80759
rect -75624 -80803 -75616 -80759
rect -75524 -80803 -75516 -80759
rect -75424 -80803 -75416 -80759
rect -50017 -80761 -49973 -80753
rect -49917 -80761 -49873 -80753
rect -49817 -80761 -49773 -80753
rect -49717 -80761 -49673 -80753
rect -49617 -80761 -49573 -80753
rect -49517 -80761 -49473 -80753
rect -49417 -80761 -49373 -80753
rect -49317 -80761 -49273 -80753
rect -49217 -80761 -49173 -80753
rect -49117 -80761 -49073 -80753
rect -49017 -80761 -48973 -80753
rect -48917 -80761 -48873 -80753
rect -48817 -80761 -48773 -80753
rect -48717 -80761 -48673 -80753
rect -48617 -80761 -48573 -80753
rect -48517 -80761 -48473 -80753
rect -48017 -80761 -47973 -80753
rect -47917 -80761 -47873 -80753
rect -47817 -80761 -47773 -80753
rect -47717 -80761 -47673 -80753
rect -47617 -80761 -47573 -80753
rect -47517 -80761 -47473 -80753
rect -47417 -80761 -47373 -80753
rect -47317 -80761 -47273 -80753
rect -47217 -80761 -47173 -80753
rect -47117 -80761 -47073 -80753
rect -47017 -80761 -46973 -80753
rect -46917 -80761 -46873 -80753
rect -46817 -80761 -46773 -80753
rect -46717 -80761 -46673 -80753
rect -46617 -80761 -46573 -80753
rect -46517 -80761 -46473 -80753
rect -46017 -80761 -45973 -80753
rect -45917 -80761 -45873 -80753
rect -45817 -80761 -45773 -80753
rect -45717 -80761 -45673 -80753
rect -45617 -80761 -45573 -80753
rect -45517 -80761 -45473 -80753
rect -45417 -80761 -45373 -80753
rect -45317 -80761 -45273 -80753
rect -45217 -80761 -45173 -80753
rect -45117 -80761 -45073 -80753
rect -45017 -80761 -44973 -80753
rect -44917 -80761 -44873 -80753
rect -44817 -80761 -44773 -80753
rect -44717 -80761 -44673 -80753
rect -44617 -80761 -44573 -80753
rect -44517 -80761 -44473 -80753
rect -44017 -80761 -43973 -80753
rect -43917 -80761 -43873 -80753
rect -43817 -80761 -43773 -80753
rect -43717 -80761 -43673 -80753
rect -43617 -80761 -43573 -80753
rect -43517 -80761 -43473 -80753
rect -43417 -80761 -43373 -80753
rect -43317 -80761 -43273 -80753
rect -43217 -80761 -43173 -80753
rect -43117 -80761 -43073 -80753
rect -43017 -80761 -42973 -80753
rect -42917 -80761 -42873 -80753
rect -42817 -80761 -42773 -80753
rect -42717 -80761 -42673 -80753
rect -42617 -80761 -42573 -80753
rect -42517 -80761 -42473 -80753
rect 80737 -80755 80781 -80747
rect 80837 -80755 80881 -80747
rect 80937 -80755 80981 -80747
rect 81037 -80755 81081 -80747
rect 81137 -80755 81181 -80747
rect 81237 -80755 81281 -80747
rect 81337 -80755 81381 -80747
rect 81437 -80755 81481 -80747
rect 81537 -80755 81581 -80747
rect 81637 -80755 81681 -80747
rect 81737 -80755 81781 -80747
rect 81837 -80755 81881 -80747
rect 81937 -80755 81981 -80747
rect 82037 -80755 82081 -80747
rect 82137 -80755 82181 -80747
rect 82237 -80755 82281 -80747
rect 82737 -80755 82781 -80747
rect 82837 -80755 82881 -80747
rect 82937 -80755 82981 -80747
rect 83037 -80755 83081 -80747
rect 83137 -80755 83181 -80747
rect 83237 -80755 83281 -80747
rect 83337 -80755 83381 -80747
rect 83437 -80755 83481 -80747
rect 83537 -80755 83581 -80747
rect 83637 -80755 83681 -80747
rect 83737 -80755 83781 -80747
rect 83837 -80755 83881 -80747
rect 83937 -80755 83981 -80747
rect 84037 -80755 84081 -80747
rect 84137 -80755 84181 -80747
rect 84237 -80755 84281 -80747
rect 84737 -80755 84781 -80747
rect 84837 -80755 84881 -80747
rect 84937 -80755 84981 -80747
rect 85037 -80755 85081 -80747
rect 85137 -80755 85181 -80747
rect 85237 -80755 85281 -80747
rect 85337 -80755 85381 -80747
rect 85437 -80755 85481 -80747
rect 85537 -80755 85581 -80747
rect 85637 -80755 85681 -80747
rect 85737 -80755 85781 -80747
rect 85837 -80755 85881 -80747
rect 85937 -80755 85981 -80747
rect 86037 -80755 86081 -80747
rect 86137 -80755 86181 -80747
rect 86237 -80755 86281 -80747
rect 86737 -80755 86781 -80747
rect 86837 -80755 86881 -80747
rect 86937 -80755 86981 -80747
rect 87037 -80755 87081 -80747
rect 87137 -80755 87181 -80747
rect 87237 -80755 87281 -80747
rect 87337 -80755 87381 -80747
rect 87437 -80755 87481 -80747
rect 87537 -80755 87581 -80747
rect 87637 -80755 87681 -80747
rect 87737 -80755 87781 -80747
rect 87837 -80755 87881 -80747
rect 87937 -80755 87981 -80747
rect 88037 -80755 88081 -80747
rect 88137 -80755 88181 -80747
rect 88237 -80755 88281 -80747
rect -49973 -80805 -49965 -80761
rect -49873 -80805 -49865 -80761
rect -49773 -80805 -49765 -80761
rect -49673 -80805 -49665 -80761
rect -49573 -80805 -49565 -80761
rect -49473 -80805 -49465 -80761
rect -49373 -80805 -49365 -80761
rect -49273 -80805 -49265 -80761
rect -49173 -80805 -49165 -80761
rect -49073 -80805 -49065 -80761
rect -48973 -80805 -48965 -80761
rect -48873 -80805 -48865 -80761
rect -48773 -80805 -48765 -80761
rect -48673 -80805 -48665 -80761
rect -48573 -80805 -48565 -80761
rect -48473 -80805 -48465 -80761
rect -47973 -80805 -47965 -80761
rect -47873 -80805 -47865 -80761
rect -47773 -80805 -47765 -80761
rect -47673 -80805 -47665 -80761
rect -47573 -80805 -47565 -80761
rect -47473 -80805 -47465 -80761
rect -47373 -80805 -47365 -80761
rect -47273 -80805 -47265 -80761
rect -47173 -80805 -47165 -80761
rect -47073 -80805 -47065 -80761
rect -46973 -80805 -46965 -80761
rect -46873 -80805 -46865 -80761
rect -46773 -80805 -46765 -80761
rect -46673 -80805 -46665 -80761
rect -46573 -80805 -46565 -80761
rect -46473 -80805 -46465 -80761
rect -45973 -80805 -45965 -80761
rect -45873 -80805 -45865 -80761
rect -45773 -80805 -45765 -80761
rect -45673 -80805 -45665 -80761
rect -45573 -80805 -45565 -80761
rect -45473 -80805 -45465 -80761
rect -45373 -80805 -45365 -80761
rect -45273 -80805 -45265 -80761
rect -45173 -80805 -45165 -80761
rect -45073 -80805 -45065 -80761
rect -44973 -80805 -44965 -80761
rect -44873 -80805 -44865 -80761
rect -44773 -80805 -44765 -80761
rect -44673 -80805 -44665 -80761
rect -44573 -80805 -44565 -80761
rect -44473 -80805 -44465 -80761
rect -43973 -80805 -43965 -80761
rect -43873 -80805 -43865 -80761
rect -43773 -80805 -43765 -80761
rect -43673 -80805 -43665 -80761
rect -43573 -80805 -43565 -80761
rect -43473 -80805 -43465 -80761
rect -43373 -80805 -43365 -80761
rect -43273 -80805 -43265 -80761
rect -43173 -80805 -43165 -80761
rect -43073 -80805 -43065 -80761
rect -42973 -80805 -42965 -80761
rect -42873 -80805 -42865 -80761
rect -42773 -80805 -42765 -80761
rect -42673 -80805 -42665 -80761
rect -42573 -80805 -42565 -80761
rect -42473 -80805 -42465 -80761
rect 80781 -80799 80789 -80755
rect 80881 -80799 80889 -80755
rect 80981 -80799 80989 -80755
rect 81081 -80799 81089 -80755
rect 81181 -80799 81189 -80755
rect 81281 -80799 81289 -80755
rect 81381 -80799 81389 -80755
rect 81481 -80799 81489 -80755
rect 81581 -80799 81589 -80755
rect 81681 -80799 81689 -80755
rect 81781 -80799 81789 -80755
rect 81881 -80799 81889 -80755
rect 81981 -80799 81989 -80755
rect 82081 -80799 82089 -80755
rect 82181 -80799 82189 -80755
rect 82281 -80799 82289 -80755
rect 82781 -80799 82789 -80755
rect 82881 -80799 82889 -80755
rect 82981 -80799 82989 -80755
rect 83081 -80799 83089 -80755
rect 83181 -80799 83189 -80755
rect 83281 -80799 83289 -80755
rect 83381 -80799 83389 -80755
rect 83481 -80799 83489 -80755
rect 83581 -80799 83589 -80755
rect 83681 -80799 83689 -80755
rect 83781 -80799 83789 -80755
rect 83881 -80799 83889 -80755
rect 83981 -80799 83989 -80755
rect 84081 -80799 84089 -80755
rect 84181 -80799 84189 -80755
rect 84281 -80799 84289 -80755
rect 84781 -80799 84789 -80755
rect 84881 -80799 84889 -80755
rect 84981 -80799 84989 -80755
rect 85081 -80799 85089 -80755
rect 85181 -80799 85189 -80755
rect 85281 -80799 85289 -80755
rect 85381 -80799 85389 -80755
rect 85481 -80799 85489 -80755
rect 85581 -80799 85589 -80755
rect 85681 -80799 85689 -80755
rect 85781 -80799 85789 -80755
rect 85881 -80799 85889 -80755
rect 85981 -80799 85989 -80755
rect 86081 -80799 86089 -80755
rect 86181 -80799 86189 -80755
rect 86281 -80799 86289 -80755
rect 86781 -80799 86789 -80755
rect 86881 -80799 86889 -80755
rect 86981 -80799 86989 -80755
rect 87081 -80799 87089 -80755
rect 87181 -80799 87189 -80755
rect 87281 -80799 87289 -80755
rect 87381 -80799 87389 -80755
rect 87481 -80799 87489 -80755
rect 87581 -80799 87589 -80755
rect 87681 -80799 87689 -80755
rect 87781 -80799 87789 -80755
rect 87881 -80799 87889 -80755
rect 87981 -80799 87989 -80755
rect 88081 -80799 88089 -80755
rect 88181 -80799 88189 -80755
rect 88281 -80799 88289 -80755
rect -82968 -80859 -82924 -80851
rect -82868 -80859 -82824 -80851
rect -82768 -80859 -82724 -80851
rect -82668 -80859 -82624 -80851
rect -82568 -80859 -82524 -80851
rect -82468 -80859 -82424 -80851
rect -82368 -80859 -82324 -80851
rect -82268 -80859 -82224 -80851
rect -82168 -80859 -82124 -80851
rect -82068 -80859 -82024 -80851
rect -81968 -80859 -81924 -80851
rect -81868 -80859 -81824 -80851
rect -81768 -80859 -81724 -80851
rect -81668 -80859 -81624 -80851
rect -81568 -80859 -81524 -80851
rect -81468 -80859 -81424 -80851
rect -80968 -80859 -80924 -80851
rect -80868 -80859 -80824 -80851
rect -80768 -80859 -80724 -80851
rect -80668 -80859 -80624 -80851
rect -80568 -80859 -80524 -80851
rect -80468 -80859 -80424 -80851
rect -80368 -80859 -80324 -80851
rect -80268 -80859 -80224 -80851
rect -80168 -80859 -80124 -80851
rect -80068 -80859 -80024 -80851
rect -79968 -80859 -79924 -80851
rect -79868 -80859 -79824 -80851
rect -79768 -80859 -79724 -80851
rect -79668 -80859 -79624 -80851
rect -79568 -80859 -79524 -80851
rect -79468 -80859 -79424 -80851
rect -78968 -80859 -78924 -80851
rect -78868 -80859 -78824 -80851
rect -78768 -80859 -78724 -80851
rect -78668 -80859 -78624 -80851
rect -78568 -80859 -78524 -80851
rect -78468 -80859 -78424 -80851
rect -78368 -80859 -78324 -80851
rect -78268 -80859 -78224 -80851
rect -78168 -80859 -78124 -80851
rect -78068 -80859 -78024 -80851
rect -77968 -80859 -77924 -80851
rect -77868 -80859 -77824 -80851
rect -77768 -80859 -77724 -80851
rect -77668 -80859 -77624 -80851
rect -77568 -80859 -77524 -80851
rect -77468 -80859 -77424 -80851
rect -76968 -80859 -76924 -80851
rect -76868 -80859 -76824 -80851
rect -76768 -80859 -76724 -80851
rect -76668 -80859 -76624 -80851
rect -76568 -80859 -76524 -80851
rect -76468 -80859 -76424 -80851
rect -76368 -80859 -76324 -80851
rect -76268 -80859 -76224 -80851
rect -76168 -80859 -76124 -80851
rect -76068 -80859 -76024 -80851
rect -75968 -80859 -75924 -80851
rect -75868 -80859 -75824 -80851
rect -75768 -80859 -75724 -80851
rect -75668 -80859 -75624 -80851
rect -75568 -80859 -75524 -80851
rect -75468 -80859 -75424 -80851
rect -82924 -80903 -82916 -80859
rect -82824 -80903 -82816 -80859
rect -82724 -80903 -82716 -80859
rect -82624 -80903 -82616 -80859
rect -82524 -80903 -82516 -80859
rect -82424 -80903 -82416 -80859
rect -82324 -80903 -82316 -80859
rect -82224 -80903 -82216 -80859
rect -82124 -80903 -82116 -80859
rect -82024 -80903 -82016 -80859
rect -81924 -80903 -81916 -80859
rect -81824 -80903 -81816 -80859
rect -81724 -80903 -81716 -80859
rect -81624 -80903 -81616 -80859
rect -81524 -80903 -81516 -80859
rect -81424 -80903 -81416 -80859
rect -80924 -80903 -80916 -80859
rect -80824 -80903 -80816 -80859
rect -80724 -80903 -80716 -80859
rect -80624 -80903 -80616 -80859
rect -80524 -80903 -80516 -80859
rect -80424 -80903 -80416 -80859
rect -80324 -80903 -80316 -80859
rect -80224 -80903 -80216 -80859
rect -80124 -80903 -80116 -80859
rect -80024 -80903 -80016 -80859
rect -79924 -80903 -79916 -80859
rect -79824 -80903 -79816 -80859
rect -79724 -80903 -79716 -80859
rect -79624 -80903 -79616 -80859
rect -79524 -80903 -79516 -80859
rect -79424 -80903 -79416 -80859
rect -78924 -80903 -78916 -80859
rect -78824 -80903 -78816 -80859
rect -78724 -80903 -78716 -80859
rect -78624 -80903 -78616 -80859
rect -78524 -80903 -78516 -80859
rect -78424 -80903 -78416 -80859
rect -78324 -80903 -78316 -80859
rect -78224 -80903 -78216 -80859
rect -78124 -80903 -78116 -80859
rect -78024 -80903 -78016 -80859
rect -77924 -80903 -77916 -80859
rect -77824 -80903 -77816 -80859
rect -77724 -80903 -77716 -80859
rect -77624 -80903 -77616 -80859
rect -77524 -80903 -77516 -80859
rect -77424 -80903 -77416 -80859
rect -76924 -80903 -76916 -80859
rect -76824 -80903 -76816 -80859
rect -76724 -80903 -76716 -80859
rect -76624 -80903 -76616 -80859
rect -76524 -80903 -76516 -80859
rect -76424 -80903 -76416 -80859
rect -76324 -80903 -76316 -80859
rect -76224 -80903 -76216 -80859
rect -76124 -80903 -76116 -80859
rect -76024 -80903 -76016 -80859
rect -75924 -80903 -75916 -80859
rect -75824 -80903 -75816 -80859
rect -75724 -80903 -75716 -80859
rect -75624 -80903 -75616 -80859
rect -75524 -80903 -75516 -80859
rect -75424 -80903 -75416 -80859
rect -50017 -80861 -49973 -80853
rect -49917 -80861 -49873 -80853
rect -49817 -80861 -49773 -80853
rect -49717 -80861 -49673 -80853
rect -49617 -80861 -49573 -80853
rect -49517 -80861 -49473 -80853
rect -49417 -80861 -49373 -80853
rect -49317 -80861 -49273 -80853
rect -49217 -80861 -49173 -80853
rect -49117 -80861 -49073 -80853
rect -49017 -80861 -48973 -80853
rect -48917 -80861 -48873 -80853
rect -48817 -80861 -48773 -80853
rect -48717 -80861 -48673 -80853
rect -48617 -80861 -48573 -80853
rect -48517 -80861 -48473 -80853
rect -48017 -80861 -47973 -80853
rect -47917 -80861 -47873 -80853
rect -47817 -80861 -47773 -80853
rect -47717 -80861 -47673 -80853
rect -47617 -80861 -47573 -80853
rect -47517 -80861 -47473 -80853
rect -47417 -80861 -47373 -80853
rect -47317 -80861 -47273 -80853
rect -47217 -80861 -47173 -80853
rect -47117 -80861 -47073 -80853
rect -47017 -80861 -46973 -80853
rect -46917 -80861 -46873 -80853
rect -46817 -80861 -46773 -80853
rect -46717 -80861 -46673 -80853
rect -46617 -80861 -46573 -80853
rect -46517 -80861 -46473 -80853
rect -46017 -80861 -45973 -80853
rect -45917 -80861 -45873 -80853
rect -45817 -80861 -45773 -80853
rect -45717 -80861 -45673 -80853
rect -45617 -80861 -45573 -80853
rect -45517 -80861 -45473 -80853
rect -45417 -80861 -45373 -80853
rect -45317 -80861 -45273 -80853
rect -45217 -80861 -45173 -80853
rect -45117 -80861 -45073 -80853
rect -45017 -80861 -44973 -80853
rect -44917 -80861 -44873 -80853
rect -44817 -80861 -44773 -80853
rect -44717 -80861 -44673 -80853
rect -44617 -80861 -44573 -80853
rect -44517 -80861 -44473 -80853
rect -44017 -80861 -43973 -80853
rect -43917 -80861 -43873 -80853
rect -43817 -80861 -43773 -80853
rect -43717 -80861 -43673 -80853
rect -43617 -80861 -43573 -80853
rect -43517 -80861 -43473 -80853
rect -43417 -80861 -43373 -80853
rect -43317 -80861 -43273 -80853
rect -43217 -80861 -43173 -80853
rect -43117 -80861 -43073 -80853
rect -43017 -80861 -42973 -80853
rect -42917 -80861 -42873 -80853
rect -42817 -80861 -42773 -80853
rect -42717 -80861 -42673 -80853
rect -42617 -80861 -42573 -80853
rect -42517 -80861 -42473 -80853
rect 80737 -80855 80781 -80847
rect 80837 -80855 80881 -80847
rect 80937 -80855 80981 -80847
rect 81037 -80855 81081 -80847
rect 81137 -80855 81181 -80847
rect 81237 -80855 81281 -80847
rect 81337 -80855 81381 -80847
rect 81437 -80855 81481 -80847
rect 81537 -80855 81581 -80847
rect 81637 -80855 81681 -80847
rect 81737 -80855 81781 -80847
rect 81837 -80855 81881 -80847
rect 81937 -80855 81981 -80847
rect 82037 -80855 82081 -80847
rect 82137 -80855 82181 -80847
rect 82237 -80855 82281 -80847
rect 82737 -80855 82781 -80847
rect 82837 -80855 82881 -80847
rect 82937 -80855 82981 -80847
rect 83037 -80855 83081 -80847
rect 83137 -80855 83181 -80847
rect 83237 -80855 83281 -80847
rect 83337 -80855 83381 -80847
rect 83437 -80855 83481 -80847
rect 83537 -80855 83581 -80847
rect 83637 -80855 83681 -80847
rect 83737 -80855 83781 -80847
rect 83837 -80855 83881 -80847
rect 83937 -80855 83981 -80847
rect 84037 -80855 84081 -80847
rect 84137 -80855 84181 -80847
rect 84237 -80855 84281 -80847
rect 84737 -80855 84781 -80847
rect 84837 -80855 84881 -80847
rect 84937 -80855 84981 -80847
rect 85037 -80855 85081 -80847
rect 85137 -80855 85181 -80847
rect 85237 -80855 85281 -80847
rect 85337 -80855 85381 -80847
rect 85437 -80855 85481 -80847
rect 85537 -80855 85581 -80847
rect 85637 -80855 85681 -80847
rect 85737 -80855 85781 -80847
rect 85837 -80855 85881 -80847
rect 85937 -80855 85981 -80847
rect 86037 -80855 86081 -80847
rect 86137 -80855 86181 -80847
rect 86237 -80855 86281 -80847
rect 86737 -80855 86781 -80847
rect 86837 -80855 86881 -80847
rect 86937 -80855 86981 -80847
rect 87037 -80855 87081 -80847
rect 87137 -80855 87181 -80847
rect 87237 -80855 87281 -80847
rect 87337 -80855 87381 -80847
rect 87437 -80855 87481 -80847
rect 87537 -80855 87581 -80847
rect 87637 -80855 87681 -80847
rect 87737 -80855 87781 -80847
rect 87837 -80855 87881 -80847
rect 87937 -80855 87981 -80847
rect 88037 -80855 88081 -80847
rect 88137 -80855 88181 -80847
rect 88237 -80855 88281 -80847
rect -49973 -80905 -49965 -80861
rect -49873 -80905 -49865 -80861
rect -49773 -80905 -49765 -80861
rect -49673 -80905 -49665 -80861
rect -49573 -80905 -49565 -80861
rect -49473 -80905 -49465 -80861
rect -49373 -80905 -49365 -80861
rect -49273 -80905 -49265 -80861
rect -49173 -80905 -49165 -80861
rect -49073 -80905 -49065 -80861
rect -48973 -80905 -48965 -80861
rect -48873 -80905 -48865 -80861
rect -48773 -80905 -48765 -80861
rect -48673 -80905 -48665 -80861
rect -48573 -80905 -48565 -80861
rect -48473 -80905 -48465 -80861
rect -47973 -80905 -47965 -80861
rect -47873 -80905 -47865 -80861
rect -47773 -80905 -47765 -80861
rect -47673 -80905 -47665 -80861
rect -47573 -80905 -47565 -80861
rect -47473 -80905 -47465 -80861
rect -47373 -80905 -47365 -80861
rect -47273 -80905 -47265 -80861
rect -47173 -80905 -47165 -80861
rect -47073 -80905 -47065 -80861
rect -46973 -80905 -46965 -80861
rect -46873 -80905 -46865 -80861
rect -46773 -80905 -46765 -80861
rect -46673 -80905 -46665 -80861
rect -46573 -80905 -46565 -80861
rect -46473 -80905 -46465 -80861
rect -45973 -80905 -45965 -80861
rect -45873 -80905 -45865 -80861
rect -45773 -80905 -45765 -80861
rect -45673 -80905 -45665 -80861
rect -45573 -80905 -45565 -80861
rect -45473 -80905 -45465 -80861
rect -45373 -80905 -45365 -80861
rect -45273 -80905 -45265 -80861
rect -45173 -80905 -45165 -80861
rect -45073 -80905 -45065 -80861
rect -44973 -80905 -44965 -80861
rect -44873 -80905 -44865 -80861
rect -44773 -80905 -44765 -80861
rect -44673 -80905 -44665 -80861
rect -44573 -80905 -44565 -80861
rect -44473 -80905 -44465 -80861
rect -43973 -80905 -43965 -80861
rect -43873 -80905 -43865 -80861
rect -43773 -80905 -43765 -80861
rect -43673 -80905 -43665 -80861
rect -43573 -80905 -43565 -80861
rect -43473 -80905 -43465 -80861
rect -43373 -80905 -43365 -80861
rect -43273 -80905 -43265 -80861
rect -43173 -80905 -43165 -80861
rect -43073 -80905 -43065 -80861
rect -42973 -80905 -42965 -80861
rect -42873 -80905 -42865 -80861
rect -42773 -80905 -42765 -80861
rect -42673 -80905 -42665 -80861
rect -42573 -80905 -42565 -80861
rect -42473 -80905 -42465 -80861
rect 80781 -80899 80789 -80855
rect 80881 -80899 80889 -80855
rect 80981 -80899 80989 -80855
rect 81081 -80899 81089 -80855
rect 81181 -80899 81189 -80855
rect 81281 -80899 81289 -80855
rect 81381 -80899 81389 -80855
rect 81481 -80899 81489 -80855
rect 81581 -80899 81589 -80855
rect 81681 -80899 81689 -80855
rect 81781 -80899 81789 -80855
rect 81881 -80899 81889 -80855
rect 81981 -80899 81989 -80855
rect 82081 -80899 82089 -80855
rect 82181 -80899 82189 -80855
rect 82281 -80899 82289 -80855
rect 82781 -80899 82789 -80855
rect 82881 -80899 82889 -80855
rect 82981 -80899 82989 -80855
rect 83081 -80899 83089 -80855
rect 83181 -80899 83189 -80855
rect 83281 -80899 83289 -80855
rect 83381 -80899 83389 -80855
rect 83481 -80899 83489 -80855
rect 83581 -80899 83589 -80855
rect 83681 -80899 83689 -80855
rect 83781 -80899 83789 -80855
rect 83881 -80899 83889 -80855
rect 83981 -80899 83989 -80855
rect 84081 -80899 84089 -80855
rect 84181 -80899 84189 -80855
rect 84281 -80899 84289 -80855
rect 84781 -80899 84789 -80855
rect 84881 -80899 84889 -80855
rect 84981 -80899 84989 -80855
rect 85081 -80899 85089 -80855
rect 85181 -80899 85189 -80855
rect 85281 -80899 85289 -80855
rect 85381 -80899 85389 -80855
rect 85481 -80899 85489 -80855
rect 85581 -80899 85589 -80855
rect 85681 -80899 85689 -80855
rect 85781 -80899 85789 -80855
rect 85881 -80899 85889 -80855
rect 85981 -80899 85989 -80855
rect 86081 -80899 86089 -80855
rect 86181 -80899 86189 -80855
rect 86281 -80899 86289 -80855
rect 86781 -80899 86789 -80855
rect 86881 -80899 86889 -80855
rect 86981 -80899 86989 -80855
rect 87081 -80899 87089 -80855
rect 87181 -80899 87189 -80855
rect 87281 -80899 87289 -80855
rect 87381 -80899 87389 -80855
rect 87481 -80899 87489 -80855
rect 87581 -80899 87589 -80855
rect 87681 -80899 87689 -80855
rect 87781 -80899 87789 -80855
rect 87881 -80899 87889 -80855
rect 87981 -80899 87989 -80855
rect 88081 -80899 88089 -80855
rect 88181 -80899 88189 -80855
rect 88281 -80899 88289 -80855
rect -82968 -80959 -82924 -80951
rect -82868 -80959 -82824 -80951
rect -82768 -80959 -82724 -80951
rect -82668 -80959 -82624 -80951
rect -82568 -80959 -82524 -80951
rect -82468 -80959 -82424 -80951
rect -82368 -80959 -82324 -80951
rect -82268 -80959 -82224 -80951
rect -82168 -80959 -82124 -80951
rect -82068 -80959 -82024 -80951
rect -81968 -80959 -81924 -80951
rect -81868 -80959 -81824 -80951
rect -81768 -80959 -81724 -80951
rect -81668 -80959 -81624 -80951
rect -81568 -80959 -81524 -80951
rect -81468 -80959 -81424 -80951
rect -80968 -80959 -80924 -80951
rect -80868 -80959 -80824 -80951
rect -80768 -80959 -80724 -80951
rect -80668 -80959 -80624 -80951
rect -80568 -80959 -80524 -80951
rect -80468 -80959 -80424 -80951
rect -80368 -80959 -80324 -80951
rect -80268 -80959 -80224 -80951
rect -80168 -80959 -80124 -80951
rect -80068 -80959 -80024 -80951
rect -79968 -80959 -79924 -80951
rect -79868 -80959 -79824 -80951
rect -79768 -80959 -79724 -80951
rect -79668 -80959 -79624 -80951
rect -79568 -80959 -79524 -80951
rect -79468 -80959 -79424 -80951
rect -78968 -80959 -78924 -80951
rect -78868 -80959 -78824 -80951
rect -78768 -80959 -78724 -80951
rect -78668 -80959 -78624 -80951
rect -78568 -80959 -78524 -80951
rect -78468 -80959 -78424 -80951
rect -78368 -80959 -78324 -80951
rect -78268 -80959 -78224 -80951
rect -78168 -80959 -78124 -80951
rect -78068 -80959 -78024 -80951
rect -77968 -80959 -77924 -80951
rect -77868 -80959 -77824 -80951
rect -77768 -80959 -77724 -80951
rect -77668 -80959 -77624 -80951
rect -77568 -80959 -77524 -80951
rect -77468 -80959 -77424 -80951
rect -76968 -80959 -76924 -80951
rect -76868 -80959 -76824 -80951
rect -76768 -80959 -76724 -80951
rect -76668 -80959 -76624 -80951
rect -76568 -80959 -76524 -80951
rect -76468 -80959 -76424 -80951
rect -76368 -80959 -76324 -80951
rect -76268 -80959 -76224 -80951
rect -76168 -80959 -76124 -80951
rect -76068 -80959 -76024 -80951
rect -75968 -80959 -75924 -80951
rect -75868 -80959 -75824 -80951
rect -75768 -80959 -75724 -80951
rect -75668 -80959 -75624 -80951
rect -75568 -80959 -75524 -80951
rect -75468 -80959 -75424 -80951
rect -82924 -81003 -82916 -80959
rect -82824 -81003 -82816 -80959
rect -82724 -81003 -82716 -80959
rect -82624 -81003 -82616 -80959
rect -82524 -81003 -82516 -80959
rect -82424 -81003 -82416 -80959
rect -82324 -81003 -82316 -80959
rect -82224 -81003 -82216 -80959
rect -82124 -81003 -82116 -80959
rect -82024 -81003 -82016 -80959
rect -81924 -81003 -81916 -80959
rect -81824 -81003 -81816 -80959
rect -81724 -81003 -81716 -80959
rect -81624 -81003 -81616 -80959
rect -81524 -81003 -81516 -80959
rect -81424 -81003 -81416 -80959
rect -80924 -81003 -80916 -80959
rect -80824 -81003 -80816 -80959
rect -80724 -81003 -80716 -80959
rect -80624 -81003 -80616 -80959
rect -80524 -81003 -80516 -80959
rect -80424 -81003 -80416 -80959
rect -80324 -81003 -80316 -80959
rect -80224 -81003 -80216 -80959
rect -80124 -81003 -80116 -80959
rect -80024 -81003 -80016 -80959
rect -79924 -81003 -79916 -80959
rect -79824 -81003 -79816 -80959
rect -79724 -81003 -79716 -80959
rect -79624 -81003 -79616 -80959
rect -79524 -81003 -79516 -80959
rect -79424 -81003 -79416 -80959
rect -78924 -81003 -78916 -80959
rect -78824 -81003 -78816 -80959
rect -78724 -81003 -78716 -80959
rect -78624 -81003 -78616 -80959
rect -78524 -81003 -78516 -80959
rect -78424 -81003 -78416 -80959
rect -78324 -81003 -78316 -80959
rect -78224 -81003 -78216 -80959
rect -78124 -81003 -78116 -80959
rect -78024 -81003 -78016 -80959
rect -77924 -81003 -77916 -80959
rect -77824 -81003 -77816 -80959
rect -77724 -81003 -77716 -80959
rect -77624 -81003 -77616 -80959
rect -77524 -81003 -77516 -80959
rect -77424 -81003 -77416 -80959
rect -76924 -81003 -76916 -80959
rect -76824 -81003 -76816 -80959
rect -76724 -81003 -76716 -80959
rect -76624 -81003 -76616 -80959
rect -76524 -81003 -76516 -80959
rect -76424 -81003 -76416 -80959
rect -76324 -81003 -76316 -80959
rect -76224 -81003 -76216 -80959
rect -76124 -81003 -76116 -80959
rect -76024 -81003 -76016 -80959
rect -75924 -81003 -75916 -80959
rect -75824 -81003 -75816 -80959
rect -75724 -81003 -75716 -80959
rect -75624 -81003 -75616 -80959
rect -75524 -81003 -75516 -80959
rect -75424 -81003 -75416 -80959
rect -50017 -80961 -49973 -80953
rect -49917 -80961 -49873 -80953
rect -49817 -80961 -49773 -80953
rect -49717 -80961 -49673 -80953
rect -49617 -80961 -49573 -80953
rect -49517 -80961 -49473 -80953
rect -49417 -80961 -49373 -80953
rect -49317 -80961 -49273 -80953
rect -49217 -80961 -49173 -80953
rect -49117 -80961 -49073 -80953
rect -49017 -80961 -48973 -80953
rect -48917 -80961 -48873 -80953
rect -48817 -80961 -48773 -80953
rect -48717 -80961 -48673 -80953
rect -48617 -80961 -48573 -80953
rect -48517 -80961 -48473 -80953
rect -48017 -80961 -47973 -80953
rect -47917 -80961 -47873 -80953
rect -47817 -80961 -47773 -80953
rect -47717 -80961 -47673 -80953
rect -47617 -80961 -47573 -80953
rect -47517 -80961 -47473 -80953
rect -47417 -80961 -47373 -80953
rect -47317 -80961 -47273 -80953
rect -47217 -80961 -47173 -80953
rect -47117 -80961 -47073 -80953
rect -47017 -80961 -46973 -80953
rect -46917 -80961 -46873 -80953
rect -46817 -80961 -46773 -80953
rect -46717 -80961 -46673 -80953
rect -46617 -80961 -46573 -80953
rect -46517 -80961 -46473 -80953
rect -46017 -80961 -45973 -80953
rect -45917 -80961 -45873 -80953
rect -45817 -80961 -45773 -80953
rect -45717 -80961 -45673 -80953
rect -45617 -80961 -45573 -80953
rect -45517 -80961 -45473 -80953
rect -45417 -80961 -45373 -80953
rect -45317 -80961 -45273 -80953
rect -45217 -80961 -45173 -80953
rect -45117 -80961 -45073 -80953
rect -45017 -80961 -44973 -80953
rect -44917 -80961 -44873 -80953
rect -44817 -80961 -44773 -80953
rect -44717 -80961 -44673 -80953
rect -44617 -80961 -44573 -80953
rect -44517 -80961 -44473 -80953
rect -44017 -80961 -43973 -80953
rect -43917 -80961 -43873 -80953
rect -43817 -80961 -43773 -80953
rect -43717 -80961 -43673 -80953
rect -43617 -80961 -43573 -80953
rect -43517 -80961 -43473 -80953
rect -43417 -80961 -43373 -80953
rect -43317 -80961 -43273 -80953
rect -43217 -80961 -43173 -80953
rect -43117 -80961 -43073 -80953
rect -43017 -80961 -42973 -80953
rect -42917 -80961 -42873 -80953
rect -42817 -80961 -42773 -80953
rect -42717 -80961 -42673 -80953
rect -42617 -80961 -42573 -80953
rect -42517 -80961 -42473 -80953
rect 80737 -80955 80781 -80947
rect 80837 -80955 80881 -80947
rect 80937 -80955 80981 -80947
rect 81037 -80955 81081 -80947
rect 81137 -80955 81181 -80947
rect 81237 -80955 81281 -80947
rect 81337 -80955 81381 -80947
rect 81437 -80955 81481 -80947
rect 81537 -80955 81581 -80947
rect 81637 -80955 81681 -80947
rect 81737 -80955 81781 -80947
rect 81837 -80955 81881 -80947
rect 81937 -80955 81981 -80947
rect 82037 -80955 82081 -80947
rect 82137 -80955 82181 -80947
rect 82237 -80955 82281 -80947
rect 82737 -80955 82781 -80947
rect 82837 -80955 82881 -80947
rect 82937 -80955 82981 -80947
rect 83037 -80955 83081 -80947
rect 83137 -80955 83181 -80947
rect 83237 -80955 83281 -80947
rect 83337 -80955 83381 -80947
rect 83437 -80955 83481 -80947
rect 83537 -80955 83581 -80947
rect 83637 -80955 83681 -80947
rect 83737 -80955 83781 -80947
rect 83837 -80955 83881 -80947
rect 83937 -80955 83981 -80947
rect 84037 -80955 84081 -80947
rect 84137 -80955 84181 -80947
rect 84237 -80955 84281 -80947
rect 84737 -80955 84781 -80947
rect 84837 -80955 84881 -80947
rect 84937 -80955 84981 -80947
rect 85037 -80955 85081 -80947
rect 85137 -80955 85181 -80947
rect 85237 -80955 85281 -80947
rect 85337 -80955 85381 -80947
rect 85437 -80955 85481 -80947
rect 85537 -80955 85581 -80947
rect 85637 -80955 85681 -80947
rect 85737 -80955 85781 -80947
rect 85837 -80955 85881 -80947
rect 85937 -80955 85981 -80947
rect 86037 -80955 86081 -80947
rect 86137 -80955 86181 -80947
rect 86237 -80955 86281 -80947
rect 86737 -80955 86781 -80947
rect 86837 -80955 86881 -80947
rect 86937 -80955 86981 -80947
rect 87037 -80955 87081 -80947
rect 87137 -80955 87181 -80947
rect 87237 -80955 87281 -80947
rect 87337 -80955 87381 -80947
rect 87437 -80955 87481 -80947
rect 87537 -80955 87581 -80947
rect 87637 -80955 87681 -80947
rect 87737 -80955 87781 -80947
rect 87837 -80955 87881 -80947
rect 87937 -80955 87981 -80947
rect 88037 -80955 88081 -80947
rect 88137 -80955 88181 -80947
rect 88237 -80955 88281 -80947
rect -49973 -81005 -49965 -80961
rect -49873 -81005 -49865 -80961
rect -49773 -81005 -49765 -80961
rect -49673 -81005 -49665 -80961
rect -49573 -81005 -49565 -80961
rect -49473 -81005 -49465 -80961
rect -49373 -81005 -49365 -80961
rect -49273 -81005 -49265 -80961
rect -49173 -81005 -49165 -80961
rect -49073 -81005 -49065 -80961
rect -48973 -81005 -48965 -80961
rect -48873 -81005 -48865 -80961
rect -48773 -81005 -48765 -80961
rect -48673 -81005 -48665 -80961
rect -48573 -81005 -48565 -80961
rect -48473 -81005 -48465 -80961
rect -47973 -81005 -47965 -80961
rect -47873 -81005 -47865 -80961
rect -47773 -81005 -47765 -80961
rect -47673 -81005 -47665 -80961
rect -47573 -81005 -47565 -80961
rect -47473 -81005 -47465 -80961
rect -47373 -81005 -47365 -80961
rect -47273 -81005 -47265 -80961
rect -47173 -81005 -47165 -80961
rect -47073 -81005 -47065 -80961
rect -46973 -81005 -46965 -80961
rect -46873 -81005 -46865 -80961
rect -46773 -81005 -46765 -80961
rect -46673 -81005 -46665 -80961
rect -46573 -81005 -46565 -80961
rect -46473 -81005 -46465 -80961
rect -45973 -81005 -45965 -80961
rect -45873 -81005 -45865 -80961
rect -45773 -81005 -45765 -80961
rect -45673 -81005 -45665 -80961
rect -45573 -81005 -45565 -80961
rect -45473 -81005 -45465 -80961
rect -45373 -81005 -45365 -80961
rect -45273 -81005 -45265 -80961
rect -45173 -81005 -45165 -80961
rect -45073 -81005 -45065 -80961
rect -44973 -81005 -44965 -80961
rect -44873 -81005 -44865 -80961
rect -44773 -81005 -44765 -80961
rect -44673 -81005 -44665 -80961
rect -44573 -81005 -44565 -80961
rect -44473 -81005 -44465 -80961
rect -43973 -81005 -43965 -80961
rect -43873 -81005 -43865 -80961
rect -43773 -81005 -43765 -80961
rect -43673 -81005 -43665 -80961
rect -43573 -81005 -43565 -80961
rect -43473 -81005 -43465 -80961
rect -43373 -81005 -43365 -80961
rect -43273 -81005 -43265 -80961
rect -43173 -81005 -43165 -80961
rect -43073 -81005 -43065 -80961
rect -42973 -81005 -42965 -80961
rect -42873 -81005 -42865 -80961
rect -42773 -81005 -42765 -80961
rect -42673 -81005 -42665 -80961
rect -42573 -81005 -42565 -80961
rect -42473 -81005 -42465 -80961
rect 80781 -80999 80789 -80955
rect 80881 -80999 80889 -80955
rect 80981 -80999 80989 -80955
rect 81081 -80999 81089 -80955
rect 81181 -80999 81189 -80955
rect 81281 -80999 81289 -80955
rect 81381 -80999 81389 -80955
rect 81481 -80999 81489 -80955
rect 81581 -80999 81589 -80955
rect 81681 -80999 81689 -80955
rect 81781 -80999 81789 -80955
rect 81881 -80999 81889 -80955
rect 81981 -80999 81989 -80955
rect 82081 -80999 82089 -80955
rect 82181 -80999 82189 -80955
rect 82281 -80999 82289 -80955
rect 82781 -80999 82789 -80955
rect 82881 -80999 82889 -80955
rect 82981 -80999 82989 -80955
rect 83081 -80999 83089 -80955
rect 83181 -80999 83189 -80955
rect 83281 -80999 83289 -80955
rect 83381 -80999 83389 -80955
rect 83481 -80999 83489 -80955
rect 83581 -80999 83589 -80955
rect 83681 -80999 83689 -80955
rect 83781 -80999 83789 -80955
rect 83881 -80999 83889 -80955
rect 83981 -80999 83989 -80955
rect 84081 -80999 84089 -80955
rect 84181 -80999 84189 -80955
rect 84281 -80999 84289 -80955
rect 84781 -80999 84789 -80955
rect 84881 -80999 84889 -80955
rect 84981 -80999 84989 -80955
rect 85081 -80999 85089 -80955
rect 85181 -80999 85189 -80955
rect 85281 -80999 85289 -80955
rect 85381 -80999 85389 -80955
rect 85481 -80999 85489 -80955
rect 85581 -80999 85589 -80955
rect 85681 -80999 85689 -80955
rect 85781 -80999 85789 -80955
rect 85881 -80999 85889 -80955
rect 85981 -80999 85989 -80955
rect 86081 -80999 86089 -80955
rect 86181 -80999 86189 -80955
rect 86281 -80999 86289 -80955
rect 86781 -80999 86789 -80955
rect 86881 -80999 86889 -80955
rect 86981 -80999 86989 -80955
rect 87081 -80999 87089 -80955
rect 87181 -80999 87189 -80955
rect 87281 -80999 87289 -80955
rect 87381 -80999 87389 -80955
rect 87481 -80999 87489 -80955
rect 87581 -80999 87589 -80955
rect 87681 -80999 87689 -80955
rect 87781 -80999 87789 -80955
rect 87881 -80999 87889 -80955
rect 87981 -80999 87989 -80955
rect 88081 -80999 88089 -80955
rect 88181 -80999 88189 -80955
rect 88281 -80999 88289 -80955
rect -82968 -81059 -82924 -81051
rect -82868 -81059 -82824 -81051
rect -82768 -81059 -82724 -81051
rect -82668 -81059 -82624 -81051
rect -82568 -81059 -82524 -81051
rect -82468 -81059 -82424 -81051
rect -82368 -81059 -82324 -81051
rect -82268 -81059 -82224 -81051
rect -82168 -81059 -82124 -81051
rect -82068 -81059 -82024 -81051
rect -81968 -81059 -81924 -81051
rect -81868 -81059 -81824 -81051
rect -81768 -81059 -81724 -81051
rect -81668 -81059 -81624 -81051
rect -81568 -81059 -81524 -81051
rect -81468 -81059 -81424 -81051
rect -80968 -81059 -80924 -81051
rect -80868 -81059 -80824 -81051
rect -80768 -81059 -80724 -81051
rect -80668 -81059 -80624 -81051
rect -80568 -81059 -80524 -81051
rect -80468 -81059 -80424 -81051
rect -80368 -81059 -80324 -81051
rect -80268 -81059 -80224 -81051
rect -80168 -81059 -80124 -81051
rect -80068 -81059 -80024 -81051
rect -79968 -81059 -79924 -81051
rect -79868 -81059 -79824 -81051
rect -79768 -81059 -79724 -81051
rect -79668 -81059 -79624 -81051
rect -79568 -81059 -79524 -81051
rect -79468 -81059 -79424 -81051
rect -78968 -81059 -78924 -81051
rect -78868 -81059 -78824 -81051
rect -78768 -81059 -78724 -81051
rect -78668 -81059 -78624 -81051
rect -78568 -81059 -78524 -81051
rect -78468 -81059 -78424 -81051
rect -78368 -81059 -78324 -81051
rect -78268 -81059 -78224 -81051
rect -78168 -81059 -78124 -81051
rect -78068 -81059 -78024 -81051
rect -77968 -81059 -77924 -81051
rect -77868 -81059 -77824 -81051
rect -77768 -81059 -77724 -81051
rect -77668 -81059 -77624 -81051
rect -77568 -81059 -77524 -81051
rect -77468 -81059 -77424 -81051
rect -76968 -81059 -76924 -81051
rect -76868 -81059 -76824 -81051
rect -76768 -81059 -76724 -81051
rect -76668 -81059 -76624 -81051
rect -76568 -81059 -76524 -81051
rect -76468 -81059 -76424 -81051
rect -76368 -81059 -76324 -81051
rect -76268 -81059 -76224 -81051
rect -76168 -81059 -76124 -81051
rect -76068 -81059 -76024 -81051
rect -75968 -81059 -75924 -81051
rect -75868 -81059 -75824 -81051
rect -75768 -81059 -75724 -81051
rect -75668 -81059 -75624 -81051
rect -75568 -81059 -75524 -81051
rect -75468 -81059 -75424 -81051
rect -82924 -81103 -82916 -81059
rect -82824 -81103 -82816 -81059
rect -82724 -81103 -82716 -81059
rect -82624 -81103 -82616 -81059
rect -82524 -81103 -82516 -81059
rect -82424 -81103 -82416 -81059
rect -82324 -81103 -82316 -81059
rect -82224 -81103 -82216 -81059
rect -82124 -81103 -82116 -81059
rect -82024 -81103 -82016 -81059
rect -81924 -81103 -81916 -81059
rect -81824 -81103 -81816 -81059
rect -81724 -81103 -81716 -81059
rect -81624 -81103 -81616 -81059
rect -81524 -81103 -81516 -81059
rect -81424 -81103 -81416 -81059
rect -80924 -81103 -80916 -81059
rect -80824 -81103 -80816 -81059
rect -80724 -81103 -80716 -81059
rect -80624 -81103 -80616 -81059
rect -80524 -81103 -80516 -81059
rect -80424 -81103 -80416 -81059
rect -80324 -81103 -80316 -81059
rect -80224 -81103 -80216 -81059
rect -80124 -81103 -80116 -81059
rect -80024 -81103 -80016 -81059
rect -79924 -81103 -79916 -81059
rect -79824 -81103 -79816 -81059
rect -79724 -81103 -79716 -81059
rect -79624 -81103 -79616 -81059
rect -79524 -81103 -79516 -81059
rect -79424 -81103 -79416 -81059
rect -78924 -81103 -78916 -81059
rect -78824 -81103 -78816 -81059
rect -78724 -81103 -78716 -81059
rect -78624 -81103 -78616 -81059
rect -78524 -81103 -78516 -81059
rect -78424 -81103 -78416 -81059
rect -78324 -81103 -78316 -81059
rect -78224 -81103 -78216 -81059
rect -78124 -81103 -78116 -81059
rect -78024 -81103 -78016 -81059
rect -77924 -81103 -77916 -81059
rect -77824 -81103 -77816 -81059
rect -77724 -81103 -77716 -81059
rect -77624 -81103 -77616 -81059
rect -77524 -81103 -77516 -81059
rect -77424 -81103 -77416 -81059
rect -76924 -81103 -76916 -81059
rect -76824 -81103 -76816 -81059
rect -76724 -81103 -76716 -81059
rect -76624 -81103 -76616 -81059
rect -76524 -81103 -76516 -81059
rect -76424 -81103 -76416 -81059
rect -76324 -81103 -76316 -81059
rect -76224 -81103 -76216 -81059
rect -76124 -81103 -76116 -81059
rect -76024 -81103 -76016 -81059
rect -75924 -81103 -75916 -81059
rect -75824 -81103 -75816 -81059
rect -75724 -81103 -75716 -81059
rect -75624 -81103 -75616 -81059
rect -75524 -81103 -75516 -81059
rect -75424 -81103 -75416 -81059
rect -50017 -81061 -49973 -81053
rect -49917 -81061 -49873 -81053
rect -49817 -81061 -49773 -81053
rect -49717 -81061 -49673 -81053
rect -49617 -81061 -49573 -81053
rect -49517 -81061 -49473 -81053
rect -49417 -81061 -49373 -81053
rect -49317 -81061 -49273 -81053
rect -49217 -81061 -49173 -81053
rect -49117 -81061 -49073 -81053
rect -49017 -81061 -48973 -81053
rect -48917 -81061 -48873 -81053
rect -48817 -81061 -48773 -81053
rect -48717 -81061 -48673 -81053
rect -48617 -81061 -48573 -81053
rect -48517 -81061 -48473 -81053
rect -48017 -81061 -47973 -81053
rect -47917 -81061 -47873 -81053
rect -47817 -81061 -47773 -81053
rect -47717 -81061 -47673 -81053
rect -47617 -81061 -47573 -81053
rect -47517 -81061 -47473 -81053
rect -47417 -81061 -47373 -81053
rect -47317 -81061 -47273 -81053
rect -47217 -81061 -47173 -81053
rect -47117 -81061 -47073 -81053
rect -47017 -81061 -46973 -81053
rect -46917 -81061 -46873 -81053
rect -46817 -81061 -46773 -81053
rect -46717 -81061 -46673 -81053
rect -46617 -81061 -46573 -81053
rect -46517 -81061 -46473 -81053
rect -46017 -81061 -45973 -81053
rect -45917 -81061 -45873 -81053
rect -45817 -81061 -45773 -81053
rect -45717 -81061 -45673 -81053
rect -45617 -81061 -45573 -81053
rect -45517 -81061 -45473 -81053
rect -45417 -81061 -45373 -81053
rect -45317 -81061 -45273 -81053
rect -45217 -81061 -45173 -81053
rect -45117 -81061 -45073 -81053
rect -45017 -81061 -44973 -81053
rect -44917 -81061 -44873 -81053
rect -44817 -81061 -44773 -81053
rect -44717 -81061 -44673 -81053
rect -44617 -81061 -44573 -81053
rect -44517 -81061 -44473 -81053
rect -44017 -81061 -43973 -81053
rect -43917 -81061 -43873 -81053
rect -43817 -81061 -43773 -81053
rect -43717 -81061 -43673 -81053
rect -43617 -81061 -43573 -81053
rect -43517 -81061 -43473 -81053
rect -43417 -81061 -43373 -81053
rect -43317 -81061 -43273 -81053
rect -43217 -81061 -43173 -81053
rect -43117 -81061 -43073 -81053
rect -43017 -81061 -42973 -81053
rect -42917 -81061 -42873 -81053
rect -42817 -81061 -42773 -81053
rect -42717 -81061 -42673 -81053
rect -42617 -81061 -42573 -81053
rect -42517 -81061 -42473 -81053
rect 80737 -81055 80781 -81047
rect 80837 -81055 80881 -81047
rect 80937 -81055 80981 -81047
rect 81037 -81055 81081 -81047
rect 81137 -81055 81181 -81047
rect 81237 -81055 81281 -81047
rect 81337 -81055 81381 -81047
rect 81437 -81055 81481 -81047
rect 81537 -81055 81581 -81047
rect 81637 -81055 81681 -81047
rect 81737 -81055 81781 -81047
rect 81837 -81055 81881 -81047
rect 81937 -81055 81981 -81047
rect 82037 -81055 82081 -81047
rect 82137 -81055 82181 -81047
rect 82237 -81055 82281 -81047
rect 82737 -81055 82781 -81047
rect 82837 -81055 82881 -81047
rect 82937 -81055 82981 -81047
rect 83037 -81055 83081 -81047
rect 83137 -81055 83181 -81047
rect 83237 -81055 83281 -81047
rect 83337 -81055 83381 -81047
rect 83437 -81055 83481 -81047
rect 83537 -81055 83581 -81047
rect 83637 -81055 83681 -81047
rect 83737 -81055 83781 -81047
rect 83837 -81055 83881 -81047
rect 83937 -81055 83981 -81047
rect 84037 -81055 84081 -81047
rect 84137 -81055 84181 -81047
rect 84237 -81055 84281 -81047
rect 84737 -81055 84781 -81047
rect 84837 -81055 84881 -81047
rect 84937 -81055 84981 -81047
rect 85037 -81055 85081 -81047
rect 85137 -81055 85181 -81047
rect 85237 -81055 85281 -81047
rect 85337 -81055 85381 -81047
rect 85437 -81055 85481 -81047
rect 85537 -81055 85581 -81047
rect 85637 -81055 85681 -81047
rect 85737 -81055 85781 -81047
rect 85837 -81055 85881 -81047
rect 85937 -81055 85981 -81047
rect 86037 -81055 86081 -81047
rect 86137 -81055 86181 -81047
rect 86237 -81055 86281 -81047
rect 86737 -81055 86781 -81047
rect 86837 -81055 86881 -81047
rect 86937 -81055 86981 -81047
rect 87037 -81055 87081 -81047
rect 87137 -81055 87181 -81047
rect 87237 -81055 87281 -81047
rect 87337 -81055 87381 -81047
rect 87437 -81055 87481 -81047
rect 87537 -81055 87581 -81047
rect 87637 -81055 87681 -81047
rect 87737 -81055 87781 -81047
rect 87837 -81055 87881 -81047
rect 87937 -81055 87981 -81047
rect 88037 -81055 88081 -81047
rect 88137 -81055 88181 -81047
rect 88237 -81055 88281 -81047
rect -49973 -81105 -49965 -81061
rect -49873 -81105 -49865 -81061
rect -49773 -81105 -49765 -81061
rect -49673 -81105 -49665 -81061
rect -49573 -81105 -49565 -81061
rect -49473 -81105 -49465 -81061
rect -49373 -81105 -49365 -81061
rect -49273 -81105 -49265 -81061
rect -49173 -81105 -49165 -81061
rect -49073 -81105 -49065 -81061
rect -48973 -81105 -48965 -81061
rect -48873 -81105 -48865 -81061
rect -48773 -81105 -48765 -81061
rect -48673 -81105 -48665 -81061
rect -48573 -81105 -48565 -81061
rect -48473 -81105 -48465 -81061
rect -47973 -81105 -47965 -81061
rect -47873 -81105 -47865 -81061
rect -47773 -81105 -47765 -81061
rect -47673 -81105 -47665 -81061
rect -47573 -81105 -47565 -81061
rect -47473 -81105 -47465 -81061
rect -47373 -81105 -47365 -81061
rect -47273 -81105 -47265 -81061
rect -47173 -81105 -47165 -81061
rect -47073 -81105 -47065 -81061
rect -46973 -81105 -46965 -81061
rect -46873 -81105 -46865 -81061
rect -46773 -81105 -46765 -81061
rect -46673 -81105 -46665 -81061
rect -46573 -81105 -46565 -81061
rect -46473 -81105 -46465 -81061
rect -45973 -81105 -45965 -81061
rect -45873 -81105 -45865 -81061
rect -45773 -81105 -45765 -81061
rect -45673 -81105 -45665 -81061
rect -45573 -81105 -45565 -81061
rect -45473 -81105 -45465 -81061
rect -45373 -81105 -45365 -81061
rect -45273 -81105 -45265 -81061
rect -45173 -81105 -45165 -81061
rect -45073 -81105 -45065 -81061
rect -44973 -81105 -44965 -81061
rect -44873 -81105 -44865 -81061
rect -44773 -81105 -44765 -81061
rect -44673 -81105 -44665 -81061
rect -44573 -81105 -44565 -81061
rect -44473 -81105 -44465 -81061
rect -43973 -81105 -43965 -81061
rect -43873 -81105 -43865 -81061
rect -43773 -81105 -43765 -81061
rect -43673 -81105 -43665 -81061
rect -43573 -81105 -43565 -81061
rect -43473 -81105 -43465 -81061
rect -43373 -81105 -43365 -81061
rect -43273 -81105 -43265 -81061
rect -43173 -81105 -43165 -81061
rect -43073 -81105 -43065 -81061
rect -42973 -81105 -42965 -81061
rect -42873 -81105 -42865 -81061
rect -42773 -81105 -42765 -81061
rect -42673 -81105 -42665 -81061
rect -42573 -81105 -42565 -81061
rect -42473 -81105 -42465 -81061
rect 80781 -81099 80789 -81055
rect 80881 -81099 80889 -81055
rect 80981 -81099 80989 -81055
rect 81081 -81099 81089 -81055
rect 81181 -81099 81189 -81055
rect 81281 -81099 81289 -81055
rect 81381 -81099 81389 -81055
rect 81481 -81099 81489 -81055
rect 81581 -81099 81589 -81055
rect 81681 -81099 81689 -81055
rect 81781 -81099 81789 -81055
rect 81881 -81099 81889 -81055
rect 81981 -81099 81989 -81055
rect 82081 -81099 82089 -81055
rect 82181 -81099 82189 -81055
rect 82281 -81099 82289 -81055
rect 82781 -81099 82789 -81055
rect 82881 -81099 82889 -81055
rect 82981 -81099 82989 -81055
rect 83081 -81099 83089 -81055
rect 83181 -81099 83189 -81055
rect 83281 -81099 83289 -81055
rect 83381 -81099 83389 -81055
rect 83481 -81099 83489 -81055
rect 83581 -81099 83589 -81055
rect 83681 -81099 83689 -81055
rect 83781 -81099 83789 -81055
rect 83881 -81099 83889 -81055
rect 83981 -81099 83989 -81055
rect 84081 -81099 84089 -81055
rect 84181 -81099 84189 -81055
rect 84281 -81099 84289 -81055
rect 84781 -81099 84789 -81055
rect 84881 -81099 84889 -81055
rect 84981 -81099 84989 -81055
rect 85081 -81099 85089 -81055
rect 85181 -81099 85189 -81055
rect 85281 -81099 85289 -81055
rect 85381 -81099 85389 -81055
rect 85481 -81099 85489 -81055
rect 85581 -81099 85589 -81055
rect 85681 -81099 85689 -81055
rect 85781 -81099 85789 -81055
rect 85881 -81099 85889 -81055
rect 85981 -81099 85989 -81055
rect 86081 -81099 86089 -81055
rect 86181 -81099 86189 -81055
rect 86281 -81099 86289 -81055
rect 86781 -81099 86789 -81055
rect 86881 -81099 86889 -81055
rect 86981 -81099 86989 -81055
rect 87081 -81099 87089 -81055
rect 87181 -81099 87189 -81055
rect 87281 -81099 87289 -81055
rect 87381 -81099 87389 -81055
rect 87481 -81099 87489 -81055
rect 87581 -81099 87589 -81055
rect 87681 -81099 87689 -81055
rect 87781 -81099 87789 -81055
rect 87881 -81099 87889 -81055
rect 87981 -81099 87989 -81055
rect 88081 -81099 88089 -81055
rect 88181 -81099 88189 -81055
rect 88281 -81099 88289 -81055
rect -82968 -81159 -82924 -81151
rect -82868 -81159 -82824 -81151
rect -82768 -81159 -82724 -81151
rect -82668 -81159 -82624 -81151
rect -82568 -81159 -82524 -81151
rect -82468 -81159 -82424 -81151
rect -82368 -81159 -82324 -81151
rect -82268 -81159 -82224 -81151
rect -82168 -81159 -82124 -81151
rect -82068 -81159 -82024 -81151
rect -81968 -81159 -81924 -81151
rect -81868 -81159 -81824 -81151
rect -81768 -81159 -81724 -81151
rect -81668 -81159 -81624 -81151
rect -81568 -81159 -81524 -81151
rect -81468 -81159 -81424 -81151
rect -80968 -81159 -80924 -81151
rect -80868 -81159 -80824 -81151
rect -80768 -81159 -80724 -81151
rect -80668 -81159 -80624 -81151
rect -80568 -81159 -80524 -81151
rect -80468 -81159 -80424 -81151
rect -80368 -81159 -80324 -81151
rect -80268 -81159 -80224 -81151
rect -80168 -81159 -80124 -81151
rect -80068 -81159 -80024 -81151
rect -79968 -81159 -79924 -81151
rect -79868 -81159 -79824 -81151
rect -79768 -81159 -79724 -81151
rect -79668 -81159 -79624 -81151
rect -79568 -81159 -79524 -81151
rect -79468 -81159 -79424 -81151
rect -78968 -81159 -78924 -81151
rect -78868 -81159 -78824 -81151
rect -78768 -81159 -78724 -81151
rect -78668 -81159 -78624 -81151
rect -78568 -81159 -78524 -81151
rect -78468 -81159 -78424 -81151
rect -78368 -81159 -78324 -81151
rect -78268 -81159 -78224 -81151
rect -78168 -81159 -78124 -81151
rect -78068 -81159 -78024 -81151
rect -77968 -81159 -77924 -81151
rect -77868 -81159 -77824 -81151
rect -77768 -81159 -77724 -81151
rect -77668 -81159 -77624 -81151
rect -77568 -81159 -77524 -81151
rect -77468 -81159 -77424 -81151
rect -76968 -81159 -76924 -81151
rect -76868 -81159 -76824 -81151
rect -76768 -81159 -76724 -81151
rect -76668 -81159 -76624 -81151
rect -76568 -81159 -76524 -81151
rect -76468 -81159 -76424 -81151
rect -76368 -81159 -76324 -81151
rect -76268 -81159 -76224 -81151
rect -76168 -81159 -76124 -81151
rect -76068 -81159 -76024 -81151
rect -75968 -81159 -75924 -81151
rect -75868 -81159 -75824 -81151
rect -75768 -81159 -75724 -81151
rect -75668 -81159 -75624 -81151
rect -75568 -81159 -75524 -81151
rect -75468 -81159 -75424 -81151
rect -82924 -81203 -82916 -81159
rect -82824 -81203 -82816 -81159
rect -82724 -81203 -82716 -81159
rect -82624 -81203 -82616 -81159
rect -82524 -81203 -82516 -81159
rect -82424 -81203 -82416 -81159
rect -82324 -81203 -82316 -81159
rect -82224 -81203 -82216 -81159
rect -82124 -81203 -82116 -81159
rect -82024 -81203 -82016 -81159
rect -81924 -81203 -81916 -81159
rect -81824 -81203 -81816 -81159
rect -81724 -81203 -81716 -81159
rect -81624 -81203 -81616 -81159
rect -81524 -81203 -81516 -81159
rect -81424 -81203 -81416 -81159
rect -80924 -81203 -80916 -81159
rect -80824 -81203 -80816 -81159
rect -80724 -81203 -80716 -81159
rect -80624 -81203 -80616 -81159
rect -80524 -81203 -80516 -81159
rect -80424 -81203 -80416 -81159
rect -80324 -81203 -80316 -81159
rect -80224 -81203 -80216 -81159
rect -80124 -81203 -80116 -81159
rect -80024 -81203 -80016 -81159
rect -79924 -81203 -79916 -81159
rect -79824 -81203 -79816 -81159
rect -79724 -81203 -79716 -81159
rect -79624 -81203 -79616 -81159
rect -79524 -81203 -79516 -81159
rect -79424 -81203 -79416 -81159
rect -78924 -81203 -78916 -81159
rect -78824 -81203 -78816 -81159
rect -78724 -81203 -78716 -81159
rect -78624 -81203 -78616 -81159
rect -78524 -81203 -78516 -81159
rect -78424 -81203 -78416 -81159
rect -78324 -81203 -78316 -81159
rect -78224 -81203 -78216 -81159
rect -78124 -81203 -78116 -81159
rect -78024 -81203 -78016 -81159
rect -77924 -81203 -77916 -81159
rect -77824 -81203 -77816 -81159
rect -77724 -81203 -77716 -81159
rect -77624 -81203 -77616 -81159
rect -77524 -81203 -77516 -81159
rect -77424 -81203 -77416 -81159
rect -76924 -81203 -76916 -81159
rect -76824 -81203 -76816 -81159
rect -76724 -81203 -76716 -81159
rect -76624 -81203 -76616 -81159
rect -76524 -81203 -76516 -81159
rect -76424 -81203 -76416 -81159
rect -76324 -81203 -76316 -81159
rect -76224 -81203 -76216 -81159
rect -76124 -81203 -76116 -81159
rect -76024 -81203 -76016 -81159
rect -75924 -81203 -75916 -81159
rect -75824 -81203 -75816 -81159
rect -75724 -81203 -75716 -81159
rect -75624 -81203 -75616 -81159
rect -75524 -81203 -75516 -81159
rect -75424 -81203 -75416 -81159
rect -50017 -81161 -49973 -81153
rect -49917 -81161 -49873 -81153
rect -49817 -81161 -49773 -81153
rect -49717 -81161 -49673 -81153
rect -49617 -81161 -49573 -81153
rect -49517 -81161 -49473 -81153
rect -49417 -81161 -49373 -81153
rect -49317 -81161 -49273 -81153
rect -49217 -81161 -49173 -81153
rect -49117 -81161 -49073 -81153
rect -49017 -81161 -48973 -81153
rect -48917 -81161 -48873 -81153
rect -48817 -81161 -48773 -81153
rect -48717 -81161 -48673 -81153
rect -48617 -81161 -48573 -81153
rect -48517 -81161 -48473 -81153
rect -48017 -81161 -47973 -81153
rect -47917 -81161 -47873 -81153
rect -47817 -81161 -47773 -81153
rect -47717 -81161 -47673 -81153
rect -47617 -81161 -47573 -81153
rect -47517 -81161 -47473 -81153
rect -47417 -81161 -47373 -81153
rect -47317 -81161 -47273 -81153
rect -47217 -81161 -47173 -81153
rect -47117 -81161 -47073 -81153
rect -47017 -81161 -46973 -81153
rect -46917 -81161 -46873 -81153
rect -46817 -81161 -46773 -81153
rect -46717 -81161 -46673 -81153
rect -46617 -81161 -46573 -81153
rect -46517 -81161 -46473 -81153
rect -46017 -81161 -45973 -81153
rect -45917 -81161 -45873 -81153
rect -45817 -81161 -45773 -81153
rect -45717 -81161 -45673 -81153
rect -45617 -81161 -45573 -81153
rect -45517 -81161 -45473 -81153
rect -45417 -81161 -45373 -81153
rect -45317 -81161 -45273 -81153
rect -45217 -81161 -45173 -81153
rect -45117 -81161 -45073 -81153
rect -45017 -81161 -44973 -81153
rect -44917 -81161 -44873 -81153
rect -44817 -81161 -44773 -81153
rect -44717 -81161 -44673 -81153
rect -44617 -81161 -44573 -81153
rect -44517 -81161 -44473 -81153
rect -44017 -81161 -43973 -81153
rect -43917 -81161 -43873 -81153
rect -43817 -81161 -43773 -81153
rect -43717 -81161 -43673 -81153
rect -43617 -81161 -43573 -81153
rect -43517 -81161 -43473 -81153
rect -43417 -81161 -43373 -81153
rect -43317 -81161 -43273 -81153
rect -43217 -81161 -43173 -81153
rect -43117 -81161 -43073 -81153
rect -43017 -81161 -42973 -81153
rect -42917 -81161 -42873 -81153
rect -42817 -81161 -42773 -81153
rect -42717 -81161 -42673 -81153
rect -42617 -81161 -42573 -81153
rect -42517 -81161 -42473 -81153
rect 80737 -81155 80781 -81147
rect 80837 -81155 80881 -81147
rect 80937 -81155 80981 -81147
rect 81037 -81155 81081 -81147
rect 81137 -81155 81181 -81147
rect 81237 -81155 81281 -81147
rect 81337 -81155 81381 -81147
rect 81437 -81155 81481 -81147
rect 81537 -81155 81581 -81147
rect 81637 -81155 81681 -81147
rect 81737 -81155 81781 -81147
rect 81837 -81155 81881 -81147
rect 81937 -81155 81981 -81147
rect 82037 -81155 82081 -81147
rect 82137 -81155 82181 -81147
rect 82237 -81155 82281 -81147
rect 82737 -81155 82781 -81147
rect 82837 -81155 82881 -81147
rect 82937 -81155 82981 -81147
rect 83037 -81155 83081 -81147
rect 83137 -81155 83181 -81147
rect 83237 -81155 83281 -81147
rect 83337 -81155 83381 -81147
rect 83437 -81155 83481 -81147
rect 83537 -81155 83581 -81147
rect 83637 -81155 83681 -81147
rect 83737 -81155 83781 -81147
rect 83837 -81155 83881 -81147
rect 83937 -81155 83981 -81147
rect 84037 -81155 84081 -81147
rect 84137 -81155 84181 -81147
rect 84237 -81155 84281 -81147
rect 84737 -81155 84781 -81147
rect 84837 -81155 84881 -81147
rect 84937 -81155 84981 -81147
rect 85037 -81155 85081 -81147
rect 85137 -81155 85181 -81147
rect 85237 -81155 85281 -81147
rect 85337 -81155 85381 -81147
rect 85437 -81155 85481 -81147
rect 85537 -81155 85581 -81147
rect 85637 -81155 85681 -81147
rect 85737 -81155 85781 -81147
rect 85837 -81155 85881 -81147
rect 85937 -81155 85981 -81147
rect 86037 -81155 86081 -81147
rect 86137 -81155 86181 -81147
rect 86237 -81155 86281 -81147
rect 86737 -81155 86781 -81147
rect 86837 -81155 86881 -81147
rect 86937 -81155 86981 -81147
rect 87037 -81155 87081 -81147
rect 87137 -81155 87181 -81147
rect 87237 -81155 87281 -81147
rect 87337 -81155 87381 -81147
rect 87437 -81155 87481 -81147
rect 87537 -81155 87581 -81147
rect 87637 -81155 87681 -81147
rect 87737 -81155 87781 -81147
rect 87837 -81155 87881 -81147
rect 87937 -81155 87981 -81147
rect 88037 -81155 88081 -81147
rect 88137 -81155 88181 -81147
rect 88237 -81155 88281 -81147
rect -49973 -81205 -49965 -81161
rect -49873 -81205 -49865 -81161
rect -49773 -81205 -49765 -81161
rect -49673 -81205 -49665 -81161
rect -49573 -81205 -49565 -81161
rect -49473 -81205 -49465 -81161
rect -49373 -81205 -49365 -81161
rect -49273 -81205 -49265 -81161
rect -49173 -81205 -49165 -81161
rect -49073 -81205 -49065 -81161
rect -48973 -81205 -48965 -81161
rect -48873 -81205 -48865 -81161
rect -48773 -81205 -48765 -81161
rect -48673 -81205 -48665 -81161
rect -48573 -81205 -48565 -81161
rect -48473 -81205 -48465 -81161
rect -47973 -81205 -47965 -81161
rect -47873 -81205 -47865 -81161
rect -47773 -81205 -47765 -81161
rect -47673 -81205 -47665 -81161
rect -47573 -81205 -47565 -81161
rect -47473 -81205 -47465 -81161
rect -47373 -81205 -47365 -81161
rect -47273 -81205 -47265 -81161
rect -47173 -81205 -47165 -81161
rect -47073 -81205 -47065 -81161
rect -46973 -81205 -46965 -81161
rect -46873 -81205 -46865 -81161
rect -46773 -81205 -46765 -81161
rect -46673 -81205 -46665 -81161
rect -46573 -81205 -46565 -81161
rect -46473 -81205 -46465 -81161
rect -45973 -81205 -45965 -81161
rect -45873 -81205 -45865 -81161
rect -45773 -81205 -45765 -81161
rect -45673 -81205 -45665 -81161
rect -45573 -81205 -45565 -81161
rect -45473 -81205 -45465 -81161
rect -45373 -81205 -45365 -81161
rect -45273 -81205 -45265 -81161
rect -45173 -81205 -45165 -81161
rect -45073 -81205 -45065 -81161
rect -44973 -81205 -44965 -81161
rect -44873 -81205 -44865 -81161
rect -44773 -81205 -44765 -81161
rect -44673 -81205 -44665 -81161
rect -44573 -81205 -44565 -81161
rect -44473 -81205 -44465 -81161
rect -43973 -81205 -43965 -81161
rect -43873 -81205 -43865 -81161
rect -43773 -81205 -43765 -81161
rect -43673 -81205 -43665 -81161
rect -43573 -81205 -43565 -81161
rect -43473 -81205 -43465 -81161
rect -43373 -81205 -43365 -81161
rect -43273 -81205 -43265 -81161
rect -43173 -81205 -43165 -81161
rect -43073 -81205 -43065 -81161
rect -42973 -81205 -42965 -81161
rect -42873 -81205 -42865 -81161
rect -42773 -81205 -42765 -81161
rect -42673 -81205 -42665 -81161
rect -42573 -81205 -42565 -81161
rect -42473 -81205 -42465 -81161
rect 80781 -81199 80789 -81155
rect 80881 -81199 80889 -81155
rect 80981 -81199 80989 -81155
rect 81081 -81199 81089 -81155
rect 81181 -81199 81189 -81155
rect 81281 -81199 81289 -81155
rect 81381 -81199 81389 -81155
rect 81481 -81199 81489 -81155
rect 81581 -81199 81589 -81155
rect 81681 -81199 81689 -81155
rect 81781 -81199 81789 -81155
rect 81881 -81199 81889 -81155
rect 81981 -81199 81989 -81155
rect 82081 -81199 82089 -81155
rect 82181 -81199 82189 -81155
rect 82281 -81199 82289 -81155
rect 82781 -81199 82789 -81155
rect 82881 -81199 82889 -81155
rect 82981 -81199 82989 -81155
rect 83081 -81199 83089 -81155
rect 83181 -81199 83189 -81155
rect 83281 -81199 83289 -81155
rect 83381 -81199 83389 -81155
rect 83481 -81199 83489 -81155
rect 83581 -81199 83589 -81155
rect 83681 -81199 83689 -81155
rect 83781 -81199 83789 -81155
rect 83881 -81199 83889 -81155
rect 83981 -81199 83989 -81155
rect 84081 -81199 84089 -81155
rect 84181 -81199 84189 -81155
rect 84281 -81199 84289 -81155
rect 84781 -81199 84789 -81155
rect 84881 -81199 84889 -81155
rect 84981 -81199 84989 -81155
rect 85081 -81199 85089 -81155
rect 85181 -81199 85189 -81155
rect 85281 -81199 85289 -81155
rect 85381 -81199 85389 -81155
rect 85481 -81199 85489 -81155
rect 85581 -81199 85589 -81155
rect 85681 -81199 85689 -81155
rect 85781 -81199 85789 -81155
rect 85881 -81199 85889 -81155
rect 85981 -81199 85989 -81155
rect 86081 -81199 86089 -81155
rect 86181 -81199 86189 -81155
rect 86281 -81199 86289 -81155
rect 86781 -81199 86789 -81155
rect 86881 -81199 86889 -81155
rect 86981 -81199 86989 -81155
rect 87081 -81199 87089 -81155
rect 87181 -81199 87189 -81155
rect 87281 -81199 87289 -81155
rect 87381 -81199 87389 -81155
rect 87481 -81199 87489 -81155
rect 87581 -81199 87589 -81155
rect 87681 -81199 87689 -81155
rect 87781 -81199 87789 -81155
rect 87881 -81199 87889 -81155
rect 87981 -81199 87989 -81155
rect 88081 -81199 88089 -81155
rect 88181 -81199 88189 -81155
rect 88281 -81199 88289 -81155
rect -82968 -81259 -82924 -81251
rect -82868 -81259 -82824 -81251
rect -82768 -81259 -82724 -81251
rect -82668 -81259 -82624 -81251
rect -82568 -81259 -82524 -81251
rect -82468 -81259 -82424 -81251
rect -82368 -81259 -82324 -81251
rect -82268 -81259 -82224 -81251
rect -82168 -81259 -82124 -81251
rect -82068 -81259 -82024 -81251
rect -81968 -81259 -81924 -81251
rect -81868 -81259 -81824 -81251
rect -81768 -81259 -81724 -81251
rect -81668 -81259 -81624 -81251
rect -81568 -81259 -81524 -81251
rect -81468 -81259 -81424 -81251
rect -80968 -81259 -80924 -81251
rect -80868 -81259 -80824 -81251
rect -80768 -81259 -80724 -81251
rect -80668 -81259 -80624 -81251
rect -80568 -81259 -80524 -81251
rect -80468 -81259 -80424 -81251
rect -80368 -81259 -80324 -81251
rect -80268 -81259 -80224 -81251
rect -80168 -81259 -80124 -81251
rect -80068 -81259 -80024 -81251
rect -79968 -81259 -79924 -81251
rect -79868 -81259 -79824 -81251
rect -79768 -81259 -79724 -81251
rect -79668 -81259 -79624 -81251
rect -79568 -81259 -79524 -81251
rect -79468 -81259 -79424 -81251
rect -78968 -81259 -78924 -81251
rect -78868 -81259 -78824 -81251
rect -78768 -81259 -78724 -81251
rect -78668 -81259 -78624 -81251
rect -78568 -81259 -78524 -81251
rect -78468 -81259 -78424 -81251
rect -78368 -81259 -78324 -81251
rect -78268 -81259 -78224 -81251
rect -78168 -81259 -78124 -81251
rect -78068 -81259 -78024 -81251
rect -77968 -81259 -77924 -81251
rect -77868 -81259 -77824 -81251
rect -77768 -81259 -77724 -81251
rect -77668 -81259 -77624 -81251
rect -77568 -81259 -77524 -81251
rect -77468 -81259 -77424 -81251
rect -76968 -81259 -76924 -81251
rect -76868 -81259 -76824 -81251
rect -76768 -81259 -76724 -81251
rect -76668 -81259 -76624 -81251
rect -76568 -81259 -76524 -81251
rect -76468 -81259 -76424 -81251
rect -76368 -81259 -76324 -81251
rect -76268 -81259 -76224 -81251
rect -76168 -81259 -76124 -81251
rect -76068 -81259 -76024 -81251
rect -75968 -81259 -75924 -81251
rect -75868 -81259 -75824 -81251
rect -75768 -81259 -75724 -81251
rect -75668 -81259 -75624 -81251
rect -75568 -81259 -75524 -81251
rect -75468 -81259 -75424 -81251
rect -82924 -81303 -82916 -81259
rect -82824 -81303 -82816 -81259
rect -82724 -81303 -82716 -81259
rect -82624 -81303 -82616 -81259
rect -82524 -81303 -82516 -81259
rect -82424 -81303 -82416 -81259
rect -82324 -81303 -82316 -81259
rect -82224 -81303 -82216 -81259
rect -82124 -81303 -82116 -81259
rect -82024 -81303 -82016 -81259
rect -81924 -81303 -81916 -81259
rect -81824 -81303 -81816 -81259
rect -81724 -81303 -81716 -81259
rect -81624 -81303 -81616 -81259
rect -81524 -81303 -81516 -81259
rect -81424 -81303 -81416 -81259
rect -80924 -81303 -80916 -81259
rect -80824 -81303 -80816 -81259
rect -80724 -81303 -80716 -81259
rect -80624 -81303 -80616 -81259
rect -80524 -81303 -80516 -81259
rect -80424 -81303 -80416 -81259
rect -80324 -81303 -80316 -81259
rect -80224 -81303 -80216 -81259
rect -80124 -81303 -80116 -81259
rect -80024 -81303 -80016 -81259
rect -79924 -81303 -79916 -81259
rect -79824 -81303 -79816 -81259
rect -79724 -81303 -79716 -81259
rect -79624 -81303 -79616 -81259
rect -79524 -81303 -79516 -81259
rect -79424 -81303 -79416 -81259
rect -78924 -81303 -78916 -81259
rect -78824 -81303 -78816 -81259
rect -78724 -81303 -78716 -81259
rect -78624 -81303 -78616 -81259
rect -78524 -81303 -78516 -81259
rect -78424 -81303 -78416 -81259
rect -78324 -81303 -78316 -81259
rect -78224 -81303 -78216 -81259
rect -78124 -81303 -78116 -81259
rect -78024 -81303 -78016 -81259
rect -77924 -81303 -77916 -81259
rect -77824 -81303 -77816 -81259
rect -77724 -81303 -77716 -81259
rect -77624 -81303 -77616 -81259
rect -77524 -81303 -77516 -81259
rect -77424 -81303 -77416 -81259
rect -76924 -81303 -76916 -81259
rect -76824 -81303 -76816 -81259
rect -76724 -81303 -76716 -81259
rect -76624 -81303 -76616 -81259
rect -76524 -81303 -76516 -81259
rect -76424 -81303 -76416 -81259
rect -76324 -81303 -76316 -81259
rect -76224 -81303 -76216 -81259
rect -76124 -81303 -76116 -81259
rect -76024 -81303 -76016 -81259
rect -75924 -81303 -75916 -81259
rect -75824 -81303 -75816 -81259
rect -75724 -81303 -75716 -81259
rect -75624 -81303 -75616 -81259
rect -75524 -81303 -75516 -81259
rect -75424 -81303 -75416 -81259
rect -50017 -81261 -49973 -81253
rect -49917 -81261 -49873 -81253
rect -49817 -81261 -49773 -81253
rect -49717 -81261 -49673 -81253
rect -49617 -81261 -49573 -81253
rect -49517 -81261 -49473 -81253
rect -49417 -81261 -49373 -81253
rect -49317 -81261 -49273 -81253
rect -49217 -81261 -49173 -81253
rect -49117 -81261 -49073 -81253
rect -49017 -81261 -48973 -81253
rect -48917 -81261 -48873 -81253
rect -48817 -81261 -48773 -81253
rect -48717 -81261 -48673 -81253
rect -48617 -81261 -48573 -81253
rect -48517 -81261 -48473 -81253
rect -48017 -81261 -47973 -81253
rect -47917 -81261 -47873 -81253
rect -47817 -81261 -47773 -81253
rect -47717 -81261 -47673 -81253
rect -47617 -81261 -47573 -81253
rect -47517 -81261 -47473 -81253
rect -47417 -81261 -47373 -81253
rect -47317 -81261 -47273 -81253
rect -47217 -81261 -47173 -81253
rect -47117 -81261 -47073 -81253
rect -47017 -81261 -46973 -81253
rect -46917 -81261 -46873 -81253
rect -46817 -81261 -46773 -81253
rect -46717 -81261 -46673 -81253
rect -46617 -81261 -46573 -81253
rect -46517 -81261 -46473 -81253
rect -46017 -81261 -45973 -81253
rect -45917 -81261 -45873 -81253
rect -45817 -81261 -45773 -81253
rect -45717 -81261 -45673 -81253
rect -45617 -81261 -45573 -81253
rect -45517 -81261 -45473 -81253
rect -45417 -81261 -45373 -81253
rect -45317 -81261 -45273 -81253
rect -45217 -81261 -45173 -81253
rect -45117 -81261 -45073 -81253
rect -45017 -81261 -44973 -81253
rect -44917 -81261 -44873 -81253
rect -44817 -81261 -44773 -81253
rect -44717 -81261 -44673 -81253
rect -44617 -81261 -44573 -81253
rect -44517 -81261 -44473 -81253
rect -44017 -81261 -43973 -81253
rect -43917 -81261 -43873 -81253
rect -43817 -81261 -43773 -81253
rect -43717 -81261 -43673 -81253
rect -43617 -81261 -43573 -81253
rect -43517 -81261 -43473 -81253
rect -43417 -81261 -43373 -81253
rect -43317 -81261 -43273 -81253
rect -43217 -81261 -43173 -81253
rect -43117 -81261 -43073 -81253
rect -43017 -81261 -42973 -81253
rect -42917 -81261 -42873 -81253
rect -42817 -81261 -42773 -81253
rect -42717 -81261 -42673 -81253
rect -42617 -81261 -42573 -81253
rect -42517 -81261 -42473 -81253
rect 80737 -81255 80781 -81247
rect 80837 -81255 80881 -81247
rect 80937 -81255 80981 -81247
rect 81037 -81255 81081 -81247
rect 81137 -81255 81181 -81247
rect 81237 -81255 81281 -81247
rect 81337 -81255 81381 -81247
rect 81437 -81255 81481 -81247
rect 81537 -81255 81581 -81247
rect 81637 -81255 81681 -81247
rect 81737 -81255 81781 -81247
rect 81837 -81255 81881 -81247
rect 81937 -81255 81981 -81247
rect 82037 -81255 82081 -81247
rect 82137 -81255 82181 -81247
rect 82237 -81255 82281 -81247
rect 82737 -81255 82781 -81247
rect 82837 -81255 82881 -81247
rect 82937 -81255 82981 -81247
rect 83037 -81255 83081 -81247
rect 83137 -81255 83181 -81247
rect 83237 -81255 83281 -81247
rect 83337 -81255 83381 -81247
rect 83437 -81255 83481 -81247
rect 83537 -81255 83581 -81247
rect 83637 -81255 83681 -81247
rect 83737 -81255 83781 -81247
rect 83837 -81255 83881 -81247
rect 83937 -81255 83981 -81247
rect 84037 -81255 84081 -81247
rect 84137 -81255 84181 -81247
rect 84237 -81255 84281 -81247
rect 84737 -81255 84781 -81247
rect 84837 -81255 84881 -81247
rect 84937 -81255 84981 -81247
rect 85037 -81255 85081 -81247
rect 85137 -81255 85181 -81247
rect 85237 -81255 85281 -81247
rect 85337 -81255 85381 -81247
rect 85437 -81255 85481 -81247
rect 85537 -81255 85581 -81247
rect 85637 -81255 85681 -81247
rect 85737 -81255 85781 -81247
rect 85837 -81255 85881 -81247
rect 85937 -81255 85981 -81247
rect 86037 -81255 86081 -81247
rect 86137 -81255 86181 -81247
rect 86237 -81255 86281 -81247
rect 86737 -81255 86781 -81247
rect 86837 -81255 86881 -81247
rect 86937 -81255 86981 -81247
rect 87037 -81255 87081 -81247
rect 87137 -81255 87181 -81247
rect 87237 -81255 87281 -81247
rect 87337 -81255 87381 -81247
rect 87437 -81255 87481 -81247
rect 87537 -81255 87581 -81247
rect 87637 -81255 87681 -81247
rect 87737 -81255 87781 -81247
rect 87837 -81255 87881 -81247
rect 87937 -81255 87981 -81247
rect 88037 -81255 88081 -81247
rect 88137 -81255 88181 -81247
rect 88237 -81255 88281 -81247
rect -49973 -81305 -49965 -81261
rect -49873 -81305 -49865 -81261
rect -49773 -81305 -49765 -81261
rect -49673 -81305 -49665 -81261
rect -49573 -81305 -49565 -81261
rect -49473 -81305 -49465 -81261
rect -49373 -81305 -49365 -81261
rect -49273 -81305 -49265 -81261
rect -49173 -81305 -49165 -81261
rect -49073 -81305 -49065 -81261
rect -48973 -81305 -48965 -81261
rect -48873 -81305 -48865 -81261
rect -48773 -81305 -48765 -81261
rect -48673 -81305 -48665 -81261
rect -48573 -81305 -48565 -81261
rect -48473 -81305 -48465 -81261
rect -47973 -81305 -47965 -81261
rect -47873 -81305 -47865 -81261
rect -47773 -81305 -47765 -81261
rect -47673 -81305 -47665 -81261
rect -47573 -81305 -47565 -81261
rect -47473 -81305 -47465 -81261
rect -47373 -81305 -47365 -81261
rect -47273 -81305 -47265 -81261
rect -47173 -81305 -47165 -81261
rect -47073 -81305 -47065 -81261
rect -46973 -81305 -46965 -81261
rect -46873 -81305 -46865 -81261
rect -46773 -81305 -46765 -81261
rect -46673 -81305 -46665 -81261
rect -46573 -81305 -46565 -81261
rect -46473 -81305 -46465 -81261
rect -45973 -81305 -45965 -81261
rect -45873 -81305 -45865 -81261
rect -45773 -81305 -45765 -81261
rect -45673 -81305 -45665 -81261
rect -45573 -81305 -45565 -81261
rect -45473 -81305 -45465 -81261
rect -45373 -81305 -45365 -81261
rect -45273 -81305 -45265 -81261
rect -45173 -81305 -45165 -81261
rect -45073 -81305 -45065 -81261
rect -44973 -81305 -44965 -81261
rect -44873 -81305 -44865 -81261
rect -44773 -81305 -44765 -81261
rect -44673 -81305 -44665 -81261
rect -44573 -81305 -44565 -81261
rect -44473 -81305 -44465 -81261
rect -43973 -81305 -43965 -81261
rect -43873 -81305 -43865 -81261
rect -43773 -81305 -43765 -81261
rect -43673 -81305 -43665 -81261
rect -43573 -81305 -43565 -81261
rect -43473 -81305 -43465 -81261
rect -43373 -81305 -43365 -81261
rect -43273 -81305 -43265 -81261
rect -43173 -81305 -43165 -81261
rect -43073 -81305 -43065 -81261
rect -42973 -81305 -42965 -81261
rect -42873 -81305 -42865 -81261
rect -42773 -81305 -42765 -81261
rect -42673 -81305 -42665 -81261
rect -42573 -81305 -42565 -81261
rect -42473 -81305 -42465 -81261
rect 80781 -81299 80789 -81255
rect 80881 -81299 80889 -81255
rect 80981 -81299 80989 -81255
rect 81081 -81299 81089 -81255
rect 81181 -81299 81189 -81255
rect 81281 -81299 81289 -81255
rect 81381 -81299 81389 -81255
rect 81481 -81299 81489 -81255
rect 81581 -81299 81589 -81255
rect 81681 -81299 81689 -81255
rect 81781 -81299 81789 -81255
rect 81881 -81299 81889 -81255
rect 81981 -81299 81989 -81255
rect 82081 -81299 82089 -81255
rect 82181 -81299 82189 -81255
rect 82281 -81299 82289 -81255
rect 82781 -81299 82789 -81255
rect 82881 -81299 82889 -81255
rect 82981 -81299 82989 -81255
rect 83081 -81299 83089 -81255
rect 83181 -81299 83189 -81255
rect 83281 -81299 83289 -81255
rect 83381 -81299 83389 -81255
rect 83481 -81299 83489 -81255
rect 83581 -81299 83589 -81255
rect 83681 -81299 83689 -81255
rect 83781 -81299 83789 -81255
rect 83881 -81299 83889 -81255
rect 83981 -81299 83989 -81255
rect 84081 -81299 84089 -81255
rect 84181 -81299 84189 -81255
rect 84281 -81299 84289 -81255
rect 84781 -81299 84789 -81255
rect 84881 -81299 84889 -81255
rect 84981 -81299 84989 -81255
rect 85081 -81299 85089 -81255
rect 85181 -81299 85189 -81255
rect 85281 -81299 85289 -81255
rect 85381 -81299 85389 -81255
rect 85481 -81299 85489 -81255
rect 85581 -81299 85589 -81255
rect 85681 -81299 85689 -81255
rect 85781 -81299 85789 -81255
rect 85881 -81299 85889 -81255
rect 85981 -81299 85989 -81255
rect 86081 -81299 86089 -81255
rect 86181 -81299 86189 -81255
rect 86281 -81299 86289 -81255
rect 86781 -81299 86789 -81255
rect 86881 -81299 86889 -81255
rect 86981 -81299 86989 -81255
rect 87081 -81299 87089 -81255
rect 87181 -81299 87189 -81255
rect 87281 -81299 87289 -81255
rect 87381 -81299 87389 -81255
rect 87481 -81299 87489 -81255
rect 87581 -81299 87589 -81255
rect 87681 -81299 87689 -81255
rect 87781 -81299 87789 -81255
rect 87881 -81299 87889 -81255
rect 87981 -81299 87989 -81255
rect 88081 -81299 88089 -81255
rect 88181 -81299 88189 -81255
rect 88281 -81299 88289 -81255
rect -82968 -81359 -82924 -81351
rect -82868 -81359 -82824 -81351
rect -82768 -81359 -82724 -81351
rect -82668 -81359 -82624 -81351
rect -82568 -81359 -82524 -81351
rect -82468 -81359 -82424 -81351
rect -82368 -81359 -82324 -81351
rect -82268 -81359 -82224 -81351
rect -82168 -81359 -82124 -81351
rect -82068 -81359 -82024 -81351
rect -81968 -81359 -81924 -81351
rect -81868 -81359 -81824 -81351
rect -81768 -81359 -81724 -81351
rect -81668 -81359 -81624 -81351
rect -81568 -81359 -81524 -81351
rect -81468 -81359 -81424 -81351
rect -80968 -81359 -80924 -81351
rect -80868 -81359 -80824 -81351
rect -80768 -81359 -80724 -81351
rect -80668 -81359 -80624 -81351
rect -80568 -81359 -80524 -81351
rect -80468 -81359 -80424 -81351
rect -80368 -81359 -80324 -81351
rect -80268 -81359 -80224 -81351
rect -80168 -81359 -80124 -81351
rect -80068 -81359 -80024 -81351
rect -79968 -81359 -79924 -81351
rect -79868 -81359 -79824 -81351
rect -79768 -81359 -79724 -81351
rect -79668 -81359 -79624 -81351
rect -79568 -81359 -79524 -81351
rect -79468 -81359 -79424 -81351
rect -78968 -81359 -78924 -81351
rect -78868 -81359 -78824 -81351
rect -78768 -81359 -78724 -81351
rect -78668 -81359 -78624 -81351
rect -78568 -81359 -78524 -81351
rect -78468 -81359 -78424 -81351
rect -78368 -81359 -78324 -81351
rect -78268 -81359 -78224 -81351
rect -78168 -81359 -78124 -81351
rect -78068 -81359 -78024 -81351
rect -77968 -81359 -77924 -81351
rect -77868 -81359 -77824 -81351
rect -77768 -81359 -77724 -81351
rect -77668 -81359 -77624 -81351
rect -77568 -81359 -77524 -81351
rect -77468 -81359 -77424 -81351
rect -76968 -81359 -76924 -81351
rect -76868 -81359 -76824 -81351
rect -76768 -81359 -76724 -81351
rect -76668 -81359 -76624 -81351
rect -76568 -81359 -76524 -81351
rect -76468 -81359 -76424 -81351
rect -76368 -81359 -76324 -81351
rect -76268 -81359 -76224 -81351
rect -76168 -81359 -76124 -81351
rect -76068 -81359 -76024 -81351
rect -75968 -81359 -75924 -81351
rect -75868 -81359 -75824 -81351
rect -75768 -81359 -75724 -81351
rect -75668 -81359 -75624 -81351
rect -75568 -81359 -75524 -81351
rect -75468 -81359 -75424 -81351
rect -82924 -81403 -82916 -81359
rect -82824 -81403 -82816 -81359
rect -82724 -81403 -82716 -81359
rect -82624 -81403 -82616 -81359
rect -82524 -81403 -82516 -81359
rect -82424 -81403 -82416 -81359
rect -82324 -81403 -82316 -81359
rect -82224 -81403 -82216 -81359
rect -82124 -81403 -82116 -81359
rect -82024 -81403 -82016 -81359
rect -81924 -81403 -81916 -81359
rect -81824 -81403 -81816 -81359
rect -81724 -81403 -81716 -81359
rect -81624 -81403 -81616 -81359
rect -81524 -81403 -81516 -81359
rect -81424 -81403 -81416 -81359
rect -80924 -81403 -80916 -81359
rect -80824 -81403 -80816 -81359
rect -80724 -81403 -80716 -81359
rect -80624 -81403 -80616 -81359
rect -80524 -81403 -80516 -81359
rect -80424 -81403 -80416 -81359
rect -80324 -81403 -80316 -81359
rect -80224 -81403 -80216 -81359
rect -80124 -81403 -80116 -81359
rect -80024 -81403 -80016 -81359
rect -79924 -81403 -79916 -81359
rect -79824 -81403 -79816 -81359
rect -79724 -81403 -79716 -81359
rect -79624 -81403 -79616 -81359
rect -79524 -81403 -79516 -81359
rect -79424 -81403 -79416 -81359
rect -78924 -81403 -78916 -81359
rect -78824 -81403 -78816 -81359
rect -78724 -81403 -78716 -81359
rect -78624 -81403 -78616 -81359
rect -78524 -81403 -78516 -81359
rect -78424 -81403 -78416 -81359
rect -78324 -81403 -78316 -81359
rect -78224 -81403 -78216 -81359
rect -78124 -81403 -78116 -81359
rect -78024 -81403 -78016 -81359
rect -77924 -81403 -77916 -81359
rect -77824 -81403 -77816 -81359
rect -77724 -81403 -77716 -81359
rect -77624 -81403 -77616 -81359
rect -77524 -81403 -77516 -81359
rect -77424 -81403 -77416 -81359
rect -76924 -81403 -76916 -81359
rect -76824 -81403 -76816 -81359
rect -76724 -81403 -76716 -81359
rect -76624 -81403 -76616 -81359
rect -76524 -81403 -76516 -81359
rect -76424 -81403 -76416 -81359
rect -76324 -81403 -76316 -81359
rect -76224 -81403 -76216 -81359
rect -76124 -81403 -76116 -81359
rect -76024 -81403 -76016 -81359
rect -75924 -81403 -75916 -81359
rect -75824 -81403 -75816 -81359
rect -75724 -81403 -75716 -81359
rect -75624 -81403 -75616 -81359
rect -75524 -81403 -75516 -81359
rect -75424 -81403 -75416 -81359
rect -50017 -81361 -49973 -81353
rect -49917 -81361 -49873 -81353
rect -49817 -81361 -49773 -81353
rect -49717 -81361 -49673 -81353
rect -49617 -81361 -49573 -81353
rect -49517 -81361 -49473 -81353
rect -49417 -81361 -49373 -81353
rect -49317 -81361 -49273 -81353
rect -49217 -81361 -49173 -81353
rect -49117 -81361 -49073 -81353
rect -49017 -81361 -48973 -81353
rect -48917 -81361 -48873 -81353
rect -48817 -81361 -48773 -81353
rect -48717 -81361 -48673 -81353
rect -48617 -81361 -48573 -81353
rect -48517 -81361 -48473 -81353
rect -48017 -81361 -47973 -81353
rect -47917 -81361 -47873 -81353
rect -47817 -81361 -47773 -81353
rect -47717 -81361 -47673 -81353
rect -47617 -81361 -47573 -81353
rect -47517 -81361 -47473 -81353
rect -47417 -81361 -47373 -81353
rect -47317 -81361 -47273 -81353
rect -47217 -81361 -47173 -81353
rect -47117 -81361 -47073 -81353
rect -47017 -81361 -46973 -81353
rect -46917 -81361 -46873 -81353
rect -46817 -81361 -46773 -81353
rect -46717 -81361 -46673 -81353
rect -46617 -81361 -46573 -81353
rect -46517 -81361 -46473 -81353
rect -46017 -81361 -45973 -81353
rect -45917 -81361 -45873 -81353
rect -45817 -81361 -45773 -81353
rect -45717 -81361 -45673 -81353
rect -45617 -81361 -45573 -81353
rect -45517 -81361 -45473 -81353
rect -45417 -81361 -45373 -81353
rect -45317 -81361 -45273 -81353
rect -45217 -81361 -45173 -81353
rect -45117 -81361 -45073 -81353
rect -45017 -81361 -44973 -81353
rect -44917 -81361 -44873 -81353
rect -44817 -81361 -44773 -81353
rect -44717 -81361 -44673 -81353
rect -44617 -81361 -44573 -81353
rect -44517 -81361 -44473 -81353
rect -44017 -81361 -43973 -81353
rect -43917 -81361 -43873 -81353
rect -43817 -81361 -43773 -81353
rect -43717 -81361 -43673 -81353
rect -43617 -81361 -43573 -81353
rect -43517 -81361 -43473 -81353
rect -43417 -81361 -43373 -81353
rect -43317 -81361 -43273 -81353
rect -43217 -81361 -43173 -81353
rect -43117 -81361 -43073 -81353
rect -43017 -81361 -42973 -81353
rect -42917 -81361 -42873 -81353
rect -42817 -81361 -42773 -81353
rect -42717 -81361 -42673 -81353
rect -42617 -81361 -42573 -81353
rect -42517 -81361 -42473 -81353
rect 80737 -81355 80781 -81347
rect 80837 -81355 80881 -81347
rect 80937 -81355 80981 -81347
rect 81037 -81355 81081 -81347
rect 81137 -81355 81181 -81347
rect 81237 -81355 81281 -81347
rect 81337 -81355 81381 -81347
rect 81437 -81355 81481 -81347
rect 81537 -81355 81581 -81347
rect 81637 -81355 81681 -81347
rect 81737 -81355 81781 -81347
rect 81837 -81355 81881 -81347
rect 81937 -81355 81981 -81347
rect 82037 -81355 82081 -81347
rect 82137 -81355 82181 -81347
rect 82237 -81355 82281 -81347
rect 82737 -81355 82781 -81347
rect 82837 -81355 82881 -81347
rect 82937 -81355 82981 -81347
rect 83037 -81355 83081 -81347
rect 83137 -81355 83181 -81347
rect 83237 -81355 83281 -81347
rect 83337 -81355 83381 -81347
rect 83437 -81355 83481 -81347
rect 83537 -81355 83581 -81347
rect 83637 -81355 83681 -81347
rect 83737 -81355 83781 -81347
rect 83837 -81355 83881 -81347
rect 83937 -81355 83981 -81347
rect 84037 -81355 84081 -81347
rect 84137 -81355 84181 -81347
rect 84237 -81355 84281 -81347
rect 84737 -81355 84781 -81347
rect 84837 -81355 84881 -81347
rect 84937 -81355 84981 -81347
rect 85037 -81355 85081 -81347
rect 85137 -81355 85181 -81347
rect 85237 -81355 85281 -81347
rect 85337 -81355 85381 -81347
rect 85437 -81355 85481 -81347
rect 85537 -81355 85581 -81347
rect 85637 -81355 85681 -81347
rect 85737 -81355 85781 -81347
rect 85837 -81355 85881 -81347
rect 85937 -81355 85981 -81347
rect 86037 -81355 86081 -81347
rect 86137 -81355 86181 -81347
rect 86237 -81355 86281 -81347
rect 86737 -81355 86781 -81347
rect 86837 -81355 86881 -81347
rect 86937 -81355 86981 -81347
rect 87037 -81355 87081 -81347
rect 87137 -81355 87181 -81347
rect 87237 -81355 87281 -81347
rect 87337 -81355 87381 -81347
rect 87437 -81355 87481 -81347
rect 87537 -81355 87581 -81347
rect 87637 -81355 87681 -81347
rect 87737 -81355 87781 -81347
rect 87837 -81355 87881 -81347
rect 87937 -81355 87981 -81347
rect 88037 -81355 88081 -81347
rect 88137 -81355 88181 -81347
rect 88237 -81355 88281 -81347
rect -49973 -81405 -49965 -81361
rect -49873 -81405 -49865 -81361
rect -49773 -81405 -49765 -81361
rect -49673 -81405 -49665 -81361
rect -49573 -81405 -49565 -81361
rect -49473 -81405 -49465 -81361
rect -49373 -81405 -49365 -81361
rect -49273 -81405 -49265 -81361
rect -49173 -81405 -49165 -81361
rect -49073 -81405 -49065 -81361
rect -48973 -81405 -48965 -81361
rect -48873 -81405 -48865 -81361
rect -48773 -81405 -48765 -81361
rect -48673 -81405 -48665 -81361
rect -48573 -81405 -48565 -81361
rect -48473 -81405 -48465 -81361
rect -47973 -81405 -47965 -81361
rect -47873 -81405 -47865 -81361
rect -47773 -81405 -47765 -81361
rect -47673 -81405 -47665 -81361
rect -47573 -81405 -47565 -81361
rect -47473 -81405 -47465 -81361
rect -47373 -81405 -47365 -81361
rect -47273 -81405 -47265 -81361
rect -47173 -81405 -47165 -81361
rect -47073 -81405 -47065 -81361
rect -46973 -81405 -46965 -81361
rect -46873 -81405 -46865 -81361
rect -46773 -81405 -46765 -81361
rect -46673 -81405 -46665 -81361
rect -46573 -81405 -46565 -81361
rect -46473 -81405 -46465 -81361
rect -45973 -81405 -45965 -81361
rect -45873 -81405 -45865 -81361
rect -45773 -81405 -45765 -81361
rect -45673 -81405 -45665 -81361
rect -45573 -81405 -45565 -81361
rect -45473 -81405 -45465 -81361
rect -45373 -81405 -45365 -81361
rect -45273 -81405 -45265 -81361
rect -45173 -81405 -45165 -81361
rect -45073 -81405 -45065 -81361
rect -44973 -81405 -44965 -81361
rect -44873 -81405 -44865 -81361
rect -44773 -81405 -44765 -81361
rect -44673 -81405 -44665 -81361
rect -44573 -81405 -44565 -81361
rect -44473 -81405 -44465 -81361
rect -43973 -81405 -43965 -81361
rect -43873 -81405 -43865 -81361
rect -43773 -81405 -43765 -81361
rect -43673 -81405 -43665 -81361
rect -43573 -81405 -43565 -81361
rect -43473 -81405 -43465 -81361
rect -43373 -81405 -43365 -81361
rect -43273 -81405 -43265 -81361
rect -43173 -81405 -43165 -81361
rect -43073 -81405 -43065 -81361
rect -42973 -81405 -42965 -81361
rect -42873 -81405 -42865 -81361
rect -42773 -81405 -42765 -81361
rect -42673 -81405 -42665 -81361
rect -42573 -81405 -42565 -81361
rect -42473 -81405 -42465 -81361
rect 80781 -81399 80789 -81355
rect 80881 -81399 80889 -81355
rect 80981 -81399 80989 -81355
rect 81081 -81399 81089 -81355
rect 81181 -81399 81189 -81355
rect 81281 -81399 81289 -81355
rect 81381 -81399 81389 -81355
rect 81481 -81399 81489 -81355
rect 81581 -81399 81589 -81355
rect 81681 -81399 81689 -81355
rect 81781 -81399 81789 -81355
rect 81881 -81399 81889 -81355
rect 81981 -81399 81989 -81355
rect 82081 -81399 82089 -81355
rect 82181 -81399 82189 -81355
rect 82281 -81399 82289 -81355
rect 82781 -81399 82789 -81355
rect 82881 -81399 82889 -81355
rect 82981 -81399 82989 -81355
rect 83081 -81399 83089 -81355
rect 83181 -81399 83189 -81355
rect 83281 -81399 83289 -81355
rect 83381 -81399 83389 -81355
rect 83481 -81399 83489 -81355
rect 83581 -81399 83589 -81355
rect 83681 -81399 83689 -81355
rect 83781 -81399 83789 -81355
rect 83881 -81399 83889 -81355
rect 83981 -81399 83989 -81355
rect 84081 -81399 84089 -81355
rect 84181 -81399 84189 -81355
rect 84281 -81399 84289 -81355
rect 84781 -81399 84789 -81355
rect 84881 -81399 84889 -81355
rect 84981 -81399 84989 -81355
rect 85081 -81399 85089 -81355
rect 85181 -81399 85189 -81355
rect 85281 -81399 85289 -81355
rect 85381 -81399 85389 -81355
rect 85481 -81399 85489 -81355
rect 85581 -81399 85589 -81355
rect 85681 -81399 85689 -81355
rect 85781 -81399 85789 -81355
rect 85881 -81399 85889 -81355
rect 85981 -81399 85989 -81355
rect 86081 -81399 86089 -81355
rect 86181 -81399 86189 -81355
rect 86281 -81399 86289 -81355
rect 86781 -81399 86789 -81355
rect 86881 -81399 86889 -81355
rect 86981 -81399 86989 -81355
rect 87081 -81399 87089 -81355
rect 87181 -81399 87189 -81355
rect 87281 -81399 87289 -81355
rect 87381 -81399 87389 -81355
rect 87481 -81399 87489 -81355
rect 87581 -81399 87589 -81355
rect 87681 -81399 87689 -81355
rect 87781 -81399 87789 -81355
rect 87881 -81399 87889 -81355
rect 87981 -81399 87989 -81355
rect 88081 -81399 88089 -81355
rect 88181 -81399 88189 -81355
rect 88281 -81399 88289 -81355
rect -82968 -81459 -82924 -81451
rect -82868 -81459 -82824 -81451
rect -82768 -81459 -82724 -81451
rect -82668 -81459 -82624 -81451
rect -82568 -81459 -82524 -81451
rect -82468 -81459 -82424 -81451
rect -82368 -81459 -82324 -81451
rect -82268 -81459 -82224 -81451
rect -82168 -81459 -82124 -81451
rect -82068 -81459 -82024 -81451
rect -81968 -81459 -81924 -81451
rect -81868 -81459 -81824 -81451
rect -81768 -81459 -81724 -81451
rect -81668 -81459 -81624 -81451
rect -81568 -81459 -81524 -81451
rect -81468 -81459 -81424 -81451
rect -80968 -81459 -80924 -81451
rect -80868 -81459 -80824 -81451
rect -80768 -81459 -80724 -81451
rect -80668 -81459 -80624 -81451
rect -80568 -81459 -80524 -81451
rect -80468 -81459 -80424 -81451
rect -80368 -81459 -80324 -81451
rect -80268 -81459 -80224 -81451
rect -80168 -81459 -80124 -81451
rect -80068 -81459 -80024 -81451
rect -79968 -81459 -79924 -81451
rect -79868 -81459 -79824 -81451
rect -79768 -81459 -79724 -81451
rect -79668 -81459 -79624 -81451
rect -79568 -81459 -79524 -81451
rect -79468 -81459 -79424 -81451
rect -78968 -81459 -78924 -81451
rect -78868 -81459 -78824 -81451
rect -78768 -81459 -78724 -81451
rect -78668 -81459 -78624 -81451
rect -78568 -81459 -78524 -81451
rect -78468 -81459 -78424 -81451
rect -78368 -81459 -78324 -81451
rect -78268 -81459 -78224 -81451
rect -78168 -81459 -78124 -81451
rect -78068 -81459 -78024 -81451
rect -77968 -81459 -77924 -81451
rect -77868 -81459 -77824 -81451
rect -77768 -81459 -77724 -81451
rect -77668 -81459 -77624 -81451
rect -77568 -81459 -77524 -81451
rect -77468 -81459 -77424 -81451
rect -76968 -81459 -76924 -81451
rect -76868 -81459 -76824 -81451
rect -76768 -81459 -76724 -81451
rect -76668 -81459 -76624 -81451
rect -76568 -81459 -76524 -81451
rect -76468 -81459 -76424 -81451
rect -76368 -81459 -76324 -81451
rect -76268 -81459 -76224 -81451
rect -76168 -81459 -76124 -81451
rect -76068 -81459 -76024 -81451
rect -75968 -81459 -75924 -81451
rect -75868 -81459 -75824 -81451
rect -75768 -81459 -75724 -81451
rect -75668 -81459 -75624 -81451
rect -75568 -81459 -75524 -81451
rect -75468 -81459 -75424 -81451
rect -82924 -81503 -82916 -81459
rect -82824 -81503 -82816 -81459
rect -82724 -81503 -82716 -81459
rect -82624 -81503 -82616 -81459
rect -82524 -81503 -82516 -81459
rect -82424 -81503 -82416 -81459
rect -82324 -81503 -82316 -81459
rect -82224 -81503 -82216 -81459
rect -82124 -81503 -82116 -81459
rect -82024 -81503 -82016 -81459
rect -81924 -81503 -81916 -81459
rect -81824 -81503 -81816 -81459
rect -81724 -81503 -81716 -81459
rect -81624 -81503 -81616 -81459
rect -81524 -81503 -81516 -81459
rect -81424 -81503 -81416 -81459
rect -80924 -81503 -80916 -81459
rect -80824 -81503 -80816 -81459
rect -80724 -81503 -80716 -81459
rect -80624 -81503 -80616 -81459
rect -80524 -81503 -80516 -81459
rect -80424 -81503 -80416 -81459
rect -80324 -81503 -80316 -81459
rect -80224 -81503 -80216 -81459
rect -80124 -81503 -80116 -81459
rect -80024 -81503 -80016 -81459
rect -79924 -81503 -79916 -81459
rect -79824 -81503 -79816 -81459
rect -79724 -81503 -79716 -81459
rect -79624 -81503 -79616 -81459
rect -79524 -81503 -79516 -81459
rect -79424 -81503 -79416 -81459
rect -78924 -81503 -78916 -81459
rect -78824 -81503 -78816 -81459
rect -78724 -81503 -78716 -81459
rect -78624 -81503 -78616 -81459
rect -78524 -81503 -78516 -81459
rect -78424 -81503 -78416 -81459
rect -78324 -81503 -78316 -81459
rect -78224 -81503 -78216 -81459
rect -78124 -81503 -78116 -81459
rect -78024 -81503 -78016 -81459
rect -77924 -81503 -77916 -81459
rect -77824 -81503 -77816 -81459
rect -77724 -81503 -77716 -81459
rect -77624 -81503 -77616 -81459
rect -77524 -81503 -77516 -81459
rect -77424 -81503 -77416 -81459
rect -76924 -81503 -76916 -81459
rect -76824 -81503 -76816 -81459
rect -76724 -81503 -76716 -81459
rect -76624 -81503 -76616 -81459
rect -76524 -81503 -76516 -81459
rect -76424 -81503 -76416 -81459
rect -76324 -81503 -76316 -81459
rect -76224 -81503 -76216 -81459
rect -76124 -81503 -76116 -81459
rect -76024 -81503 -76016 -81459
rect -75924 -81503 -75916 -81459
rect -75824 -81503 -75816 -81459
rect -75724 -81503 -75716 -81459
rect -75624 -81503 -75616 -81459
rect -75524 -81503 -75516 -81459
rect -75424 -81503 -75416 -81459
rect -50017 -81461 -49973 -81453
rect -49917 -81461 -49873 -81453
rect -49817 -81461 -49773 -81453
rect -49717 -81461 -49673 -81453
rect -49617 -81461 -49573 -81453
rect -49517 -81461 -49473 -81453
rect -49417 -81461 -49373 -81453
rect -49317 -81461 -49273 -81453
rect -49217 -81461 -49173 -81453
rect -49117 -81461 -49073 -81453
rect -49017 -81461 -48973 -81453
rect -48917 -81461 -48873 -81453
rect -48817 -81461 -48773 -81453
rect -48717 -81461 -48673 -81453
rect -48617 -81461 -48573 -81453
rect -48517 -81461 -48473 -81453
rect -48017 -81461 -47973 -81453
rect -47917 -81461 -47873 -81453
rect -47817 -81461 -47773 -81453
rect -47717 -81461 -47673 -81453
rect -47617 -81461 -47573 -81453
rect -47517 -81461 -47473 -81453
rect -47417 -81461 -47373 -81453
rect -47317 -81461 -47273 -81453
rect -47217 -81461 -47173 -81453
rect -47117 -81461 -47073 -81453
rect -47017 -81461 -46973 -81453
rect -46917 -81461 -46873 -81453
rect -46817 -81461 -46773 -81453
rect -46717 -81461 -46673 -81453
rect -46617 -81461 -46573 -81453
rect -46517 -81461 -46473 -81453
rect -46017 -81461 -45973 -81453
rect -45917 -81461 -45873 -81453
rect -45817 -81461 -45773 -81453
rect -45717 -81461 -45673 -81453
rect -45617 -81461 -45573 -81453
rect -45517 -81461 -45473 -81453
rect -45417 -81461 -45373 -81453
rect -45317 -81461 -45273 -81453
rect -45217 -81461 -45173 -81453
rect -45117 -81461 -45073 -81453
rect -45017 -81461 -44973 -81453
rect -44917 -81461 -44873 -81453
rect -44817 -81461 -44773 -81453
rect -44717 -81461 -44673 -81453
rect -44617 -81461 -44573 -81453
rect -44517 -81461 -44473 -81453
rect -44017 -81461 -43973 -81453
rect -43917 -81461 -43873 -81453
rect -43817 -81461 -43773 -81453
rect -43717 -81461 -43673 -81453
rect -43617 -81461 -43573 -81453
rect -43517 -81461 -43473 -81453
rect -43417 -81461 -43373 -81453
rect -43317 -81461 -43273 -81453
rect -43217 -81461 -43173 -81453
rect -43117 -81461 -43073 -81453
rect -43017 -81461 -42973 -81453
rect -42917 -81461 -42873 -81453
rect -42817 -81461 -42773 -81453
rect -42717 -81461 -42673 -81453
rect -42617 -81461 -42573 -81453
rect -42517 -81461 -42473 -81453
rect 80737 -81455 80781 -81447
rect 80837 -81455 80881 -81447
rect 80937 -81455 80981 -81447
rect 81037 -81455 81081 -81447
rect 81137 -81455 81181 -81447
rect 81237 -81455 81281 -81447
rect 81337 -81455 81381 -81447
rect 81437 -81455 81481 -81447
rect 81537 -81455 81581 -81447
rect 81637 -81455 81681 -81447
rect 81737 -81455 81781 -81447
rect 81837 -81455 81881 -81447
rect 81937 -81455 81981 -81447
rect 82037 -81455 82081 -81447
rect 82137 -81455 82181 -81447
rect 82237 -81455 82281 -81447
rect 82737 -81455 82781 -81447
rect 82837 -81455 82881 -81447
rect 82937 -81455 82981 -81447
rect 83037 -81455 83081 -81447
rect 83137 -81455 83181 -81447
rect 83237 -81455 83281 -81447
rect 83337 -81455 83381 -81447
rect 83437 -81455 83481 -81447
rect 83537 -81455 83581 -81447
rect 83637 -81455 83681 -81447
rect 83737 -81455 83781 -81447
rect 83837 -81455 83881 -81447
rect 83937 -81455 83981 -81447
rect 84037 -81455 84081 -81447
rect 84137 -81455 84181 -81447
rect 84237 -81455 84281 -81447
rect 84737 -81455 84781 -81447
rect 84837 -81455 84881 -81447
rect 84937 -81455 84981 -81447
rect 85037 -81455 85081 -81447
rect 85137 -81455 85181 -81447
rect 85237 -81455 85281 -81447
rect 85337 -81455 85381 -81447
rect 85437 -81455 85481 -81447
rect 85537 -81455 85581 -81447
rect 85637 -81455 85681 -81447
rect 85737 -81455 85781 -81447
rect 85837 -81455 85881 -81447
rect 85937 -81455 85981 -81447
rect 86037 -81455 86081 -81447
rect 86137 -81455 86181 -81447
rect 86237 -81455 86281 -81447
rect 86737 -81455 86781 -81447
rect 86837 -81455 86881 -81447
rect 86937 -81455 86981 -81447
rect 87037 -81455 87081 -81447
rect 87137 -81455 87181 -81447
rect 87237 -81455 87281 -81447
rect 87337 -81455 87381 -81447
rect 87437 -81455 87481 -81447
rect 87537 -81455 87581 -81447
rect 87637 -81455 87681 -81447
rect 87737 -81455 87781 -81447
rect 87837 -81455 87881 -81447
rect 87937 -81455 87981 -81447
rect 88037 -81455 88081 -81447
rect 88137 -81455 88181 -81447
rect 88237 -81455 88281 -81447
rect -49973 -81505 -49965 -81461
rect -49873 -81505 -49865 -81461
rect -49773 -81505 -49765 -81461
rect -49673 -81505 -49665 -81461
rect -49573 -81505 -49565 -81461
rect -49473 -81505 -49465 -81461
rect -49373 -81505 -49365 -81461
rect -49273 -81505 -49265 -81461
rect -49173 -81505 -49165 -81461
rect -49073 -81505 -49065 -81461
rect -48973 -81505 -48965 -81461
rect -48873 -81505 -48865 -81461
rect -48773 -81505 -48765 -81461
rect -48673 -81505 -48665 -81461
rect -48573 -81505 -48565 -81461
rect -48473 -81505 -48465 -81461
rect -47973 -81505 -47965 -81461
rect -47873 -81505 -47865 -81461
rect -47773 -81505 -47765 -81461
rect -47673 -81505 -47665 -81461
rect -47573 -81505 -47565 -81461
rect -47473 -81505 -47465 -81461
rect -47373 -81505 -47365 -81461
rect -47273 -81505 -47265 -81461
rect -47173 -81505 -47165 -81461
rect -47073 -81505 -47065 -81461
rect -46973 -81505 -46965 -81461
rect -46873 -81505 -46865 -81461
rect -46773 -81505 -46765 -81461
rect -46673 -81505 -46665 -81461
rect -46573 -81505 -46565 -81461
rect -46473 -81505 -46465 -81461
rect -45973 -81505 -45965 -81461
rect -45873 -81505 -45865 -81461
rect -45773 -81505 -45765 -81461
rect -45673 -81505 -45665 -81461
rect -45573 -81505 -45565 -81461
rect -45473 -81505 -45465 -81461
rect -45373 -81505 -45365 -81461
rect -45273 -81505 -45265 -81461
rect -45173 -81505 -45165 -81461
rect -45073 -81505 -45065 -81461
rect -44973 -81505 -44965 -81461
rect -44873 -81505 -44865 -81461
rect -44773 -81505 -44765 -81461
rect -44673 -81505 -44665 -81461
rect -44573 -81505 -44565 -81461
rect -44473 -81505 -44465 -81461
rect -43973 -81505 -43965 -81461
rect -43873 -81505 -43865 -81461
rect -43773 -81505 -43765 -81461
rect -43673 -81505 -43665 -81461
rect -43573 -81505 -43565 -81461
rect -43473 -81505 -43465 -81461
rect -43373 -81505 -43365 -81461
rect -43273 -81505 -43265 -81461
rect -43173 -81505 -43165 -81461
rect -43073 -81505 -43065 -81461
rect -42973 -81505 -42965 -81461
rect -42873 -81505 -42865 -81461
rect -42773 -81505 -42765 -81461
rect -42673 -81505 -42665 -81461
rect -42573 -81505 -42565 -81461
rect -42473 -81505 -42465 -81461
rect 80781 -81499 80789 -81455
rect 80881 -81499 80889 -81455
rect 80981 -81499 80989 -81455
rect 81081 -81499 81089 -81455
rect 81181 -81499 81189 -81455
rect 81281 -81499 81289 -81455
rect 81381 -81499 81389 -81455
rect 81481 -81499 81489 -81455
rect 81581 -81499 81589 -81455
rect 81681 -81499 81689 -81455
rect 81781 -81499 81789 -81455
rect 81881 -81499 81889 -81455
rect 81981 -81499 81989 -81455
rect 82081 -81499 82089 -81455
rect 82181 -81499 82189 -81455
rect 82281 -81499 82289 -81455
rect 82781 -81499 82789 -81455
rect 82881 -81499 82889 -81455
rect 82981 -81499 82989 -81455
rect 83081 -81499 83089 -81455
rect 83181 -81499 83189 -81455
rect 83281 -81499 83289 -81455
rect 83381 -81499 83389 -81455
rect 83481 -81499 83489 -81455
rect 83581 -81499 83589 -81455
rect 83681 -81499 83689 -81455
rect 83781 -81499 83789 -81455
rect 83881 -81499 83889 -81455
rect 83981 -81499 83989 -81455
rect 84081 -81499 84089 -81455
rect 84181 -81499 84189 -81455
rect 84281 -81499 84289 -81455
rect 84781 -81499 84789 -81455
rect 84881 -81499 84889 -81455
rect 84981 -81499 84989 -81455
rect 85081 -81499 85089 -81455
rect 85181 -81499 85189 -81455
rect 85281 -81499 85289 -81455
rect 85381 -81499 85389 -81455
rect 85481 -81499 85489 -81455
rect 85581 -81499 85589 -81455
rect 85681 -81499 85689 -81455
rect 85781 -81499 85789 -81455
rect 85881 -81499 85889 -81455
rect 85981 -81499 85989 -81455
rect 86081 -81499 86089 -81455
rect 86181 -81499 86189 -81455
rect 86281 -81499 86289 -81455
rect 86781 -81499 86789 -81455
rect 86881 -81499 86889 -81455
rect 86981 -81499 86989 -81455
rect 87081 -81499 87089 -81455
rect 87181 -81499 87189 -81455
rect 87281 -81499 87289 -81455
rect 87381 -81499 87389 -81455
rect 87481 -81499 87489 -81455
rect 87581 -81499 87589 -81455
rect 87681 -81499 87689 -81455
rect 87781 -81499 87789 -81455
rect 87881 -81499 87889 -81455
rect 87981 -81499 87989 -81455
rect 88081 -81499 88089 -81455
rect 88181 -81499 88189 -81455
rect 88281 -81499 88289 -81455
rect -82968 -81559 -82924 -81551
rect -82868 -81559 -82824 -81551
rect -82768 -81559 -82724 -81551
rect -82668 -81559 -82624 -81551
rect -82568 -81559 -82524 -81551
rect -82468 -81559 -82424 -81551
rect -82368 -81559 -82324 -81551
rect -82268 -81559 -82224 -81551
rect -82168 -81559 -82124 -81551
rect -82068 -81559 -82024 -81551
rect -81968 -81559 -81924 -81551
rect -81868 -81559 -81824 -81551
rect -81768 -81559 -81724 -81551
rect -81668 -81559 -81624 -81551
rect -81568 -81559 -81524 -81551
rect -81468 -81559 -81424 -81551
rect -80968 -81559 -80924 -81551
rect -80868 -81559 -80824 -81551
rect -80768 -81559 -80724 -81551
rect -80668 -81559 -80624 -81551
rect -80568 -81559 -80524 -81551
rect -80468 -81559 -80424 -81551
rect -80368 -81559 -80324 -81551
rect -80268 -81559 -80224 -81551
rect -80168 -81559 -80124 -81551
rect -80068 -81559 -80024 -81551
rect -79968 -81559 -79924 -81551
rect -79868 -81559 -79824 -81551
rect -79768 -81559 -79724 -81551
rect -79668 -81559 -79624 -81551
rect -79568 -81559 -79524 -81551
rect -79468 -81559 -79424 -81551
rect -78968 -81559 -78924 -81551
rect -78868 -81559 -78824 -81551
rect -78768 -81559 -78724 -81551
rect -78668 -81559 -78624 -81551
rect -78568 -81559 -78524 -81551
rect -78468 -81559 -78424 -81551
rect -78368 -81559 -78324 -81551
rect -78268 -81559 -78224 -81551
rect -78168 -81559 -78124 -81551
rect -78068 -81559 -78024 -81551
rect -77968 -81559 -77924 -81551
rect -77868 -81559 -77824 -81551
rect -77768 -81559 -77724 -81551
rect -77668 -81559 -77624 -81551
rect -77568 -81559 -77524 -81551
rect -77468 -81559 -77424 -81551
rect -76968 -81559 -76924 -81551
rect -76868 -81559 -76824 -81551
rect -76768 -81559 -76724 -81551
rect -76668 -81559 -76624 -81551
rect -76568 -81559 -76524 -81551
rect -76468 -81559 -76424 -81551
rect -76368 -81559 -76324 -81551
rect -76268 -81559 -76224 -81551
rect -76168 -81559 -76124 -81551
rect -76068 -81559 -76024 -81551
rect -75968 -81559 -75924 -81551
rect -75868 -81559 -75824 -81551
rect -75768 -81559 -75724 -81551
rect -75668 -81559 -75624 -81551
rect -75568 -81559 -75524 -81551
rect -75468 -81559 -75424 -81551
rect -82924 -81603 -82916 -81559
rect -82824 -81603 -82816 -81559
rect -82724 -81603 -82716 -81559
rect -82624 -81603 -82616 -81559
rect -82524 -81603 -82516 -81559
rect -82424 -81603 -82416 -81559
rect -82324 -81603 -82316 -81559
rect -82224 -81603 -82216 -81559
rect -82124 -81603 -82116 -81559
rect -82024 -81603 -82016 -81559
rect -81924 -81603 -81916 -81559
rect -81824 -81603 -81816 -81559
rect -81724 -81603 -81716 -81559
rect -81624 -81603 -81616 -81559
rect -81524 -81603 -81516 -81559
rect -81424 -81603 -81416 -81559
rect -80924 -81603 -80916 -81559
rect -80824 -81603 -80816 -81559
rect -80724 -81603 -80716 -81559
rect -80624 -81603 -80616 -81559
rect -80524 -81603 -80516 -81559
rect -80424 -81603 -80416 -81559
rect -80324 -81603 -80316 -81559
rect -80224 -81603 -80216 -81559
rect -80124 -81603 -80116 -81559
rect -80024 -81603 -80016 -81559
rect -79924 -81603 -79916 -81559
rect -79824 -81603 -79816 -81559
rect -79724 -81603 -79716 -81559
rect -79624 -81603 -79616 -81559
rect -79524 -81603 -79516 -81559
rect -79424 -81603 -79416 -81559
rect -78924 -81603 -78916 -81559
rect -78824 -81603 -78816 -81559
rect -78724 -81603 -78716 -81559
rect -78624 -81603 -78616 -81559
rect -78524 -81603 -78516 -81559
rect -78424 -81603 -78416 -81559
rect -78324 -81603 -78316 -81559
rect -78224 -81603 -78216 -81559
rect -78124 -81603 -78116 -81559
rect -78024 -81603 -78016 -81559
rect -77924 -81603 -77916 -81559
rect -77824 -81603 -77816 -81559
rect -77724 -81603 -77716 -81559
rect -77624 -81603 -77616 -81559
rect -77524 -81603 -77516 -81559
rect -77424 -81603 -77416 -81559
rect -76924 -81603 -76916 -81559
rect -76824 -81603 -76816 -81559
rect -76724 -81603 -76716 -81559
rect -76624 -81603 -76616 -81559
rect -76524 -81603 -76516 -81559
rect -76424 -81603 -76416 -81559
rect -76324 -81603 -76316 -81559
rect -76224 -81603 -76216 -81559
rect -76124 -81603 -76116 -81559
rect -76024 -81603 -76016 -81559
rect -75924 -81603 -75916 -81559
rect -75824 -81603 -75816 -81559
rect -75724 -81603 -75716 -81559
rect -75624 -81603 -75616 -81559
rect -75524 -81603 -75516 -81559
rect -75424 -81603 -75416 -81559
rect -50017 -81561 -49973 -81553
rect -49917 -81561 -49873 -81553
rect -49817 -81561 -49773 -81553
rect -49717 -81561 -49673 -81553
rect -49617 -81561 -49573 -81553
rect -49517 -81561 -49473 -81553
rect -49417 -81561 -49373 -81553
rect -49317 -81561 -49273 -81553
rect -49217 -81561 -49173 -81553
rect -49117 -81561 -49073 -81553
rect -49017 -81561 -48973 -81553
rect -48917 -81561 -48873 -81553
rect -48817 -81561 -48773 -81553
rect -48717 -81561 -48673 -81553
rect -48617 -81561 -48573 -81553
rect -48517 -81561 -48473 -81553
rect -48017 -81561 -47973 -81553
rect -47917 -81561 -47873 -81553
rect -47817 -81561 -47773 -81553
rect -47717 -81561 -47673 -81553
rect -47617 -81561 -47573 -81553
rect -47517 -81561 -47473 -81553
rect -47417 -81561 -47373 -81553
rect -47317 -81561 -47273 -81553
rect -47217 -81561 -47173 -81553
rect -47117 -81561 -47073 -81553
rect -47017 -81561 -46973 -81553
rect -46917 -81561 -46873 -81553
rect -46817 -81561 -46773 -81553
rect -46717 -81561 -46673 -81553
rect -46617 -81561 -46573 -81553
rect -46517 -81561 -46473 -81553
rect -46017 -81561 -45973 -81553
rect -45917 -81561 -45873 -81553
rect -45817 -81561 -45773 -81553
rect -45717 -81561 -45673 -81553
rect -45617 -81561 -45573 -81553
rect -45517 -81561 -45473 -81553
rect -45417 -81561 -45373 -81553
rect -45317 -81561 -45273 -81553
rect -45217 -81561 -45173 -81553
rect -45117 -81561 -45073 -81553
rect -45017 -81561 -44973 -81553
rect -44917 -81561 -44873 -81553
rect -44817 -81561 -44773 -81553
rect -44717 -81561 -44673 -81553
rect -44617 -81561 -44573 -81553
rect -44517 -81561 -44473 -81553
rect -44017 -81561 -43973 -81553
rect -43917 -81561 -43873 -81553
rect -43817 -81561 -43773 -81553
rect -43717 -81561 -43673 -81553
rect -43617 -81561 -43573 -81553
rect -43517 -81561 -43473 -81553
rect -43417 -81561 -43373 -81553
rect -43317 -81561 -43273 -81553
rect -43217 -81561 -43173 -81553
rect -43117 -81561 -43073 -81553
rect -43017 -81561 -42973 -81553
rect -42917 -81561 -42873 -81553
rect -42817 -81561 -42773 -81553
rect -42717 -81561 -42673 -81553
rect -42617 -81561 -42573 -81553
rect -42517 -81561 -42473 -81553
rect 80737 -81555 80781 -81547
rect 80837 -81555 80881 -81547
rect 80937 -81555 80981 -81547
rect 81037 -81555 81081 -81547
rect 81137 -81555 81181 -81547
rect 81237 -81555 81281 -81547
rect 81337 -81555 81381 -81547
rect 81437 -81555 81481 -81547
rect 81537 -81555 81581 -81547
rect 81637 -81555 81681 -81547
rect 81737 -81555 81781 -81547
rect 81837 -81555 81881 -81547
rect 81937 -81555 81981 -81547
rect 82037 -81555 82081 -81547
rect 82137 -81555 82181 -81547
rect 82237 -81555 82281 -81547
rect 82737 -81555 82781 -81547
rect 82837 -81555 82881 -81547
rect 82937 -81555 82981 -81547
rect 83037 -81555 83081 -81547
rect 83137 -81555 83181 -81547
rect 83237 -81555 83281 -81547
rect 83337 -81555 83381 -81547
rect 83437 -81555 83481 -81547
rect 83537 -81555 83581 -81547
rect 83637 -81555 83681 -81547
rect 83737 -81555 83781 -81547
rect 83837 -81555 83881 -81547
rect 83937 -81555 83981 -81547
rect 84037 -81555 84081 -81547
rect 84137 -81555 84181 -81547
rect 84237 -81555 84281 -81547
rect 84737 -81555 84781 -81547
rect 84837 -81555 84881 -81547
rect 84937 -81555 84981 -81547
rect 85037 -81555 85081 -81547
rect 85137 -81555 85181 -81547
rect 85237 -81555 85281 -81547
rect 85337 -81555 85381 -81547
rect 85437 -81555 85481 -81547
rect 85537 -81555 85581 -81547
rect 85637 -81555 85681 -81547
rect 85737 -81555 85781 -81547
rect 85837 -81555 85881 -81547
rect 85937 -81555 85981 -81547
rect 86037 -81555 86081 -81547
rect 86137 -81555 86181 -81547
rect 86237 -81555 86281 -81547
rect 86737 -81555 86781 -81547
rect 86837 -81555 86881 -81547
rect 86937 -81555 86981 -81547
rect 87037 -81555 87081 -81547
rect 87137 -81555 87181 -81547
rect 87237 -81555 87281 -81547
rect 87337 -81555 87381 -81547
rect 87437 -81555 87481 -81547
rect 87537 -81555 87581 -81547
rect 87637 -81555 87681 -81547
rect 87737 -81555 87781 -81547
rect 87837 -81555 87881 -81547
rect 87937 -81555 87981 -81547
rect 88037 -81555 88081 -81547
rect 88137 -81555 88181 -81547
rect 88237 -81555 88281 -81547
rect -49973 -81605 -49965 -81561
rect -49873 -81605 -49865 -81561
rect -49773 -81605 -49765 -81561
rect -49673 -81605 -49665 -81561
rect -49573 -81605 -49565 -81561
rect -49473 -81605 -49465 -81561
rect -49373 -81605 -49365 -81561
rect -49273 -81605 -49265 -81561
rect -49173 -81605 -49165 -81561
rect -49073 -81605 -49065 -81561
rect -48973 -81605 -48965 -81561
rect -48873 -81605 -48865 -81561
rect -48773 -81605 -48765 -81561
rect -48673 -81605 -48665 -81561
rect -48573 -81605 -48565 -81561
rect -48473 -81605 -48465 -81561
rect -47973 -81605 -47965 -81561
rect -47873 -81605 -47865 -81561
rect -47773 -81605 -47765 -81561
rect -47673 -81605 -47665 -81561
rect -47573 -81605 -47565 -81561
rect -47473 -81605 -47465 -81561
rect -47373 -81605 -47365 -81561
rect -47273 -81605 -47265 -81561
rect -47173 -81605 -47165 -81561
rect -47073 -81605 -47065 -81561
rect -46973 -81605 -46965 -81561
rect -46873 -81605 -46865 -81561
rect -46773 -81605 -46765 -81561
rect -46673 -81605 -46665 -81561
rect -46573 -81605 -46565 -81561
rect -46473 -81605 -46465 -81561
rect -45973 -81605 -45965 -81561
rect -45873 -81605 -45865 -81561
rect -45773 -81605 -45765 -81561
rect -45673 -81605 -45665 -81561
rect -45573 -81605 -45565 -81561
rect -45473 -81605 -45465 -81561
rect -45373 -81605 -45365 -81561
rect -45273 -81605 -45265 -81561
rect -45173 -81605 -45165 -81561
rect -45073 -81605 -45065 -81561
rect -44973 -81605 -44965 -81561
rect -44873 -81605 -44865 -81561
rect -44773 -81605 -44765 -81561
rect -44673 -81605 -44665 -81561
rect -44573 -81605 -44565 -81561
rect -44473 -81605 -44465 -81561
rect -43973 -81605 -43965 -81561
rect -43873 -81605 -43865 -81561
rect -43773 -81605 -43765 -81561
rect -43673 -81605 -43665 -81561
rect -43573 -81605 -43565 -81561
rect -43473 -81605 -43465 -81561
rect -43373 -81605 -43365 -81561
rect -43273 -81605 -43265 -81561
rect -43173 -81605 -43165 -81561
rect -43073 -81605 -43065 -81561
rect -42973 -81605 -42965 -81561
rect -42873 -81605 -42865 -81561
rect -42773 -81605 -42765 -81561
rect -42673 -81605 -42665 -81561
rect -42573 -81605 -42565 -81561
rect -42473 -81605 -42465 -81561
rect 80781 -81599 80789 -81555
rect 80881 -81599 80889 -81555
rect 80981 -81599 80989 -81555
rect 81081 -81599 81089 -81555
rect 81181 -81599 81189 -81555
rect 81281 -81599 81289 -81555
rect 81381 -81599 81389 -81555
rect 81481 -81599 81489 -81555
rect 81581 -81599 81589 -81555
rect 81681 -81599 81689 -81555
rect 81781 -81599 81789 -81555
rect 81881 -81599 81889 -81555
rect 81981 -81599 81989 -81555
rect 82081 -81599 82089 -81555
rect 82181 -81599 82189 -81555
rect 82281 -81599 82289 -81555
rect 82781 -81599 82789 -81555
rect 82881 -81599 82889 -81555
rect 82981 -81599 82989 -81555
rect 83081 -81599 83089 -81555
rect 83181 -81599 83189 -81555
rect 83281 -81599 83289 -81555
rect 83381 -81599 83389 -81555
rect 83481 -81599 83489 -81555
rect 83581 -81599 83589 -81555
rect 83681 -81599 83689 -81555
rect 83781 -81599 83789 -81555
rect 83881 -81599 83889 -81555
rect 83981 -81599 83989 -81555
rect 84081 -81599 84089 -81555
rect 84181 -81599 84189 -81555
rect 84281 -81599 84289 -81555
rect 84781 -81599 84789 -81555
rect 84881 -81599 84889 -81555
rect 84981 -81599 84989 -81555
rect 85081 -81599 85089 -81555
rect 85181 -81599 85189 -81555
rect 85281 -81599 85289 -81555
rect 85381 -81599 85389 -81555
rect 85481 -81599 85489 -81555
rect 85581 -81599 85589 -81555
rect 85681 -81599 85689 -81555
rect 85781 -81599 85789 -81555
rect 85881 -81599 85889 -81555
rect 85981 -81599 85989 -81555
rect 86081 -81599 86089 -81555
rect 86181 -81599 86189 -81555
rect 86281 -81599 86289 -81555
rect 86781 -81599 86789 -81555
rect 86881 -81599 86889 -81555
rect 86981 -81599 86989 -81555
rect 87081 -81599 87089 -81555
rect 87181 -81599 87189 -81555
rect 87281 -81599 87289 -81555
rect 87381 -81599 87389 -81555
rect 87481 -81599 87489 -81555
rect 87581 -81599 87589 -81555
rect 87681 -81599 87689 -81555
rect 87781 -81599 87789 -81555
rect 87881 -81599 87889 -81555
rect 87981 -81599 87989 -81555
rect 88081 -81599 88089 -81555
rect 88181 -81599 88189 -81555
rect 88281 -81599 88289 -81555
rect -82968 -81659 -82924 -81651
rect -82868 -81659 -82824 -81651
rect -82768 -81659 -82724 -81651
rect -82668 -81659 -82624 -81651
rect -82568 -81659 -82524 -81651
rect -82468 -81659 -82424 -81651
rect -82368 -81659 -82324 -81651
rect -82268 -81659 -82224 -81651
rect -82168 -81659 -82124 -81651
rect -82068 -81659 -82024 -81651
rect -81968 -81659 -81924 -81651
rect -81868 -81659 -81824 -81651
rect -81768 -81659 -81724 -81651
rect -81668 -81659 -81624 -81651
rect -81568 -81659 -81524 -81651
rect -81468 -81659 -81424 -81651
rect -80968 -81659 -80924 -81651
rect -80868 -81659 -80824 -81651
rect -80768 -81659 -80724 -81651
rect -80668 -81659 -80624 -81651
rect -80568 -81659 -80524 -81651
rect -80468 -81659 -80424 -81651
rect -80368 -81659 -80324 -81651
rect -80268 -81659 -80224 -81651
rect -80168 -81659 -80124 -81651
rect -80068 -81659 -80024 -81651
rect -79968 -81659 -79924 -81651
rect -79868 -81659 -79824 -81651
rect -79768 -81659 -79724 -81651
rect -79668 -81659 -79624 -81651
rect -79568 -81659 -79524 -81651
rect -79468 -81659 -79424 -81651
rect -78968 -81659 -78924 -81651
rect -78868 -81659 -78824 -81651
rect -78768 -81659 -78724 -81651
rect -78668 -81659 -78624 -81651
rect -78568 -81659 -78524 -81651
rect -78468 -81659 -78424 -81651
rect -78368 -81659 -78324 -81651
rect -78268 -81659 -78224 -81651
rect -78168 -81659 -78124 -81651
rect -78068 -81659 -78024 -81651
rect -77968 -81659 -77924 -81651
rect -77868 -81659 -77824 -81651
rect -77768 -81659 -77724 -81651
rect -77668 -81659 -77624 -81651
rect -77568 -81659 -77524 -81651
rect -77468 -81659 -77424 -81651
rect -76968 -81659 -76924 -81651
rect -76868 -81659 -76824 -81651
rect -76768 -81659 -76724 -81651
rect -76668 -81659 -76624 -81651
rect -76568 -81659 -76524 -81651
rect -76468 -81659 -76424 -81651
rect -76368 -81659 -76324 -81651
rect -76268 -81659 -76224 -81651
rect -76168 -81659 -76124 -81651
rect -76068 -81659 -76024 -81651
rect -75968 -81659 -75924 -81651
rect -75868 -81659 -75824 -81651
rect -75768 -81659 -75724 -81651
rect -75668 -81659 -75624 -81651
rect -75568 -81659 -75524 -81651
rect -75468 -81659 -75424 -81651
rect -82924 -81703 -82916 -81659
rect -82824 -81703 -82816 -81659
rect -82724 -81703 -82716 -81659
rect -82624 -81703 -82616 -81659
rect -82524 -81703 -82516 -81659
rect -82424 -81703 -82416 -81659
rect -82324 -81703 -82316 -81659
rect -82224 -81703 -82216 -81659
rect -82124 -81703 -82116 -81659
rect -82024 -81703 -82016 -81659
rect -81924 -81703 -81916 -81659
rect -81824 -81703 -81816 -81659
rect -81724 -81703 -81716 -81659
rect -81624 -81703 -81616 -81659
rect -81524 -81703 -81516 -81659
rect -81424 -81703 -81416 -81659
rect -80924 -81703 -80916 -81659
rect -80824 -81703 -80816 -81659
rect -80724 -81703 -80716 -81659
rect -80624 -81703 -80616 -81659
rect -80524 -81703 -80516 -81659
rect -80424 -81703 -80416 -81659
rect -80324 -81703 -80316 -81659
rect -80224 -81703 -80216 -81659
rect -80124 -81703 -80116 -81659
rect -80024 -81703 -80016 -81659
rect -79924 -81703 -79916 -81659
rect -79824 -81703 -79816 -81659
rect -79724 -81703 -79716 -81659
rect -79624 -81703 -79616 -81659
rect -79524 -81703 -79516 -81659
rect -79424 -81703 -79416 -81659
rect -78924 -81703 -78916 -81659
rect -78824 -81703 -78816 -81659
rect -78724 -81703 -78716 -81659
rect -78624 -81703 -78616 -81659
rect -78524 -81703 -78516 -81659
rect -78424 -81703 -78416 -81659
rect -78324 -81703 -78316 -81659
rect -78224 -81703 -78216 -81659
rect -78124 -81703 -78116 -81659
rect -78024 -81703 -78016 -81659
rect -77924 -81703 -77916 -81659
rect -77824 -81703 -77816 -81659
rect -77724 -81703 -77716 -81659
rect -77624 -81703 -77616 -81659
rect -77524 -81703 -77516 -81659
rect -77424 -81703 -77416 -81659
rect -76924 -81703 -76916 -81659
rect -76824 -81703 -76816 -81659
rect -76724 -81703 -76716 -81659
rect -76624 -81703 -76616 -81659
rect -76524 -81703 -76516 -81659
rect -76424 -81703 -76416 -81659
rect -76324 -81703 -76316 -81659
rect -76224 -81703 -76216 -81659
rect -76124 -81703 -76116 -81659
rect -76024 -81703 -76016 -81659
rect -75924 -81703 -75916 -81659
rect -75824 -81703 -75816 -81659
rect -75724 -81703 -75716 -81659
rect -75624 -81703 -75616 -81659
rect -75524 -81703 -75516 -81659
rect -75424 -81703 -75416 -81659
rect -50017 -81661 -49973 -81653
rect -49917 -81661 -49873 -81653
rect -49817 -81661 -49773 -81653
rect -49717 -81661 -49673 -81653
rect -49617 -81661 -49573 -81653
rect -49517 -81661 -49473 -81653
rect -49417 -81661 -49373 -81653
rect -49317 -81661 -49273 -81653
rect -49217 -81661 -49173 -81653
rect -49117 -81661 -49073 -81653
rect -49017 -81661 -48973 -81653
rect -48917 -81661 -48873 -81653
rect -48817 -81661 -48773 -81653
rect -48717 -81661 -48673 -81653
rect -48617 -81661 -48573 -81653
rect -48517 -81661 -48473 -81653
rect -48017 -81661 -47973 -81653
rect -47917 -81661 -47873 -81653
rect -47817 -81661 -47773 -81653
rect -47717 -81661 -47673 -81653
rect -47617 -81661 -47573 -81653
rect -47517 -81661 -47473 -81653
rect -47417 -81661 -47373 -81653
rect -47317 -81661 -47273 -81653
rect -47217 -81661 -47173 -81653
rect -47117 -81661 -47073 -81653
rect -47017 -81661 -46973 -81653
rect -46917 -81661 -46873 -81653
rect -46817 -81661 -46773 -81653
rect -46717 -81661 -46673 -81653
rect -46617 -81661 -46573 -81653
rect -46517 -81661 -46473 -81653
rect -46017 -81661 -45973 -81653
rect -45917 -81661 -45873 -81653
rect -45817 -81661 -45773 -81653
rect -45717 -81661 -45673 -81653
rect -45617 -81661 -45573 -81653
rect -45517 -81661 -45473 -81653
rect -45417 -81661 -45373 -81653
rect -45317 -81661 -45273 -81653
rect -45217 -81661 -45173 -81653
rect -45117 -81661 -45073 -81653
rect -45017 -81661 -44973 -81653
rect -44917 -81661 -44873 -81653
rect -44817 -81661 -44773 -81653
rect -44717 -81661 -44673 -81653
rect -44617 -81661 -44573 -81653
rect -44517 -81661 -44473 -81653
rect -44017 -81661 -43973 -81653
rect -43917 -81661 -43873 -81653
rect -43817 -81661 -43773 -81653
rect -43717 -81661 -43673 -81653
rect -43617 -81661 -43573 -81653
rect -43517 -81661 -43473 -81653
rect -43417 -81661 -43373 -81653
rect -43317 -81661 -43273 -81653
rect -43217 -81661 -43173 -81653
rect -43117 -81661 -43073 -81653
rect -43017 -81661 -42973 -81653
rect -42917 -81661 -42873 -81653
rect -42817 -81661 -42773 -81653
rect -42717 -81661 -42673 -81653
rect -42617 -81661 -42573 -81653
rect -42517 -81661 -42473 -81653
rect 80737 -81655 80781 -81647
rect 80837 -81655 80881 -81647
rect 80937 -81655 80981 -81647
rect 81037 -81655 81081 -81647
rect 81137 -81655 81181 -81647
rect 81237 -81655 81281 -81647
rect 81337 -81655 81381 -81647
rect 81437 -81655 81481 -81647
rect 81537 -81655 81581 -81647
rect 81637 -81655 81681 -81647
rect 81737 -81655 81781 -81647
rect 81837 -81655 81881 -81647
rect 81937 -81655 81981 -81647
rect 82037 -81655 82081 -81647
rect 82137 -81655 82181 -81647
rect 82237 -81655 82281 -81647
rect 82737 -81655 82781 -81647
rect 82837 -81655 82881 -81647
rect 82937 -81655 82981 -81647
rect 83037 -81655 83081 -81647
rect 83137 -81655 83181 -81647
rect 83237 -81655 83281 -81647
rect 83337 -81655 83381 -81647
rect 83437 -81655 83481 -81647
rect 83537 -81655 83581 -81647
rect 83637 -81655 83681 -81647
rect 83737 -81655 83781 -81647
rect 83837 -81655 83881 -81647
rect 83937 -81655 83981 -81647
rect 84037 -81655 84081 -81647
rect 84137 -81655 84181 -81647
rect 84237 -81655 84281 -81647
rect 84737 -81655 84781 -81647
rect 84837 -81655 84881 -81647
rect 84937 -81655 84981 -81647
rect 85037 -81655 85081 -81647
rect 85137 -81655 85181 -81647
rect 85237 -81655 85281 -81647
rect 85337 -81655 85381 -81647
rect 85437 -81655 85481 -81647
rect 85537 -81655 85581 -81647
rect 85637 -81655 85681 -81647
rect 85737 -81655 85781 -81647
rect 85837 -81655 85881 -81647
rect 85937 -81655 85981 -81647
rect 86037 -81655 86081 -81647
rect 86137 -81655 86181 -81647
rect 86237 -81655 86281 -81647
rect 86737 -81655 86781 -81647
rect 86837 -81655 86881 -81647
rect 86937 -81655 86981 -81647
rect 87037 -81655 87081 -81647
rect 87137 -81655 87181 -81647
rect 87237 -81655 87281 -81647
rect 87337 -81655 87381 -81647
rect 87437 -81655 87481 -81647
rect 87537 -81655 87581 -81647
rect 87637 -81655 87681 -81647
rect 87737 -81655 87781 -81647
rect 87837 -81655 87881 -81647
rect 87937 -81655 87981 -81647
rect 88037 -81655 88081 -81647
rect 88137 -81655 88181 -81647
rect 88237 -81655 88281 -81647
rect -49973 -81705 -49965 -81661
rect -49873 -81705 -49865 -81661
rect -49773 -81705 -49765 -81661
rect -49673 -81705 -49665 -81661
rect -49573 -81705 -49565 -81661
rect -49473 -81705 -49465 -81661
rect -49373 -81705 -49365 -81661
rect -49273 -81705 -49265 -81661
rect -49173 -81705 -49165 -81661
rect -49073 -81705 -49065 -81661
rect -48973 -81705 -48965 -81661
rect -48873 -81705 -48865 -81661
rect -48773 -81705 -48765 -81661
rect -48673 -81705 -48665 -81661
rect -48573 -81705 -48565 -81661
rect -48473 -81705 -48465 -81661
rect -47973 -81705 -47965 -81661
rect -47873 -81705 -47865 -81661
rect -47773 -81705 -47765 -81661
rect -47673 -81705 -47665 -81661
rect -47573 -81705 -47565 -81661
rect -47473 -81705 -47465 -81661
rect -47373 -81705 -47365 -81661
rect -47273 -81705 -47265 -81661
rect -47173 -81705 -47165 -81661
rect -47073 -81705 -47065 -81661
rect -46973 -81705 -46965 -81661
rect -46873 -81705 -46865 -81661
rect -46773 -81705 -46765 -81661
rect -46673 -81705 -46665 -81661
rect -46573 -81705 -46565 -81661
rect -46473 -81705 -46465 -81661
rect -45973 -81705 -45965 -81661
rect -45873 -81705 -45865 -81661
rect -45773 -81705 -45765 -81661
rect -45673 -81705 -45665 -81661
rect -45573 -81705 -45565 -81661
rect -45473 -81705 -45465 -81661
rect -45373 -81705 -45365 -81661
rect -45273 -81705 -45265 -81661
rect -45173 -81705 -45165 -81661
rect -45073 -81705 -45065 -81661
rect -44973 -81705 -44965 -81661
rect -44873 -81705 -44865 -81661
rect -44773 -81705 -44765 -81661
rect -44673 -81705 -44665 -81661
rect -44573 -81705 -44565 -81661
rect -44473 -81705 -44465 -81661
rect -43973 -81705 -43965 -81661
rect -43873 -81705 -43865 -81661
rect -43773 -81705 -43765 -81661
rect -43673 -81705 -43665 -81661
rect -43573 -81705 -43565 -81661
rect -43473 -81705 -43465 -81661
rect -43373 -81705 -43365 -81661
rect -43273 -81705 -43265 -81661
rect -43173 -81705 -43165 -81661
rect -43073 -81705 -43065 -81661
rect -42973 -81705 -42965 -81661
rect -42873 -81705 -42865 -81661
rect -42773 -81705 -42765 -81661
rect -42673 -81705 -42665 -81661
rect -42573 -81705 -42565 -81661
rect -42473 -81705 -42465 -81661
rect 80781 -81699 80789 -81655
rect 80881 -81699 80889 -81655
rect 80981 -81699 80989 -81655
rect 81081 -81699 81089 -81655
rect 81181 -81699 81189 -81655
rect 81281 -81699 81289 -81655
rect 81381 -81699 81389 -81655
rect 81481 -81699 81489 -81655
rect 81581 -81699 81589 -81655
rect 81681 -81699 81689 -81655
rect 81781 -81699 81789 -81655
rect 81881 -81699 81889 -81655
rect 81981 -81699 81989 -81655
rect 82081 -81699 82089 -81655
rect 82181 -81699 82189 -81655
rect 82281 -81699 82289 -81655
rect 82781 -81699 82789 -81655
rect 82881 -81699 82889 -81655
rect 82981 -81699 82989 -81655
rect 83081 -81699 83089 -81655
rect 83181 -81699 83189 -81655
rect 83281 -81699 83289 -81655
rect 83381 -81699 83389 -81655
rect 83481 -81699 83489 -81655
rect 83581 -81699 83589 -81655
rect 83681 -81699 83689 -81655
rect 83781 -81699 83789 -81655
rect 83881 -81699 83889 -81655
rect 83981 -81699 83989 -81655
rect 84081 -81699 84089 -81655
rect 84181 -81699 84189 -81655
rect 84281 -81699 84289 -81655
rect 84781 -81699 84789 -81655
rect 84881 -81699 84889 -81655
rect 84981 -81699 84989 -81655
rect 85081 -81699 85089 -81655
rect 85181 -81699 85189 -81655
rect 85281 -81699 85289 -81655
rect 85381 -81699 85389 -81655
rect 85481 -81699 85489 -81655
rect 85581 -81699 85589 -81655
rect 85681 -81699 85689 -81655
rect 85781 -81699 85789 -81655
rect 85881 -81699 85889 -81655
rect 85981 -81699 85989 -81655
rect 86081 -81699 86089 -81655
rect 86181 -81699 86189 -81655
rect 86281 -81699 86289 -81655
rect 86781 -81699 86789 -81655
rect 86881 -81699 86889 -81655
rect 86981 -81699 86989 -81655
rect 87081 -81699 87089 -81655
rect 87181 -81699 87189 -81655
rect 87281 -81699 87289 -81655
rect 87381 -81699 87389 -81655
rect 87481 -81699 87489 -81655
rect 87581 -81699 87589 -81655
rect 87681 -81699 87689 -81655
rect 87781 -81699 87789 -81655
rect 87881 -81699 87889 -81655
rect 87981 -81699 87989 -81655
rect 88081 -81699 88089 -81655
rect 88181 -81699 88189 -81655
rect 88281 -81699 88289 -81655
rect -82968 -81759 -82924 -81751
rect -82868 -81759 -82824 -81751
rect -82768 -81759 -82724 -81751
rect -82668 -81759 -82624 -81751
rect -82568 -81759 -82524 -81751
rect -82468 -81759 -82424 -81751
rect -82368 -81759 -82324 -81751
rect -82268 -81759 -82224 -81751
rect -82168 -81759 -82124 -81751
rect -82068 -81759 -82024 -81751
rect -81968 -81759 -81924 -81751
rect -81868 -81759 -81824 -81751
rect -81768 -81759 -81724 -81751
rect -81668 -81759 -81624 -81751
rect -81568 -81759 -81524 -81751
rect -81468 -81759 -81424 -81751
rect -80968 -81759 -80924 -81751
rect -80868 -81759 -80824 -81751
rect -80768 -81759 -80724 -81751
rect -80668 -81759 -80624 -81751
rect -80568 -81759 -80524 -81751
rect -80468 -81759 -80424 -81751
rect -80368 -81759 -80324 -81751
rect -80268 -81759 -80224 -81751
rect -80168 -81759 -80124 -81751
rect -80068 -81759 -80024 -81751
rect -79968 -81759 -79924 -81751
rect -79868 -81759 -79824 -81751
rect -79768 -81759 -79724 -81751
rect -79668 -81759 -79624 -81751
rect -79568 -81759 -79524 -81751
rect -79468 -81759 -79424 -81751
rect -78968 -81759 -78924 -81751
rect -78868 -81759 -78824 -81751
rect -78768 -81759 -78724 -81751
rect -78668 -81759 -78624 -81751
rect -78568 -81759 -78524 -81751
rect -78468 -81759 -78424 -81751
rect -78368 -81759 -78324 -81751
rect -78268 -81759 -78224 -81751
rect -78168 -81759 -78124 -81751
rect -78068 -81759 -78024 -81751
rect -77968 -81759 -77924 -81751
rect -77868 -81759 -77824 -81751
rect -77768 -81759 -77724 -81751
rect -77668 -81759 -77624 -81751
rect -77568 -81759 -77524 -81751
rect -77468 -81759 -77424 -81751
rect -76968 -81759 -76924 -81751
rect -76868 -81759 -76824 -81751
rect -76768 -81759 -76724 -81751
rect -76668 -81759 -76624 -81751
rect -76568 -81759 -76524 -81751
rect -76468 -81759 -76424 -81751
rect -76368 -81759 -76324 -81751
rect -76268 -81759 -76224 -81751
rect -76168 -81759 -76124 -81751
rect -76068 -81759 -76024 -81751
rect -75968 -81759 -75924 -81751
rect -75868 -81759 -75824 -81751
rect -75768 -81759 -75724 -81751
rect -75668 -81759 -75624 -81751
rect -75568 -81759 -75524 -81751
rect -75468 -81759 -75424 -81751
rect -82924 -81803 -82916 -81759
rect -82824 -81803 -82816 -81759
rect -82724 -81803 -82716 -81759
rect -82624 -81803 -82616 -81759
rect -82524 -81803 -82516 -81759
rect -82424 -81803 -82416 -81759
rect -82324 -81803 -82316 -81759
rect -82224 -81803 -82216 -81759
rect -82124 -81803 -82116 -81759
rect -82024 -81803 -82016 -81759
rect -81924 -81803 -81916 -81759
rect -81824 -81803 -81816 -81759
rect -81724 -81803 -81716 -81759
rect -81624 -81803 -81616 -81759
rect -81524 -81803 -81516 -81759
rect -81424 -81803 -81416 -81759
rect -80924 -81803 -80916 -81759
rect -80824 -81803 -80816 -81759
rect -80724 -81803 -80716 -81759
rect -80624 -81803 -80616 -81759
rect -80524 -81803 -80516 -81759
rect -80424 -81803 -80416 -81759
rect -80324 -81803 -80316 -81759
rect -80224 -81803 -80216 -81759
rect -80124 -81803 -80116 -81759
rect -80024 -81803 -80016 -81759
rect -79924 -81803 -79916 -81759
rect -79824 -81803 -79816 -81759
rect -79724 -81803 -79716 -81759
rect -79624 -81803 -79616 -81759
rect -79524 -81803 -79516 -81759
rect -79424 -81803 -79416 -81759
rect -78924 -81803 -78916 -81759
rect -78824 -81803 -78816 -81759
rect -78724 -81803 -78716 -81759
rect -78624 -81803 -78616 -81759
rect -78524 -81803 -78516 -81759
rect -78424 -81803 -78416 -81759
rect -78324 -81803 -78316 -81759
rect -78224 -81803 -78216 -81759
rect -78124 -81803 -78116 -81759
rect -78024 -81803 -78016 -81759
rect -77924 -81803 -77916 -81759
rect -77824 -81803 -77816 -81759
rect -77724 -81803 -77716 -81759
rect -77624 -81803 -77616 -81759
rect -77524 -81803 -77516 -81759
rect -77424 -81803 -77416 -81759
rect -76924 -81803 -76916 -81759
rect -76824 -81803 -76816 -81759
rect -76724 -81803 -76716 -81759
rect -76624 -81803 -76616 -81759
rect -76524 -81803 -76516 -81759
rect -76424 -81803 -76416 -81759
rect -76324 -81803 -76316 -81759
rect -76224 -81803 -76216 -81759
rect -76124 -81803 -76116 -81759
rect -76024 -81803 -76016 -81759
rect -75924 -81803 -75916 -81759
rect -75824 -81803 -75816 -81759
rect -75724 -81803 -75716 -81759
rect -75624 -81803 -75616 -81759
rect -75524 -81803 -75516 -81759
rect -75424 -81803 -75416 -81759
rect -50017 -81761 -49973 -81753
rect -49917 -81761 -49873 -81753
rect -49817 -81761 -49773 -81753
rect -49717 -81761 -49673 -81753
rect -49617 -81761 -49573 -81753
rect -49517 -81761 -49473 -81753
rect -49417 -81761 -49373 -81753
rect -49317 -81761 -49273 -81753
rect -49217 -81761 -49173 -81753
rect -49117 -81761 -49073 -81753
rect -49017 -81761 -48973 -81753
rect -48917 -81761 -48873 -81753
rect -48817 -81761 -48773 -81753
rect -48717 -81761 -48673 -81753
rect -48617 -81761 -48573 -81753
rect -48517 -81761 -48473 -81753
rect -48017 -81761 -47973 -81753
rect -47917 -81761 -47873 -81753
rect -47817 -81761 -47773 -81753
rect -47717 -81761 -47673 -81753
rect -47617 -81761 -47573 -81753
rect -47517 -81761 -47473 -81753
rect -47417 -81761 -47373 -81753
rect -47317 -81761 -47273 -81753
rect -47217 -81761 -47173 -81753
rect -47117 -81761 -47073 -81753
rect -47017 -81761 -46973 -81753
rect -46917 -81761 -46873 -81753
rect -46817 -81761 -46773 -81753
rect -46717 -81761 -46673 -81753
rect -46617 -81761 -46573 -81753
rect -46517 -81761 -46473 -81753
rect -46017 -81761 -45973 -81753
rect -45917 -81761 -45873 -81753
rect -45817 -81761 -45773 -81753
rect -45717 -81761 -45673 -81753
rect -45617 -81761 -45573 -81753
rect -45517 -81761 -45473 -81753
rect -45417 -81761 -45373 -81753
rect -45317 -81761 -45273 -81753
rect -45217 -81761 -45173 -81753
rect -45117 -81761 -45073 -81753
rect -45017 -81761 -44973 -81753
rect -44917 -81761 -44873 -81753
rect -44817 -81761 -44773 -81753
rect -44717 -81761 -44673 -81753
rect -44617 -81761 -44573 -81753
rect -44517 -81761 -44473 -81753
rect -44017 -81761 -43973 -81753
rect -43917 -81761 -43873 -81753
rect -43817 -81761 -43773 -81753
rect -43717 -81761 -43673 -81753
rect -43617 -81761 -43573 -81753
rect -43517 -81761 -43473 -81753
rect -43417 -81761 -43373 -81753
rect -43317 -81761 -43273 -81753
rect -43217 -81761 -43173 -81753
rect -43117 -81761 -43073 -81753
rect -43017 -81761 -42973 -81753
rect -42917 -81761 -42873 -81753
rect -42817 -81761 -42773 -81753
rect -42717 -81761 -42673 -81753
rect -42617 -81761 -42573 -81753
rect -42517 -81761 -42473 -81753
rect 80737 -81755 80781 -81747
rect 80837 -81755 80881 -81747
rect 80937 -81755 80981 -81747
rect 81037 -81755 81081 -81747
rect 81137 -81755 81181 -81747
rect 81237 -81755 81281 -81747
rect 81337 -81755 81381 -81747
rect 81437 -81755 81481 -81747
rect 81537 -81755 81581 -81747
rect 81637 -81755 81681 -81747
rect 81737 -81755 81781 -81747
rect 81837 -81755 81881 -81747
rect 81937 -81755 81981 -81747
rect 82037 -81755 82081 -81747
rect 82137 -81755 82181 -81747
rect 82237 -81755 82281 -81747
rect 82737 -81755 82781 -81747
rect 82837 -81755 82881 -81747
rect 82937 -81755 82981 -81747
rect 83037 -81755 83081 -81747
rect 83137 -81755 83181 -81747
rect 83237 -81755 83281 -81747
rect 83337 -81755 83381 -81747
rect 83437 -81755 83481 -81747
rect 83537 -81755 83581 -81747
rect 83637 -81755 83681 -81747
rect 83737 -81755 83781 -81747
rect 83837 -81755 83881 -81747
rect 83937 -81755 83981 -81747
rect 84037 -81755 84081 -81747
rect 84137 -81755 84181 -81747
rect 84237 -81755 84281 -81747
rect 84737 -81755 84781 -81747
rect 84837 -81755 84881 -81747
rect 84937 -81755 84981 -81747
rect 85037 -81755 85081 -81747
rect 85137 -81755 85181 -81747
rect 85237 -81755 85281 -81747
rect 85337 -81755 85381 -81747
rect 85437 -81755 85481 -81747
rect 85537 -81755 85581 -81747
rect 85637 -81755 85681 -81747
rect 85737 -81755 85781 -81747
rect 85837 -81755 85881 -81747
rect 85937 -81755 85981 -81747
rect 86037 -81755 86081 -81747
rect 86137 -81755 86181 -81747
rect 86237 -81755 86281 -81747
rect 86737 -81755 86781 -81747
rect 86837 -81755 86881 -81747
rect 86937 -81755 86981 -81747
rect 87037 -81755 87081 -81747
rect 87137 -81755 87181 -81747
rect 87237 -81755 87281 -81747
rect 87337 -81755 87381 -81747
rect 87437 -81755 87481 -81747
rect 87537 -81755 87581 -81747
rect 87637 -81755 87681 -81747
rect 87737 -81755 87781 -81747
rect 87837 -81755 87881 -81747
rect 87937 -81755 87981 -81747
rect 88037 -81755 88081 -81747
rect 88137 -81755 88181 -81747
rect 88237 -81755 88281 -81747
rect -49973 -81805 -49965 -81761
rect -49873 -81805 -49865 -81761
rect -49773 -81805 -49765 -81761
rect -49673 -81805 -49665 -81761
rect -49573 -81805 -49565 -81761
rect -49473 -81805 -49465 -81761
rect -49373 -81805 -49365 -81761
rect -49273 -81805 -49265 -81761
rect -49173 -81805 -49165 -81761
rect -49073 -81805 -49065 -81761
rect -48973 -81805 -48965 -81761
rect -48873 -81805 -48865 -81761
rect -48773 -81805 -48765 -81761
rect -48673 -81805 -48665 -81761
rect -48573 -81805 -48565 -81761
rect -48473 -81805 -48465 -81761
rect -47973 -81805 -47965 -81761
rect -47873 -81805 -47865 -81761
rect -47773 -81805 -47765 -81761
rect -47673 -81805 -47665 -81761
rect -47573 -81805 -47565 -81761
rect -47473 -81805 -47465 -81761
rect -47373 -81805 -47365 -81761
rect -47273 -81805 -47265 -81761
rect -47173 -81805 -47165 -81761
rect -47073 -81805 -47065 -81761
rect -46973 -81805 -46965 -81761
rect -46873 -81805 -46865 -81761
rect -46773 -81805 -46765 -81761
rect -46673 -81805 -46665 -81761
rect -46573 -81805 -46565 -81761
rect -46473 -81805 -46465 -81761
rect -45973 -81805 -45965 -81761
rect -45873 -81805 -45865 -81761
rect -45773 -81805 -45765 -81761
rect -45673 -81805 -45665 -81761
rect -45573 -81805 -45565 -81761
rect -45473 -81805 -45465 -81761
rect -45373 -81805 -45365 -81761
rect -45273 -81805 -45265 -81761
rect -45173 -81805 -45165 -81761
rect -45073 -81805 -45065 -81761
rect -44973 -81805 -44965 -81761
rect -44873 -81805 -44865 -81761
rect -44773 -81805 -44765 -81761
rect -44673 -81805 -44665 -81761
rect -44573 -81805 -44565 -81761
rect -44473 -81805 -44465 -81761
rect -43973 -81805 -43965 -81761
rect -43873 -81805 -43865 -81761
rect -43773 -81805 -43765 -81761
rect -43673 -81805 -43665 -81761
rect -43573 -81805 -43565 -81761
rect -43473 -81805 -43465 -81761
rect -43373 -81805 -43365 -81761
rect -43273 -81805 -43265 -81761
rect -43173 -81805 -43165 -81761
rect -43073 -81805 -43065 -81761
rect -42973 -81805 -42965 -81761
rect -42873 -81805 -42865 -81761
rect -42773 -81805 -42765 -81761
rect -42673 -81805 -42665 -81761
rect -42573 -81805 -42565 -81761
rect -42473 -81805 -42465 -81761
rect 80781 -81799 80789 -81755
rect 80881 -81799 80889 -81755
rect 80981 -81799 80989 -81755
rect 81081 -81799 81089 -81755
rect 81181 -81799 81189 -81755
rect 81281 -81799 81289 -81755
rect 81381 -81799 81389 -81755
rect 81481 -81799 81489 -81755
rect 81581 -81799 81589 -81755
rect 81681 -81799 81689 -81755
rect 81781 -81799 81789 -81755
rect 81881 -81799 81889 -81755
rect 81981 -81799 81989 -81755
rect 82081 -81799 82089 -81755
rect 82181 -81799 82189 -81755
rect 82281 -81799 82289 -81755
rect 82781 -81799 82789 -81755
rect 82881 -81799 82889 -81755
rect 82981 -81799 82989 -81755
rect 83081 -81799 83089 -81755
rect 83181 -81799 83189 -81755
rect 83281 -81799 83289 -81755
rect 83381 -81799 83389 -81755
rect 83481 -81799 83489 -81755
rect 83581 -81799 83589 -81755
rect 83681 -81799 83689 -81755
rect 83781 -81799 83789 -81755
rect 83881 -81799 83889 -81755
rect 83981 -81799 83989 -81755
rect 84081 -81799 84089 -81755
rect 84181 -81799 84189 -81755
rect 84281 -81799 84289 -81755
rect 84781 -81799 84789 -81755
rect 84881 -81799 84889 -81755
rect 84981 -81799 84989 -81755
rect 85081 -81799 85089 -81755
rect 85181 -81799 85189 -81755
rect 85281 -81799 85289 -81755
rect 85381 -81799 85389 -81755
rect 85481 -81799 85489 -81755
rect 85581 -81799 85589 -81755
rect 85681 -81799 85689 -81755
rect 85781 -81799 85789 -81755
rect 85881 -81799 85889 -81755
rect 85981 -81799 85989 -81755
rect 86081 -81799 86089 -81755
rect 86181 -81799 86189 -81755
rect 86281 -81799 86289 -81755
rect 86781 -81799 86789 -81755
rect 86881 -81799 86889 -81755
rect 86981 -81799 86989 -81755
rect 87081 -81799 87089 -81755
rect 87181 -81799 87189 -81755
rect 87281 -81799 87289 -81755
rect 87381 -81799 87389 -81755
rect 87481 -81799 87489 -81755
rect 87581 -81799 87589 -81755
rect 87681 -81799 87689 -81755
rect 87781 -81799 87789 -81755
rect 87881 -81799 87889 -81755
rect 87981 -81799 87989 -81755
rect 88081 -81799 88089 -81755
rect 88181 -81799 88189 -81755
rect 88281 -81799 88289 -81755
rect -82968 -81859 -82924 -81851
rect -82868 -81859 -82824 -81851
rect -82768 -81859 -82724 -81851
rect -82668 -81859 -82624 -81851
rect -82568 -81859 -82524 -81851
rect -82468 -81859 -82424 -81851
rect -82368 -81859 -82324 -81851
rect -82268 -81859 -82224 -81851
rect -82168 -81859 -82124 -81851
rect -82068 -81859 -82024 -81851
rect -81968 -81859 -81924 -81851
rect -81868 -81859 -81824 -81851
rect -81768 -81859 -81724 -81851
rect -81668 -81859 -81624 -81851
rect -81568 -81859 -81524 -81851
rect -81468 -81859 -81424 -81851
rect -80968 -81859 -80924 -81851
rect -80868 -81859 -80824 -81851
rect -80768 -81859 -80724 -81851
rect -80668 -81859 -80624 -81851
rect -80568 -81859 -80524 -81851
rect -80468 -81859 -80424 -81851
rect -80368 -81859 -80324 -81851
rect -80268 -81859 -80224 -81851
rect -80168 -81859 -80124 -81851
rect -80068 -81859 -80024 -81851
rect -79968 -81859 -79924 -81851
rect -79868 -81859 -79824 -81851
rect -79768 -81859 -79724 -81851
rect -79668 -81859 -79624 -81851
rect -79568 -81859 -79524 -81851
rect -79468 -81859 -79424 -81851
rect -78968 -81859 -78924 -81851
rect -78868 -81859 -78824 -81851
rect -78768 -81859 -78724 -81851
rect -78668 -81859 -78624 -81851
rect -78568 -81859 -78524 -81851
rect -78468 -81859 -78424 -81851
rect -78368 -81859 -78324 -81851
rect -78268 -81859 -78224 -81851
rect -78168 -81859 -78124 -81851
rect -78068 -81859 -78024 -81851
rect -77968 -81859 -77924 -81851
rect -77868 -81859 -77824 -81851
rect -77768 -81859 -77724 -81851
rect -77668 -81859 -77624 -81851
rect -77568 -81859 -77524 -81851
rect -77468 -81859 -77424 -81851
rect -76968 -81859 -76924 -81851
rect -76868 -81859 -76824 -81851
rect -76768 -81859 -76724 -81851
rect -76668 -81859 -76624 -81851
rect -76568 -81859 -76524 -81851
rect -76468 -81859 -76424 -81851
rect -76368 -81859 -76324 -81851
rect -76268 -81859 -76224 -81851
rect -76168 -81859 -76124 -81851
rect -76068 -81859 -76024 -81851
rect -75968 -81859 -75924 -81851
rect -75868 -81859 -75824 -81851
rect -75768 -81859 -75724 -81851
rect -75668 -81859 -75624 -81851
rect -75568 -81859 -75524 -81851
rect -75468 -81859 -75424 -81851
rect -82924 -81903 -82916 -81859
rect -82824 -81903 -82816 -81859
rect -82724 -81903 -82716 -81859
rect -82624 -81903 -82616 -81859
rect -82524 -81903 -82516 -81859
rect -82424 -81903 -82416 -81859
rect -82324 -81903 -82316 -81859
rect -82224 -81903 -82216 -81859
rect -82124 -81903 -82116 -81859
rect -82024 -81903 -82016 -81859
rect -81924 -81903 -81916 -81859
rect -81824 -81903 -81816 -81859
rect -81724 -81903 -81716 -81859
rect -81624 -81903 -81616 -81859
rect -81524 -81903 -81516 -81859
rect -81424 -81903 -81416 -81859
rect -80924 -81903 -80916 -81859
rect -80824 -81903 -80816 -81859
rect -80724 -81903 -80716 -81859
rect -80624 -81903 -80616 -81859
rect -80524 -81903 -80516 -81859
rect -80424 -81903 -80416 -81859
rect -80324 -81903 -80316 -81859
rect -80224 -81903 -80216 -81859
rect -80124 -81903 -80116 -81859
rect -80024 -81903 -80016 -81859
rect -79924 -81903 -79916 -81859
rect -79824 -81903 -79816 -81859
rect -79724 -81903 -79716 -81859
rect -79624 -81903 -79616 -81859
rect -79524 -81903 -79516 -81859
rect -79424 -81903 -79416 -81859
rect -78924 -81903 -78916 -81859
rect -78824 -81903 -78816 -81859
rect -78724 -81903 -78716 -81859
rect -78624 -81903 -78616 -81859
rect -78524 -81903 -78516 -81859
rect -78424 -81903 -78416 -81859
rect -78324 -81903 -78316 -81859
rect -78224 -81903 -78216 -81859
rect -78124 -81903 -78116 -81859
rect -78024 -81903 -78016 -81859
rect -77924 -81903 -77916 -81859
rect -77824 -81903 -77816 -81859
rect -77724 -81903 -77716 -81859
rect -77624 -81903 -77616 -81859
rect -77524 -81903 -77516 -81859
rect -77424 -81903 -77416 -81859
rect -76924 -81903 -76916 -81859
rect -76824 -81903 -76816 -81859
rect -76724 -81903 -76716 -81859
rect -76624 -81903 -76616 -81859
rect -76524 -81903 -76516 -81859
rect -76424 -81903 -76416 -81859
rect -76324 -81903 -76316 -81859
rect -76224 -81903 -76216 -81859
rect -76124 -81903 -76116 -81859
rect -76024 -81903 -76016 -81859
rect -75924 -81903 -75916 -81859
rect -75824 -81903 -75816 -81859
rect -75724 -81903 -75716 -81859
rect -75624 -81903 -75616 -81859
rect -75524 -81903 -75516 -81859
rect -75424 -81903 -75416 -81859
rect -50017 -81861 -49973 -81853
rect -49917 -81861 -49873 -81853
rect -49817 -81861 -49773 -81853
rect -49717 -81861 -49673 -81853
rect -49617 -81861 -49573 -81853
rect -49517 -81861 -49473 -81853
rect -49417 -81861 -49373 -81853
rect -49317 -81861 -49273 -81853
rect -49217 -81861 -49173 -81853
rect -49117 -81861 -49073 -81853
rect -49017 -81861 -48973 -81853
rect -48917 -81861 -48873 -81853
rect -48817 -81861 -48773 -81853
rect -48717 -81861 -48673 -81853
rect -48617 -81861 -48573 -81853
rect -48517 -81861 -48473 -81853
rect -48017 -81861 -47973 -81853
rect -47917 -81861 -47873 -81853
rect -47817 -81861 -47773 -81853
rect -47717 -81861 -47673 -81853
rect -47617 -81861 -47573 -81853
rect -47517 -81861 -47473 -81853
rect -47417 -81861 -47373 -81853
rect -47317 -81861 -47273 -81853
rect -47217 -81861 -47173 -81853
rect -47117 -81861 -47073 -81853
rect -47017 -81861 -46973 -81853
rect -46917 -81861 -46873 -81853
rect -46817 -81861 -46773 -81853
rect -46717 -81861 -46673 -81853
rect -46617 -81861 -46573 -81853
rect -46517 -81861 -46473 -81853
rect -46017 -81861 -45973 -81853
rect -45917 -81861 -45873 -81853
rect -45817 -81861 -45773 -81853
rect -45717 -81861 -45673 -81853
rect -45617 -81861 -45573 -81853
rect -45517 -81861 -45473 -81853
rect -45417 -81861 -45373 -81853
rect -45317 -81861 -45273 -81853
rect -45217 -81861 -45173 -81853
rect -45117 -81861 -45073 -81853
rect -45017 -81861 -44973 -81853
rect -44917 -81861 -44873 -81853
rect -44817 -81861 -44773 -81853
rect -44717 -81861 -44673 -81853
rect -44617 -81861 -44573 -81853
rect -44517 -81861 -44473 -81853
rect -44017 -81861 -43973 -81853
rect -43917 -81861 -43873 -81853
rect -43817 -81861 -43773 -81853
rect -43717 -81861 -43673 -81853
rect -43617 -81861 -43573 -81853
rect -43517 -81861 -43473 -81853
rect -43417 -81861 -43373 -81853
rect -43317 -81861 -43273 -81853
rect -43217 -81861 -43173 -81853
rect -43117 -81861 -43073 -81853
rect -43017 -81861 -42973 -81853
rect -42917 -81861 -42873 -81853
rect -42817 -81861 -42773 -81853
rect -42717 -81861 -42673 -81853
rect -42617 -81861 -42573 -81853
rect -42517 -81861 -42473 -81853
rect 80737 -81855 80781 -81847
rect 80837 -81855 80881 -81847
rect 80937 -81855 80981 -81847
rect 81037 -81855 81081 -81847
rect 81137 -81855 81181 -81847
rect 81237 -81855 81281 -81847
rect 81337 -81855 81381 -81847
rect 81437 -81855 81481 -81847
rect 81537 -81855 81581 -81847
rect 81637 -81855 81681 -81847
rect 81737 -81855 81781 -81847
rect 81837 -81855 81881 -81847
rect 81937 -81855 81981 -81847
rect 82037 -81855 82081 -81847
rect 82137 -81855 82181 -81847
rect 82237 -81855 82281 -81847
rect 82737 -81855 82781 -81847
rect 82837 -81855 82881 -81847
rect 82937 -81855 82981 -81847
rect 83037 -81855 83081 -81847
rect 83137 -81855 83181 -81847
rect 83237 -81855 83281 -81847
rect 83337 -81855 83381 -81847
rect 83437 -81855 83481 -81847
rect 83537 -81855 83581 -81847
rect 83637 -81855 83681 -81847
rect 83737 -81855 83781 -81847
rect 83837 -81855 83881 -81847
rect 83937 -81855 83981 -81847
rect 84037 -81855 84081 -81847
rect 84137 -81855 84181 -81847
rect 84237 -81855 84281 -81847
rect 84737 -81855 84781 -81847
rect 84837 -81855 84881 -81847
rect 84937 -81855 84981 -81847
rect 85037 -81855 85081 -81847
rect 85137 -81855 85181 -81847
rect 85237 -81855 85281 -81847
rect 85337 -81855 85381 -81847
rect 85437 -81855 85481 -81847
rect 85537 -81855 85581 -81847
rect 85637 -81855 85681 -81847
rect 85737 -81855 85781 -81847
rect 85837 -81855 85881 -81847
rect 85937 -81855 85981 -81847
rect 86037 -81855 86081 -81847
rect 86137 -81855 86181 -81847
rect 86237 -81855 86281 -81847
rect 86737 -81855 86781 -81847
rect 86837 -81855 86881 -81847
rect 86937 -81855 86981 -81847
rect 87037 -81855 87081 -81847
rect 87137 -81855 87181 -81847
rect 87237 -81855 87281 -81847
rect 87337 -81855 87381 -81847
rect 87437 -81855 87481 -81847
rect 87537 -81855 87581 -81847
rect 87637 -81855 87681 -81847
rect 87737 -81855 87781 -81847
rect 87837 -81855 87881 -81847
rect 87937 -81855 87981 -81847
rect 88037 -81855 88081 -81847
rect 88137 -81855 88181 -81847
rect 88237 -81855 88281 -81847
rect -49973 -81905 -49965 -81861
rect -49873 -81905 -49865 -81861
rect -49773 -81905 -49765 -81861
rect -49673 -81905 -49665 -81861
rect -49573 -81905 -49565 -81861
rect -49473 -81905 -49465 -81861
rect -49373 -81905 -49365 -81861
rect -49273 -81905 -49265 -81861
rect -49173 -81905 -49165 -81861
rect -49073 -81905 -49065 -81861
rect -48973 -81905 -48965 -81861
rect -48873 -81905 -48865 -81861
rect -48773 -81905 -48765 -81861
rect -48673 -81905 -48665 -81861
rect -48573 -81905 -48565 -81861
rect -48473 -81905 -48465 -81861
rect -47973 -81905 -47965 -81861
rect -47873 -81905 -47865 -81861
rect -47773 -81905 -47765 -81861
rect -47673 -81905 -47665 -81861
rect -47573 -81905 -47565 -81861
rect -47473 -81905 -47465 -81861
rect -47373 -81905 -47365 -81861
rect -47273 -81905 -47265 -81861
rect -47173 -81905 -47165 -81861
rect -47073 -81905 -47065 -81861
rect -46973 -81905 -46965 -81861
rect -46873 -81905 -46865 -81861
rect -46773 -81905 -46765 -81861
rect -46673 -81905 -46665 -81861
rect -46573 -81905 -46565 -81861
rect -46473 -81905 -46465 -81861
rect -45973 -81905 -45965 -81861
rect -45873 -81905 -45865 -81861
rect -45773 -81905 -45765 -81861
rect -45673 -81905 -45665 -81861
rect -45573 -81905 -45565 -81861
rect -45473 -81905 -45465 -81861
rect -45373 -81905 -45365 -81861
rect -45273 -81905 -45265 -81861
rect -45173 -81905 -45165 -81861
rect -45073 -81905 -45065 -81861
rect -44973 -81905 -44965 -81861
rect -44873 -81905 -44865 -81861
rect -44773 -81905 -44765 -81861
rect -44673 -81905 -44665 -81861
rect -44573 -81905 -44565 -81861
rect -44473 -81905 -44465 -81861
rect -43973 -81905 -43965 -81861
rect -43873 -81905 -43865 -81861
rect -43773 -81905 -43765 -81861
rect -43673 -81905 -43665 -81861
rect -43573 -81905 -43565 -81861
rect -43473 -81905 -43465 -81861
rect -43373 -81905 -43365 -81861
rect -43273 -81905 -43265 -81861
rect -43173 -81905 -43165 -81861
rect -43073 -81905 -43065 -81861
rect -42973 -81905 -42965 -81861
rect -42873 -81905 -42865 -81861
rect -42773 -81905 -42765 -81861
rect -42673 -81905 -42665 -81861
rect -42573 -81905 -42565 -81861
rect -42473 -81905 -42465 -81861
rect 80781 -81899 80789 -81855
rect 80881 -81899 80889 -81855
rect 80981 -81899 80989 -81855
rect 81081 -81899 81089 -81855
rect 81181 -81899 81189 -81855
rect 81281 -81899 81289 -81855
rect 81381 -81899 81389 -81855
rect 81481 -81899 81489 -81855
rect 81581 -81899 81589 -81855
rect 81681 -81899 81689 -81855
rect 81781 -81899 81789 -81855
rect 81881 -81899 81889 -81855
rect 81981 -81899 81989 -81855
rect 82081 -81899 82089 -81855
rect 82181 -81899 82189 -81855
rect 82281 -81899 82289 -81855
rect 82781 -81899 82789 -81855
rect 82881 -81899 82889 -81855
rect 82981 -81899 82989 -81855
rect 83081 -81899 83089 -81855
rect 83181 -81899 83189 -81855
rect 83281 -81899 83289 -81855
rect 83381 -81899 83389 -81855
rect 83481 -81899 83489 -81855
rect 83581 -81899 83589 -81855
rect 83681 -81899 83689 -81855
rect 83781 -81899 83789 -81855
rect 83881 -81899 83889 -81855
rect 83981 -81899 83989 -81855
rect 84081 -81899 84089 -81855
rect 84181 -81899 84189 -81855
rect 84281 -81899 84289 -81855
rect 84781 -81899 84789 -81855
rect 84881 -81899 84889 -81855
rect 84981 -81899 84989 -81855
rect 85081 -81899 85089 -81855
rect 85181 -81899 85189 -81855
rect 85281 -81899 85289 -81855
rect 85381 -81899 85389 -81855
rect 85481 -81899 85489 -81855
rect 85581 -81899 85589 -81855
rect 85681 -81899 85689 -81855
rect 85781 -81899 85789 -81855
rect 85881 -81899 85889 -81855
rect 85981 -81899 85989 -81855
rect 86081 -81899 86089 -81855
rect 86181 -81899 86189 -81855
rect 86281 -81899 86289 -81855
rect 86781 -81899 86789 -81855
rect 86881 -81899 86889 -81855
rect 86981 -81899 86989 -81855
rect 87081 -81899 87089 -81855
rect 87181 -81899 87189 -81855
rect 87281 -81899 87289 -81855
rect 87381 -81899 87389 -81855
rect 87481 -81899 87489 -81855
rect 87581 -81899 87589 -81855
rect 87681 -81899 87689 -81855
rect 87781 -81899 87789 -81855
rect 87881 -81899 87889 -81855
rect 87981 -81899 87989 -81855
rect 88081 -81899 88089 -81855
rect 88181 -81899 88189 -81855
rect 88281 -81899 88289 -81855
rect -82968 -81959 -82924 -81951
rect -82868 -81959 -82824 -81951
rect -82768 -81959 -82724 -81951
rect -82668 -81959 -82624 -81951
rect -82568 -81959 -82524 -81951
rect -82468 -81959 -82424 -81951
rect -82368 -81959 -82324 -81951
rect -82268 -81959 -82224 -81951
rect -82168 -81959 -82124 -81951
rect -82068 -81959 -82024 -81951
rect -81968 -81959 -81924 -81951
rect -81868 -81959 -81824 -81951
rect -81768 -81959 -81724 -81951
rect -81668 -81959 -81624 -81951
rect -81568 -81959 -81524 -81951
rect -81468 -81959 -81424 -81951
rect -80968 -81959 -80924 -81951
rect -80868 -81959 -80824 -81951
rect -80768 -81959 -80724 -81951
rect -80668 -81959 -80624 -81951
rect -80568 -81959 -80524 -81951
rect -80468 -81959 -80424 -81951
rect -80368 -81959 -80324 -81951
rect -80268 -81959 -80224 -81951
rect -80168 -81959 -80124 -81951
rect -80068 -81959 -80024 -81951
rect -79968 -81959 -79924 -81951
rect -79868 -81959 -79824 -81951
rect -79768 -81959 -79724 -81951
rect -79668 -81959 -79624 -81951
rect -79568 -81959 -79524 -81951
rect -79468 -81959 -79424 -81951
rect -78968 -81959 -78924 -81951
rect -78868 -81959 -78824 -81951
rect -78768 -81959 -78724 -81951
rect -78668 -81959 -78624 -81951
rect -78568 -81959 -78524 -81951
rect -78468 -81959 -78424 -81951
rect -78368 -81959 -78324 -81951
rect -78268 -81959 -78224 -81951
rect -78168 -81959 -78124 -81951
rect -78068 -81959 -78024 -81951
rect -77968 -81959 -77924 -81951
rect -77868 -81959 -77824 -81951
rect -77768 -81959 -77724 -81951
rect -77668 -81959 -77624 -81951
rect -77568 -81959 -77524 -81951
rect -77468 -81959 -77424 -81951
rect -76968 -81959 -76924 -81951
rect -76868 -81959 -76824 -81951
rect -76768 -81959 -76724 -81951
rect -76668 -81959 -76624 -81951
rect -76568 -81959 -76524 -81951
rect -76468 -81959 -76424 -81951
rect -76368 -81959 -76324 -81951
rect -76268 -81959 -76224 -81951
rect -76168 -81959 -76124 -81951
rect -76068 -81959 -76024 -81951
rect -75968 -81959 -75924 -81951
rect -75868 -81959 -75824 -81951
rect -75768 -81959 -75724 -81951
rect -75668 -81959 -75624 -81951
rect -75568 -81959 -75524 -81951
rect -75468 -81959 -75424 -81951
rect -82924 -82003 -82916 -81959
rect -82824 -82003 -82816 -81959
rect -82724 -82003 -82716 -81959
rect -82624 -82003 -82616 -81959
rect -82524 -82003 -82516 -81959
rect -82424 -82003 -82416 -81959
rect -82324 -82003 -82316 -81959
rect -82224 -82003 -82216 -81959
rect -82124 -82003 -82116 -81959
rect -82024 -82003 -82016 -81959
rect -81924 -82003 -81916 -81959
rect -81824 -82003 -81816 -81959
rect -81724 -82003 -81716 -81959
rect -81624 -82003 -81616 -81959
rect -81524 -82003 -81516 -81959
rect -81424 -82003 -81416 -81959
rect -80924 -82003 -80916 -81959
rect -80824 -82003 -80816 -81959
rect -80724 -82003 -80716 -81959
rect -80624 -82003 -80616 -81959
rect -80524 -82003 -80516 -81959
rect -80424 -82003 -80416 -81959
rect -80324 -82003 -80316 -81959
rect -80224 -82003 -80216 -81959
rect -80124 -82003 -80116 -81959
rect -80024 -82003 -80016 -81959
rect -79924 -82003 -79916 -81959
rect -79824 -82003 -79816 -81959
rect -79724 -82003 -79716 -81959
rect -79624 -82003 -79616 -81959
rect -79524 -82003 -79516 -81959
rect -79424 -82003 -79416 -81959
rect -78924 -82003 -78916 -81959
rect -78824 -82003 -78816 -81959
rect -78724 -82003 -78716 -81959
rect -78624 -82003 -78616 -81959
rect -78524 -82003 -78516 -81959
rect -78424 -82003 -78416 -81959
rect -78324 -82003 -78316 -81959
rect -78224 -82003 -78216 -81959
rect -78124 -82003 -78116 -81959
rect -78024 -82003 -78016 -81959
rect -77924 -82003 -77916 -81959
rect -77824 -82003 -77816 -81959
rect -77724 -82003 -77716 -81959
rect -77624 -82003 -77616 -81959
rect -77524 -82003 -77516 -81959
rect -77424 -82003 -77416 -81959
rect -76924 -82003 -76916 -81959
rect -76824 -82003 -76816 -81959
rect -76724 -82003 -76716 -81959
rect -76624 -82003 -76616 -81959
rect -76524 -82003 -76516 -81959
rect -76424 -82003 -76416 -81959
rect -76324 -82003 -76316 -81959
rect -76224 -82003 -76216 -81959
rect -76124 -82003 -76116 -81959
rect -76024 -82003 -76016 -81959
rect -75924 -82003 -75916 -81959
rect -75824 -82003 -75816 -81959
rect -75724 -82003 -75716 -81959
rect -75624 -82003 -75616 -81959
rect -75524 -82003 -75516 -81959
rect -75424 -82003 -75416 -81959
rect -50017 -81961 -49973 -81953
rect -49917 -81961 -49873 -81953
rect -49817 -81961 -49773 -81953
rect -49717 -81961 -49673 -81953
rect -49617 -81961 -49573 -81953
rect -49517 -81961 -49473 -81953
rect -49417 -81961 -49373 -81953
rect -49317 -81961 -49273 -81953
rect -49217 -81961 -49173 -81953
rect -49117 -81961 -49073 -81953
rect -49017 -81961 -48973 -81953
rect -48917 -81961 -48873 -81953
rect -48817 -81961 -48773 -81953
rect -48717 -81961 -48673 -81953
rect -48617 -81961 -48573 -81953
rect -48517 -81961 -48473 -81953
rect -48017 -81961 -47973 -81953
rect -47917 -81961 -47873 -81953
rect -47817 -81961 -47773 -81953
rect -47717 -81961 -47673 -81953
rect -47617 -81961 -47573 -81953
rect -47517 -81961 -47473 -81953
rect -47417 -81961 -47373 -81953
rect -47317 -81961 -47273 -81953
rect -47217 -81961 -47173 -81953
rect -47117 -81961 -47073 -81953
rect -47017 -81961 -46973 -81953
rect -46917 -81961 -46873 -81953
rect -46817 -81961 -46773 -81953
rect -46717 -81961 -46673 -81953
rect -46617 -81961 -46573 -81953
rect -46517 -81961 -46473 -81953
rect -46017 -81961 -45973 -81953
rect -45917 -81961 -45873 -81953
rect -45817 -81961 -45773 -81953
rect -45717 -81961 -45673 -81953
rect -45617 -81961 -45573 -81953
rect -45517 -81961 -45473 -81953
rect -45417 -81961 -45373 -81953
rect -45317 -81961 -45273 -81953
rect -45217 -81961 -45173 -81953
rect -45117 -81961 -45073 -81953
rect -45017 -81961 -44973 -81953
rect -44917 -81961 -44873 -81953
rect -44817 -81961 -44773 -81953
rect -44717 -81961 -44673 -81953
rect -44617 -81961 -44573 -81953
rect -44517 -81961 -44473 -81953
rect -44017 -81961 -43973 -81953
rect -43917 -81961 -43873 -81953
rect -43817 -81961 -43773 -81953
rect -43717 -81961 -43673 -81953
rect -43617 -81961 -43573 -81953
rect -43517 -81961 -43473 -81953
rect -43417 -81961 -43373 -81953
rect -43317 -81961 -43273 -81953
rect -43217 -81961 -43173 -81953
rect -43117 -81961 -43073 -81953
rect -43017 -81961 -42973 -81953
rect -42917 -81961 -42873 -81953
rect -42817 -81961 -42773 -81953
rect -42717 -81961 -42673 -81953
rect -42617 -81961 -42573 -81953
rect -42517 -81961 -42473 -81953
rect 80737 -81955 80781 -81947
rect 80837 -81955 80881 -81947
rect 80937 -81955 80981 -81947
rect 81037 -81955 81081 -81947
rect 81137 -81955 81181 -81947
rect 81237 -81955 81281 -81947
rect 81337 -81955 81381 -81947
rect 81437 -81955 81481 -81947
rect 81537 -81955 81581 -81947
rect 81637 -81955 81681 -81947
rect 81737 -81955 81781 -81947
rect 81837 -81955 81881 -81947
rect 81937 -81955 81981 -81947
rect 82037 -81955 82081 -81947
rect 82137 -81955 82181 -81947
rect 82237 -81955 82281 -81947
rect 82737 -81955 82781 -81947
rect 82837 -81955 82881 -81947
rect 82937 -81955 82981 -81947
rect 83037 -81955 83081 -81947
rect 83137 -81955 83181 -81947
rect 83237 -81955 83281 -81947
rect 83337 -81955 83381 -81947
rect 83437 -81955 83481 -81947
rect 83537 -81955 83581 -81947
rect 83637 -81955 83681 -81947
rect 83737 -81955 83781 -81947
rect 83837 -81955 83881 -81947
rect 83937 -81955 83981 -81947
rect 84037 -81955 84081 -81947
rect 84137 -81955 84181 -81947
rect 84237 -81955 84281 -81947
rect 84737 -81955 84781 -81947
rect 84837 -81955 84881 -81947
rect 84937 -81955 84981 -81947
rect 85037 -81955 85081 -81947
rect 85137 -81955 85181 -81947
rect 85237 -81955 85281 -81947
rect 85337 -81955 85381 -81947
rect 85437 -81955 85481 -81947
rect 85537 -81955 85581 -81947
rect 85637 -81955 85681 -81947
rect 85737 -81955 85781 -81947
rect 85837 -81955 85881 -81947
rect 85937 -81955 85981 -81947
rect 86037 -81955 86081 -81947
rect 86137 -81955 86181 -81947
rect 86237 -81955 86281 -81947
rect 86737 -81955 86781 -81947
rect 86837 -81955 86881 -81947
rect 86937 -81955 86981 -81947
rect 87037 -81955 87081 -81947
rect 87137 -81955 87181 -81947
rect 87237 -81955 87281 -81947
rect 87337 -81955 87381 -81947
rect 87437 -81955 87481 -81947
rect 87537 -81955 87581 -81947
rect 87637 -81955 87681 -81947
rect 87737 -81955 87781 -81947
rect 87837 -81955 87881 -81947
rect 87937 -81955 87981 -81947
rect 88037 -81955 88081 -81947
rect 88137 -81955 88181 -81947
rect 88237 -81955 88281 -81947
rect -49973 -82005 -49965 -81961
rect -49873 -82005 -49865 -81961
rect -49773 -82005 -49765 -81961
rect -49673 -82005 -49665 -81961
rect -49573 -82005 -49565 -81961
rect -49473 -82005 -49465 -81961
rect -49373 -82005 -49365 -81961
rect -49273 -82005 -49265 -81961
rect -49173 -82005 -49165 -81961
rect -49073 -82005 -49065 -81961
rect -48973 -82005 -48965 -81961
rect -48873 -82005 -48865 -81961
rect -48773 -82005 -48765 -81961
rect -48673 -82005 -48665 -81961
rect -48573 -82005 -48565 -81961
rect -48473 -82005 -48465 -81961
rect -47973 -82005 -47965 -81961
rect -47873 -82005 -47865 -81961
rect -47773 -82005 -47765 -81961
rect -47673 -82005 -47665 -81961
rect -47573 -82005 -47565 -81961
rect -47473 -82005 -47465 -81961
rect -47373 -82005 -47365 -81961
rect -47273 -82005 -47265 -81961
rect -47173 -82005 -47165 -81961
rect -47073 -82005 -47065 -81961
rect -46973 -82005 -46965 -81961
rect -46873 -82005 -46865 -81961
rect -46773 -82005 -46765 -81961
rect -46673 -82005 -46665 -81961
rect -46573 -82005 -46565 -81961
rect -46473 -82005 -46465 -81961
rect -45973 -82005 -45965 -81961
rect -45873 -82005 -45865 -81961
rect -45773 -82005 -45765 -81961
rect -45673 -82005 -45665 -81961
rect -45573 -82005 -45565 -81961
rect -45473 -82005 -45465 -81961
rect -45373 -82005 -45365 -81961
rect -45273 -82005 -45265 -81961
rect -45173 -82005 -45165 -81961
rect -45073 -82005 -45065 -81961
rect -44973 -82005 -44965 -81961
rect -44873 -82005 -44865 -81961
rect -44773 -82005 -44765 -81961
rect -44673 -82005 -44665 -81961
rect -44573 -82005 -44565 -81961
rect -44473 -82005 -44465 -81961
rect -43973 -82005 -43965 -81961
rect -43873 -82005 -43865 -81961
rect -43773 -82005 -43765 -81961
rect -43673 -82005 -43665 -81961
rect -43573 -82005 -43565 -81961
rect -43473 -82005 -43465 -81961
rect -43373 -82005 -43365 -81961
rect -43273 -82005 -43265 -81961
rect -43173 -82005 -43165 -81961
rect -43073 -82005 -43065 -81961
rect -42973 -82005 -42965 -81961
rect -42873 -82005 -42865 -81961
rect -42773 -82005 -42765 -81961
rect -42673 -82005 -42665 -81961
rect -42573 -82005 -42565 -81961
rect -42473 -82005 -42465 -81961
rect 80781 -81999 80789 -81955
rect 80881 -81999 80889 -81955
rect 80981 -81999 80989 -81955
rect 81081 -81999 81089 -81955
rect 81181 -81999 81189 -81955
rect 81281 -81999 81289 -81955
rect 81381 -81999 81389 -81955
rect 81481 -81999 81489 -81955
rect 81581 -81999 81589 -81955
rect 81681 -81999 81689 -81955
rect 81781 -81999 81789 -81955
rect 81881 -81999 81889 -81955
rect 81981 -81999 81989 -81955
rect 82081 -81999 82089 -81955
rect 82181 -81999 82189 -81955
rect 82281 -81999 82289 -81955
rect 82781 -81999 82789 -81955
rect 82881 -81999 82889 -81955
rect 82981 -81999 82989 -81955
rect 83081 -81999 83089 -81955
rect 83181 -81999 83189 -81955
rect 83281 -81999 83289 -81955
rect 83381 -81999 83389 -81955
rect 83481 -81999 83489 -81955
rect 83581 -81999 83589 -81955
rect 83681 -81999 83689 -81955
rect 83781 -81999 83789 -81955
rect 83881 -81999 83889 -81955
rect 83981 -81999 83989 -81955
rect 84081 -81999 84089 -81955
rect 84181 -81999 84189 -81955
rect 84281 -81999 84289 -81955
rect 84781 -81999 84789 -81955
rect 84881 -81999 84889 -81955
rect 84981 -81999 84989 -81955
rect 85081 -81999 85089 -81955
rect 85181 -81999 85189 -81955
rect 85281 -81999 85289 -81955
rect 85381 -81999 85389 -81955
rect 85481 -81999 85489 -81955
rect 85581 -81999 85589 -81955
rect 85681 -81999 85689 -81955
rect 85781 -81999 85789 -81955
rect 85881 -81999 85889 -81955
rect 85981 -81999 85989 -81955
rect 86081 -81999 86089 -81955
rect 86181 -81999 86189 -81955
rect 86281 -81999 86289 -81955
rect 86781 -81999 86789 -81955
rect 86881 -81999 86889 -81955
rect 86981 -81999 86989 -81955
rect 87081 -81999 87089 -81955
rect 87181 -81999 87189 -81955
rect 87281 -81999 87289 -81955
rect 87381 -81999 87389 -81955
rect 87481 -81999 87489 -81955
rect 87581 -81999 87589 -81955
rect 87681 -81999 87689 -81955
rect 87781 -81999 87789 -81955
rect 87881 -81999 87889 -81955
rect 87981 -81999 87989 -81955
rect 88081 -81999 88089 -81955
rect 88181 -81999 88189 -81955
rect 88281 -81999 88289 -81955
rect -109180 -103119 -109178 -83119
rect -109114 -103119 -109112 -83119
rect -77180 -103119 -77178 -83119
rect -77114 -103119 -77112 -83119
rect -45180 -103119 -45178 -83119
rect -45114 -103119 -45112 -83119
rect -13180 -103119 -13178 -83119
rect -13114 -103119 -13112 -83119
rect 18820 -103119 18822 -83119
rect 18886 -103119 18888 -83119
rect 50820 -103119 50822 -83119
rect 50886 -103119 50888 -83119
rect 82820 -103119 82822 -83119
rect 82886 -103119 82888 -83119
rect 114820 -103119 114822 -83119
rect 114886 -103119 114888 -83119
rect 146820 -103119 146822 -83119
rect 146886 -103119 146888 -83119
rect -50075 -106193 -50031 -106185
rect -49975 -106193 -49931 -106185
rect -49875 -106193 -49831 -106185
rect -49775 -106193 -49731 -106185
rect -49675 -106193 -49631 -106185
rect -49575 -106193 -49531 -106185
rect -49475 -106193 -49431 -106185
rect -49375 -106193 -49331 -106185
rect -49275 -106193 -49231 -106185
rect -49175 -106193 -49131 -106185
rect -49075 -106193 -49031 -106185
rect -48975 -106193 -48931 -106185
rect -48875 -106193 -48831 -106185
rect -48775 -106193 -48731 -106185
rect -48675 -106193 -48631 -106185
rect -48575 -106193 -48531 -106185
rect -48075 -106193 -48031 -106185
rect -47975 -106193 -47931 -106185
rect -47875 -106193 -47831 -106185
rect -47775 -106193 -47731 -106185
rect -47675 -106193 -47631 -106185
rect -47575 -106193 -47531 -106185
rect -47475 -106193 -47431 -106185
rect -47375 -106193 -47331 -106185
rect -47275 -106193 -47231 -106185
rect -47175 -106193 -47131 -106185
rect -47075 -106193 -47031 -106185
rect -46975 -106193 -46931 -106185
rect -46875 -106193 -46831 -106185
rect -46775 -106193 -46731 -106185
rect -46675 -106193 -46631 -106185
rect -46575 -106193 -46531 -106185
rect -46075 -106193 -46031 -106185
rect -45975 -106193 -45931 -106185
rect -45875 -106193 -45831 -106185
rect -45775 -106193 -45731 -106185
rect -45675 -106193 -45631 -106185
rect -45575 -106193 -45531 -106185
rect -45475 -106193 -45431 -106185
rect -45375 -106193 -45331 -106185
rect -45275 -106193 -45231 -106185
rect -45175 -106193 -45131 -106185
rect -45075 -106193 -45031 -106185
rect -44975 -106193 -44931 -106185
rect -44875 -106193 -44831 -106185
rect -44775 -106193 -44731 -106185
rect -44675 -106193 -44631 -106185
rect -44575 -106193 -44531 -106185
rect -44075 -106193 -44031 -106185
rect -43975 -106193 -43931 -106185
rect -43875 -106193 -43831 -106185
rect -43775 -106193 -43731 -106185
rect -43675 -106193 -43631 -106185
rect -43575 -106193 -43531 -106185
rect -43475 -106193 -43431 -106185
rect -43375 -106193 -43331 -106185
rect -43275 -106193 -43231 -106185
rect -43175 -106193 -43131 -106185
rect -43075 -106193 -43031 -106185
rect -42975 -106193 -42931 -106185
rect -42875 -106193 -42831 -106185
rect -42775 -106193 -42731 -106185
rect -42675 -106193 -42631 -106185
rect -42575 -106193 -42531 -106185
rect -50031 -106237 -50023 -106193
rect -49931 -106237 -49923 -106193
rect -49831 -106237 -49823 -106193
rect -49731 -106237 -49723 -106193
rect -49631 -106237 -49623 -106193
rect -49531 -106237 -49523 -106193
rect -49431 -106237 -49423 -106193
rect -49331 -106237 -49323 -106193
rect -49231 -106237 -49223 -106193
rect -49131 -106237 -49123 -106193
rect -49031 -106237 -49023 -106193
rect -48931 -106237 -48923 -106193
rect -48831 -106237 -48823 -106193
rect -48731 -106237 -48723 -106193
rect -48631 -106237 -48623 -106193
rect -48531 -106237 -48523 -106193
rect -48031 -106237 -48023 -106193
rect -47931 -106237 -47923 -106193
rect -47831 -106237 -47823 -106193
rect -47731 -106237 -47723 -106193
rect -47631 -106237 -47623 -106193
rect -47531 -106237 -47523 -106193
rect -47431 -106237 -47423 -106193
rect -47331 -106237 -47323 -106193
rect -47231 -106237 -47223 -106193
rect -47131 -106237 -47123 -106193
rect -47031 -106237 -47023 -106193
rect -46931 -106237 -46923 -106193
rect -46831 -106237 -46823 -106193
rect -46731 -106237 -46723 -106193
rect -46631 -106237 -46623 -106193
rect -46531 -106237 -46523 -106193
rect -46031 -106237 -46023 -106193
rect -45931 -106237 -45923 -106193
rect -45831 -106237 -45823 -106193
rect -45731 -106237 -45723 -106193
rect -45631 -106237 -45623 -106193
rect -45531 -106237 -45523 -106193
rect -45431 -106237 -45423 -106193
rect -45331 -106237 -45323 -106193
rect -45231 -106237 -45223 -106193
rect -45131 -106237 -45123 -106193
rect -45031 -106237 -45023 -106193
rect -44931 -106237 -44923 -106193
rect -44831 -106237 -44823 -106193
rect -44731 -106237 -44723 -106193
rect -44631 -106237 -44623 -106193
rect -44531 -106237 -44523 -106193
rect -44031 -106237 -44023 -106193
rect -43931 -106237 -43923 -106193
rect -43831 -106237 -43823 -106193
rect -43731 -106237 -43723 -106193
rect -43631 -106237 -43623 -106193
rect -43531 -106237 -43523 -106193
rect -43431 -106237 -43423 -106193
rect -43331 -106237 -43323 -106193
rect -43231 -106237 -43223 -106193
rect -43131 -106237 -43123 -106193
rect -43031 -106237 -43023 -106193
rect -42931 -106237 -42923 -106193
rect -42831 -106237 -42823 -106193
rect -42731 -106237 -42723 -106193
rect -42631 -106237 -42623 -106193
rect -42531 -106237 -42523 -106193
rect -50075 -106293 -50031 -106285
rect -49975 -106293 -49931 -106285
rect -49875 -106293 -49831 -106285
rect -49775 -106293 -49731 -106285
rect -49675 -106293 -49631 -106285
rect -49575 -106293 -49531 -106285
rect -49475 -106293 -49431 -106285
rect -49375 -106293 -49331 -106285
rect -49275 -106293 -49231 -106285
rect -49175 -106293 -49131 -106285
rect -49075 -106293 -49031 -106285
rect -48975 -106293 -48931 -106285
rect -48875 -106293 -48831 -106285
rect -48775 -106293 -48731 -106285
rect -48675 -106293 -48631 -106285
rect -48575 -106293 -48531 -106285
rect -48075 -106293 -48031 -106285
rect -47975 -106293 -47931 -106285
rect -47875 -106293 -47831 -106285
rect -47775 -106293 -47731 -106285
rect -47675 -106293 -47631 -106285
rect -47575 -106293 -47531 -106285
rect -47475 -106293 -47431 -106285
rect -47375 -106293 -47331 -106285
rect -47275 -106293 -47231 -106285
rect -47175 -106293 -47131 -106285
rect -47075 -106293 -47031 -106285
rect -46975 -106293 -46931 -106285
rect -46875 -106293 -46831 -106285
rect -46775 -106293 -46731 -106285
rect -46675 -106293 -46631 -106285
rect -46575 -106293 -46531 -106285
rect -46075 -106293 -46031 -106285
rect -45975 -106293 -45931 -106285
rect -45875 -106293 -45831 -106285
rect -45775 -106293 -45731 -106285
rect -45675 -106293 -45631 -106285
rect -45575 -106293 -45531 -106285
rect -45475 -106293 -45431 -106285
rect -45375 -106293 -45331 -106285
rect -45275 -106293 -45231 -106285
rect -45175 -106293 -45131 -106285
rect -45075 -106293 -45031 -106285
rect -44975 -106293 -44931 -106285
rect -44875 -106293 -44831 -106285
rect -44775 -106293 -44731 -106285
rect -44675 -106293 -44631 -106285
rect -44575 -106293 -44531 -106285
rect -44075 -106293 -44031 -106285
rect -43975 -106293 -43931 -106285
rect -43875 -106293 -43831 -106285
rect -43775 -106293 -43731 -106285
rect -43675 -106293 -43631 -106285
rect -43575 -106293 -43531 -106285
rect -43475 -106293 -43431 -106285
rect -43375 -106293 -43331 -106285
rect -43275 -106293 -43231 -106285
rect -43175 -106293 -43131 -106285
rect -43075 -106293 -43031 -106285
rect -42975 -106293 -42931 -106285
rect -42875 -106293 -42831 -106285
rect -42775 -106293 -42731 -106285
rect -42675 -106293 -42631 -106285
rect -42575 -106293 -42531 -106285
rect -50031 -106337 -50023 -106293
rect -49931 -106337 -49923 -106293
rect -49831 -106337 -49823 -106293
rect -49731 -106337 -49723 -106293
rect -49631 -106337 -49623 -106293
rect -49531 -106337 -49523 -106293
rect -49431 -106337 -49423 -106293
rect -49331 -106337 -49323 -106293
rect -49231 -106337 -49223 -106293
rect -49131 -106337 -49123 -106293
rect -49031 -106337 -49023 -106293
rect -48931 -106337 -48923 -106293
rect -48831 -106337 -48823 -106293
rect -48731 -106337 -48723 -106293
rect -48631 -106337 -48623 -106293
rect -48531 -106337 -48523 -106293
rect -48031 -106337 -48023 -106293
rect -47931 -106337 -47923 -106293
rect -47831 -106337 -47823 -106293
rect -47731 -106337 -47723 -106293
rect -47631 -106337 -47623 -106293
rect -47531 -106337 -47523 -106293
rect -47431 -106337 -47423 -106293
rect -47331 -106337 -47323 -106293
rect -47231 -106337 -47223 -106293
rect -47131 -106337 -47123 -106293
rect -47031 -106337 -47023 -106293
rect -46931 -106337 -46923 -106293
rect -46831 -106337 -46823 -106293
rect -46731 -106337 -46723 -106293
rect -46631 -106337 -46623 -106293
rect -46531 -106337 -46523 -106293
rect -46031 -106337 -46023 -106293
rect -45931 -106337 -45923 -106293
rect -45831 -106337 -45823 -106293
rect -45731 -106337 -45723 -106293
rect -45631 -106337 -45623 -106293
rect -45531 -106337 -45523 -106293
rect -45431 -106337 -45423 -106293
rect -45331 -106337 -45323 -106293
rect -45231 -106337 -45223 -106293
rect -45131 -106337 -45123 -106293
rect -45031 -106337 -45023 -106293
rect -44931 -106337 -44923 -106293
rect -44831 -106337 -44823 -106293
rect -44731 -106337 -44723 -106293
rect -44631 -106337 -44623 -106293
rect -44531 -106337 -44523 -106293
rect -44031 -106337 -44023 -106293
rect -43931 -106337 -43923 -106293
rect -43831 -106337 -43823 -106293
rect -43731 -106337 -43723 -106293
rect -43631 -106337 -43623 -106293
rect -43531 -106337 -43523 -106293
rect -43431 -106337 -43423 -106293
rect -43331 -106337 -43323 -106293
rect -43231 -106337 -43223 -106293
rect -43131 -106337 -43123 -106293
rect -43031 -106337 -43023 -106293
rect -42931 -106337 -42923 -106293
rect -42831 -106337 -42823 -106293
rect -42731 -106337 -42723 -106293
rect -42631 -106337 -42623 -106293
rect -42531 -106337 -42523 -106293
rect -50075 -106393 -50031 -106385
rect -49975 -106393 -49931 -106385
rect -49875 -106393 -49831 -106385
rect -49775 -106393 -49731 -106385
rect -49675 -106393 -49631 -106385
rect -49575 -106393 -49531 -106385
rect -49475 -106393 -49431 -106385
rect -49375 -106393 -49331 -106385
rect -49275 -106393 -49231 -106385
rect -49175 -106393 -49131 -106385
rect -49075 -106393 -49031 -106385
rect -48975 -106393 -48931 -106385
rect -48875 -106393 -48831 -106385
rect -48775 -106393 -48731 -106385
rect -48675 -106393 -48631 -106385
rect -48575 -106393 -48531 -106385
rect -48075 -106393 -48031 -106385
rect -47975 -106393 -47931 -106385
rect -47875 -106393 -47831 -106385
rect -47775 -106393 -47731 -106385
rect -47675 -106393 -47631 -106385
rect -47575 -106393 -47531 -106385
rect -47475 -106393 -47431 -106385
rect -47375 -106393 -47331 -106385
rect -47275 -106393 -47231 -106385
rect -47175 -106393 -47131 -106385
rect -47075 -106393 -47031 -106385
rect -46975 -106393 -46931 -106385
rect -46875 -106393 -46831 -106385
rect -46775 -106393 -46731 -106385
rect -46675 -106393 -46631 -106385
rect -46575 -106393 -46531 -106385
rect -46075 -106393 -46031 -106385
rect -45975 -106393 -45931 -106385
rect -45875 -106393 -45831 -106385
rect -45775 -106393 -45731 -106385
rect -45675 -106393 -45631 -106385
rect -45575 -106393 -45531 -106385
rect -45475 -106393 -45431 -106385
rect -45375 -106393 -45331 -106385
rect -45275 -106393 -45231 -106385
rect -45175 -106393 -45131 -106385
rect -45075 -106393 -45031 -106385
rect -44975 -106393 -44931 -106385
rect -44875 -106393 -44831 -106385
rect -44775 -106393 -44731 -106385
rect -44675 -106393 -44631 -106385
rect -44575 -106393 -44531 -106385
rect -44075 -106393 -44031 -106385
rect -43975 -106393 -43931 -106385
rect -43875 -106393 -43831 -106385
rect -43775 -106393 -43731 -106385
rect -43675 -106393 -43631 -106385
rect -43575 -106393 -43531 -106385
rect -43475 -106393 -43431 -106385
rect -43375 -106393 -43331 -106385
rect -43275 -106393 -43231 -106385
rect -43175 -106393 -43131 -106385
rect -43075 -106393 -43031 -106385
rect -42975 -106393 -42931 -106385
rect -42875 -106393 -42831 -106385
rect -42775 -106393 -42731 -106385
rect -42675 -106393 -42631 -106385
rect -42575 -106393 -42531 -106385
rect -50031 -106437 -50023 -106393
rect -49931 -106437 -49923 -106393
rect -49831 -106437 -49823 -106393
rect -49731 -106437 -49723 -106393
rect -49631 -106437 -49623 -106393
rect -49531 -106437 -49523 -106393
rect -49431 -106437 -49423 -106393
rect -49331 -106437 -49323 -106393
rect -49231 -106437 -49223 -106393
rect -49131 -106437 -49123 -106393
rect -49031 -106437 -49023 -106393
rect -48931 -106437 -48923 -106393
rect -48831 -106437 -48823 -106393
rect -48731 -106437 -48723 -106393
rect -48631 -106437 -48623 -106393
rect -48531 -106437 -48523 -106393
rect -48031 -106437 -48023 -106393
rect -47931 -106437 -47923 -106393
rect -47831 -106437 -47823 -106393
rect -47731 -106437 -47723 -106393
rect -47631 -106437 -47623 -106393
rect -47531 -106437 -47523 -106393
rect -47431 -106437 -47423 -106393
rect -47331 -106437 -47323 -106393
rect -47231 -106437 -47223 -106393
rect -47131 -106437 -47123 -106393
rect -47031 -106437 -47023 -106393
rect -46931 -106437 -46923 -106393
rect -46831 -106437 -46823 -106393
rect -46731 -106437 -46723 -106393
rect -46631 -106437 -46623 -106393
rect -46531 -106437 -46523 -106393
rect -46031 -106437 -46023 -106393
rect -45931 -106437 -45923 -106393
rect -45831 -106437 -45823 -106393
rect -45731 -106437 -45723 -106393
rect -45631 -106437 -45623 -106393
rect -45531 -106437 -45523 -106393
rect -45431 -106437 -45423 -106393
rect -45331 -106437 -45323 -106393
rect -45231 -106437 -45223 -106393
rect -45131 -106437 -45123 -106393
rect -45031 -106437 -45023 -106393
rect -44931 -106437 -44923 -106393
rect -44831 -106437 -44823 -106393
rect -44731 -106437 -44723 -106393
rect -44631 -106437 -44623 -106393
rect -44531 -106437 -44523 -106393
rect -44031 -106437 -44023 -106393
rect -43931 -106437 -43923 -106393
rect -43831 -106437 -43823 -106393
rect -43731 -106437 -43723 -106393
rect -43631 -106437 -43623 -106393
rect -43531 -106437 -43523 -106393
rect -43431 -106437 -43423 -106393
rect -43331 -106437 -43323 -106393
rect -43231 -106437 -43223 -106393
rect -43131 -106437 -43123 -106393
rect -43031 -106437 -43023 -106393
rect -42931 -106437 -42923 -106393
rect -42831 -106437 -42823 -106393
rect -42731 -106437 -42723 -106393
rect -42631 -106437 -42623 -106393
rect -42531 -106437 -42523 -106393
rect -50075 -106493 -50031 -106485
rect -49975 -106493 -49931 -106485
rect -49875 -106493 -49831 -106485
rect -49775 -106493 -49731 -106485
rect -49675 -106493 -49631 -106485
rect -49575 -106493 -49531 -106485
rect -49475 -106493 -49431 -106485
rect -49375 -106493 -49331 -106485
rect -49275 -106493 -49231 -106485
rect -49175 -106493 -49131 -106485
rect -49075 -106493 -49031 -106485
rect -48975 -106493 -48931 -106485
rect -48875 -106493 -48831 -106485
rect -48775 -106493 -48731 -106485
rect -48675 -106493 -48631 -106485
rect -48575 -106493 -48531 -106485
rect -48075 -106493 -48031 -106485
rect -47975 -106493 -47931 -106485
rect -47875 -106493 -47831 -106485
rect -47775 -106493 -47731 -106485
rect -47675 -106493 -47631 -106485
rect -47575 -106493 -47531 -106485
rect -47475 -106493 -47431 -106485
rect -47375 -106493 -47331 -106485
rect -47275 -106493 -47231 -106485
rect -47175 -106493 -47131 -106485
rect -47075 -106493 -47031 -106485
rect -46975 -106493 -46931 -106485
rect -46875 -106493 -46831 -106485
rect -46775 -106493 -46731 -106485
rect -46675 -106493 -46631 -106485
rect -46575 -106493 -46531 -106485
rect -46075 -106493 -46031 -106485
rect -45975 -106493 -45931 -106485
rect -45875 -106493 -45831 -106485
rect -45775 -106493 -45731 -106485
rect -45675 -106493 -45631 -106485
rect -45575 -106493 -45531 -106485
rect -45475 -106493 -45431 -106485
rect -45375 -106493 -45331 -106485
rect -45275 -106493 -45231 -106485
rect -45175 -106493 -45131 -106485
rect -45075 -106493 -45031 -106485
rect -44975 -106493 -44931 -106485
rect -44875 -106493 -44831 -106485
rect -44775 -106493 -44731 -106485
rect -44675 -106493 -44631 -106485
rect -44575 -106493 -44531 -106485
rect -44075 -106493 -44031 -106485
rect -43975 -106493 -43931 -106485
rect -43875 -106493 -43831 -106485
rect -43775 -106493 -43731 -106485
rect -43675 -106493 -43631 -106485
rect -43575 -106493 -43531 -106485
rect -43475 -106493 -43431 -106485
rect -43375 -106493 -43331 -106485
rect -43275 -106493 -43231 -106485
rect -43175 -106493 -43131 -106485
rect -43075 -106493 -43031 -106485
rect -42975 -106493 -42931 -106485
rect -42875 -106493 -42831 -106485
rect -42775 -106493 -42731 -106485
rect -42675 -106493 -42631 -106485
rect -42575 -106493 -42531 -106485
rect -50031 -106537 -50023 -106493
rect -49931 -106537 -49923 -106493
rect -49831 -106537 -49823 -106493
rect -49731 -106537 -49723 -106493
rect -49631 -106537 -49623 -106493
rect -49531 -106537 -49523 -106493
rect -49431 -106537 -49423 -106493
rect -49331 -106537 -49323 -106493
rect -49231 -106537 -49223 -106493
rect -49131 -106537 -49123 -106493
rect -49031 -106537 -49023 -106493
rect -48931 -106537 -48923 -106493
rect -48831 -106537 -48823 -106493
rect -48731 -106537 -48723 -106493
rect -48631 -106537 -48623 -106493
rect -48531 -106537 -48523 -106493
rect -48031 -106537 -48023 -106493
rect -47931 -106537 -47923 -106493
rect -47831 -106537 -47823 -106493
rect -47731 -106537 -47723 -106493
rect -47631 -106537 -47623 -106493
rect -47531 -106537 -47523 -106493
rect -47431 -106537 -47423 -106493
rect -47331 -106537 -47323 -106493
rect -47231 -106537 -47223 -106493
rect -47131 -106537 -47123 -106493
rect -47031 -106537 -47023 -106493
rect -46931 -106537 -46923 -106493
rect -46831 -106537 -46823 -106493
rect -46731 -106537 -46723 -106493
rect -46631 -106537 -46623 -106493
rect -46531 -106537 -46523 -106493
rect -46031 -106537 -46023 -106493
rect -45931 -106537 -45923 -106493
rect -45831 -106537 -45823 -106493
rect -45731 -106537 -45723 -106493
rect -45631 -106537 -45623 -106493
rect -45531 -106537 -45523 -106493
rect -45431 -106537 -45423 -106493
rect -45331 -106537 -45323 -106493
rect -45231 -106537 -45223 -106493
rect -45131 -106537 -45123 -106493
rect -45031 -106537 -45023 -106493
rect -44931 -106537 -44923 -106493
rect -44831 -106537 -44823 -106493
rect -44731 -106537 -44723 -106493
rect -44631 -106537 -44623 -106493
rect -44531 -106537 -44523 -106493
rect -44031 -106537 -44023 -106493
rect -43931 -106537 -43923 -106493
rect -43831 -106537 -43823 -106493
rect -43731 -106537 -43723 -106493
rect -43631 -106537 -43623 -106493
rect -43531 -106537 -43523 -106493
rect -43431 -106537 -43423 -106493
rect -43331 -106537 -43323 -106493
rect -43231 -106537 -43223 -106493
rect -43131 -106537 -43123 -106493
rect -43031 -106537 -43023 -106493
rect -42931 -106537 -42923 -106493
rect -42831 -106537 -42823 -106493
rect -42731 -106537 -42723 -106493
rect -42631 -106537 -42623 -106493
rect -42531 -106537 -42523 -106493
rect -50075 -106593 -50031 -106585
rect -49975 -106593 -49931 -106585
rect -49875 -106593 -49831 -106585
rect -49775 -106593 -49731 -106585
rect -49675 -106593 -49631 -106585
rect -49575 -106593 -49531 -106585
rect -49475 -106593 -49431 -106585
rect -49375 -106593 -49331 -106585
rect -49275 -106593 -49231 -106585
rect -49175 -106593 -49131 -106585
rect -49075 -106593 -49031 -106585
rect -48975 -106593 -48931 -106585
rect -48875 -106593 -48831 -106585
rect -48775 -106593 -48731 -106585
rect -48675 -106593 -48631 -106585
rect -48575 -106593 -48531 -106585
rect -48075 -106593 -48031 -106585
rect -47975 -106593 -47931 -106585
rect -47875 -106593 -47831 -106585
rect -47775 -106593 -47731 -106585
rect -47675 -106593 -47631 -106585
rect -47575 -106593 -47531 -106585
rect -47475 -106593 -47431 -106585
rect -47375 -106593 -47331 -106585
rect -47275 -106593 -47231 -106585
rect -47175 -106593 -47131 -106585
rect -47075 -106593 -47031 -106585
rect -46975 -106593 -46931 -106585
rect -46875 -106593 -46831 -106585
rect -46775 -106593 -46731 -106585
rect -46675 -106593 -46631 -106585
rect -46575 -106593 -46531 -106585
rect -46075 -106593 -46031 -106585
rect -45975 -106593 -45931 -106585
rect -45875 -106593 -45831 -106585
rect -45775 -106593 -45731 -106585
rect -45675 -106593 -45631 -106585
rect -45575 -106593 -45531 -106585
rect -45475 -106593 -45431 -106585
rect -45375 -106593 -45331 -106585
rect -45275 -106593 -45231 -106585
rect -45175 -106593 -45131 -106585
rect -45075 -106593 -45031 -106585
rect -44975 -106593 -44931 -106585
rect -44875 -106593 -44831 -106585
rect -44775 -106593 -44731 -106585
rect -44675 -106593 -44631 -106585
rect -44575 -106593 -44531 -106585
rect -44075 -106593 -44031 -106585
rect -43975 -106593 -43931 -106585
rect -43875 -106593 -43831 -106585
rect -43775 -106593 -43731 -106585
rect -43675 -106593 -43631 -106585
rect -43575 -106593 -43531 -106585
rect -43475 -106593 -43431 -106585
rect -43375 -106593 -43331 -106585
rect -43275 -106593 -43231 -106585
rect -43175 -106593 -43131 -106585
rect -43075 -106593 -43031 -106585
rect -42975 -106593 -42931 -106585
rect -42875 -106593 -42831 -106585
rect -42775 -106593 -42731 -106585
rect -42675 -106593 -42631 -106585
rect -42575 -106593 -42531 -106585
rect -50031 -106637 -50023 -106593
rect -49931 -106637 -49923 -106593
rect -49831 -106637 -49823 -106593
rect -49731 -106637 -49723 -106593
rect -49631 -106637 -49623 -106593
rect -49531 -106637 -49523 -106593
rect -49431 -106637 -49423 -106593
rect -49331 -106637 -49323 -106593
rect -49231 -106637 -49223 -106593
rect -49131 -106637 -49123 -106593
rect -49031 -106637 -49023 -106593
rect -48931 -106637 -48923 -106593
rect -48831 -106637 -48823 -106593
rect -48731 -106637 -48723 -106593
rect -48631 -106637 -48623 -106593
rect -48531 -106637 -48523 -106593
rect -48031 -106637 -48023 -106593
rect -47931 -106637 -47923 -106593
rect -47831 -106637 -47823 -106593
rect -47731 -106637 -47723 -106593
rect -47631 -106637 -47623 -106593
rect -47531 -106637 -47523 -106593
rect -47431 -106637 -47423 -106593
rect -47331 -106637 -47323 -106593
rect -47231 -106637 -47223 -106593
rect -47131 -106637 -47123 -106593
rect -47031 -106637 -47023 -106593
rect -46931 -106637 -46923 -106593
rect -46831 -106637 -46823 -106593
rect -46731 -106637 -46723 -106593
rect -46631 -106637 -46623 -106593
rect -46531 -106637 -46523 -106593
rect -46031 -106637 -46023 -106593
rect -45931 -106637 -45923 -106593
rect -45831 -106637 -45823 -106593
rect -45731 -106637 -45723 -106593
rect -45631 -106637 -45623 -106593
rect -45531 -106637 -45523 -106593
rect -45431 -106637 -45423 -106593
rect -45331 -106637 -45323 -106593
rect -45231 -106637 -45223 -106593
rect -45131 -106637 -45123 -106593
rect -45031 -106637 -45023 -106593
rect -44931 -106637 -44923 -106593
rect -44831 -106637 -44823 -106593
rect -44731 -106637 -44723 -106593
rect -44631 -106637 -44623 -106593
rect -44531 -106637 -44523 -106593
rect -44031 -106637 -44023 -106593
rect -43931 -106637 -43923 -106593
rect -43831 -106637 -43823 -106593
rect -43731 -106637 -43723 -106593
rect -43631 -106637 -43623 -106593
rect -43531 -106637 -43523 -106593
rect -43431 -106637 -43423 -106593
rect -43331 -106637 -43323 -106593
rect -43231 -106637 -43223 -106593
rect -43131 -106637 -43123 -106593
rect -43031 -106637 -43023 -106593
rect -42931 -106637 -42923 -106593
rect -42831 -106637 -42823 -106593
rect -42731 -106637 -42723 -106593
rect -42631 -106637 -42623 -106593
rect -42531 -106637 -42523 -106593
rect -50075 -106693 -50031 -106685
rect -49975 -106693 -49931 -106685
rect -49875 -106693 -49831 -106685
rect -49775 -106693 -49731 -106685
rect -49675 -106693 -49631 -106685
rect -49575 -106693 -49531 -106685
rect -49475 -106693 -49431 -106685
rect -49375 -106693 -49331 -106685
rect -49275 -106693 -49231 -106685
rect -49175 -106693 -49131 -106685
rect -49075 -106693 -49031 -106685
rect -48975 -106693 -48931 -106685
rect -48875 -106693 -48831 -106685
rect -48775 -106693 -48731 -106685
rect -48675 -106693 -48631 -106685
rect -48575 -106693 -48531 -106685
rect -48075 -106693 -48031 -106685
rect -47975 -106693 -47931 -106685
rect -47875 -106693 -47831 -106685
rect -47775 -106693 -47731 -106685
rect -47675 -106693 -47631 -106685
rect -47575 -106693 -47531 -106685
rect -47475 -106693 -47431 -106685
rect -47375 -106693 -47331 -106685
rect -47275 -106693 -47231 -106685
rect -47175 -106693 -47131 -106685
rect -47075 -106693 -47031 -106685
rect -46975 -106693 -46931 -106685
rect -46875 -106693 -46831 -106685
rect -46775 -106693 -46731 -106685
rect -46675 -106693 -46631 -106685
rect -46575 -106693 -46531 -106685
rect -46075 -106693 -46031 -106685
rect -45975 -106693 -45931 -106685
rect -45875 -106693 -45831 -106685
rect -45775 -106693 -45731 -106685
rect -45675 -106693 -45631 -106685
rect -45575 -106693 -45531 -106685
rect -45475 -106693 -45431 -106685
rect -45375 -106693 -45331 -106685
rect -45275 -106693 -45231 -106685
rect -45175 -106693 -45131 -106685
rect -45075 -106693 -45031 -106685
rect -44975 -106693 -44931 -106685
rect -44875 -106693 -44831 -106685
rect -44775 -106693 -44731 -106685
rect -44675 -106693 -44631 -106685
rect -44575 -106693 -44531 -106685
rect -44075 -106693 -44031 -106685
rect -43975 -106693 -43931 -106685
rect -43875 -106693 -43831 -106685
rect -43775 -106693 -43731 -106685
rect -43675 -106693 -43631 -106685
rect -43575 -106693 -43531 -106685
rect -43475 -106693 -43431 -106685
rect -43375 -106693 -43331 -106685
rect -43275 -106693 -43231 -106685
rect -43175 -106693 -43131 -106685
rect -43075 -106693 -43031 -106685
rect -42975 -106693 -42931 -106685
rect -42875 -106693 -42831 -106685
rect -42775 -106693 -42731 -106685
rect -42675 -106693 -42631 -106685
rect -42575 -106693 -42531 -106685
rect -50031 -106737 -50023 -106693
rect -49931 -106737 -49923 -106693
rect -49831 -106737 -49823 -106693
rect -49731 -106737 -49723 -106693
rect -49631 -106737 -49623 -106693
rect -49531 -106737 -49523 -106693
rect -49431 -106737 -49423 -106693
rect -49331 -106737 -49323 -106693
rect -49231 -106737 -49223 -106693
rect -49131 -106737 -49123 -106693
rect -49031 -106737 -49023 -106693
rect -48931 -106737 -48923 -106693
rect -48831 -106737 -48823 -106693
rect -48731 -106737 -48723 -106693
rect -48631 -106737 -48623 -106693
rect -48531 -106737 -48523 -106693
rect -48031 -106737 -48023 -106693
rect -47931 -106737 -47923 -106693
rect -47831 -106737 -47823 -106693
rect -47731 -106737 -47723 -106693
rect -47631 -106737 -47623 -106693
rect -47531 -106737 -47523 -106693
rect -47431 -106737 -47423 -106693
rect -47331 -106737 -47323 -106693
rect -47231 -106737 -47223 -106693
rect -47131 -106737 -47123 -106693
rect -47031 -106737 -47023 -106693
rect -46931 -106737 -46923 -106693
rect -46831 -106737 -46823 -106693
rect -46731 -106737 -46723 -106693
rect -46631 -106737 -46623 -106693
rect -46531 -106737 -46523 -106693
rect -46031 -106737 -46023 -106693
rect -45931 -106737 -45923 -106693
rect -45831 -106737 -45823 -106693
rect -45731 -106737 -45723 -106693
rect -45631 -106737 -45623 -106693
rect -45531 -106737 -45523 -106693
rect -45431 -106737 -45423 -106693
rect -45331 -106737 -45323 -106693
rect -45231 -106737 -45223 -106693
rect -45131 -106737 -45123 -106693
rect -45031 -106737 -45023 -106693
rect -44931 -106737 -44923 -106693
rect -44831 -106737 -44823 -106693
rect -44731 -106737 -44723 -106693
rect -44631 -106737 -44623 -106693
rect -44531 -106737 -44523 -106693
rect -44031 -106737 -44023 -106693
rect -43931 -106737 -43923 -106693
rect -43831 -106737 -43823 -106693
rect -43731 -106737 -43723 -106693
rect -43631 -106737 -43623 -106693
rect -43531 -106737 -43523 -106693
rect -43431 -106737 -43423 -106693
rect -43331 -106737 -43323 -106693
rect -43231 -106737 -43223 -106693
rect -43131 -106737 -43123 -106693
rect -43031 -106737 -43023 -106693
rect -42931 -106737 -42923 -106693
rect -42831 -106737 -42823 -106693
rect -42731 -106737 -42723 -106693
rect -42631 -106737 -42623 -106693
rect -42531 -106737 -42523 -106693
rect -50075 -106793 -50031 -106785
rect -49975 -106793 -49931 -106785
rect -49875 -106793 -49831 -106785
rect -49775 -106793 -49731 -106785
rect -49675 -106793 -49631 -106785
rect -49575 -106793 -49531 -106785
rect -49475 -106793 -49431 -106785
rect -49375 -106793 -49331 -106785
rect -49275 -106793 -49231 -106785
rect -49175 -106793 -49131 -106785
rect -49075 -106793 -49031 -106785
rect -48975 -106793 -48931 -106785
rect -48875 -106793 -48831 -106785
rect -48775 -106793 -48731 -106785
rect -48675 -106793 -48631 -106785
rect -48575 -106793 -48531 -106785
rect -48075 -106793 -48031 -106785
rect -47975 -106793 -47931 -106785
rect -47875 -106793 -47831 -106785
rect -47775 -106793 -47731 -106785
rect -47675 -106793 -47631 -106785
rect -47575 -106793 -47531 -106785
rect -47475 -106793 -47431 -106785
rect -47375 -106793 -47331 -106785
rect -47275 -106793 -47231 -106785
rect -47175 -106793 -47131 -106785
rect -47075 -106793 -47031 -106785
rect -46975 -106793 -46931 -106785
rect -46875 -106793 -46831 -106785
rect -46775 -106793 -46731 -106785
rect -46675 -106793 -46631 -106785
rect -46575 -106793 -46531 -106785
rect -46075 -106793 -46031 -106785
rect -45975 -106793 -45931 -106785
rect -45875 -106793 -45831 -106785
rect -45775 -106793 -45731 -106785
rect -45675 -106793 -45631 -106785
rect -45575 -106793 -45531 -106785
rect -45475 -106793 -45431 -106785
rect -45375 -106793 -45331 -106785
rect -45275 -106793 -45231 -106785
rect -45175 -106793 -45131 -106785
rect -45075 -106793 -45031 -106785
rect -44975 -106793 -44931 -106785
rect -44875 -106793 -44831 -106785
rect -44775 -106793 -44731 -106785
rect -44675 -106793 -44631 -106785
rect -44575 -106793 -44531 -106785
rect -44075 -106793 -44031 -106785
rect -43975 -106793 -43931 -106785
rect -43875 -106793 -43831 -106785
rect -43775 -106793 -43731 -106785
rect -43675 -106793 -43631 -106785
rect -43575 -106793 -43531 -106785
rect -43475 -106793 -43431 -106785
rect -43375 -106793 -43331 -106785
rect -43275 -106793 -43231 -106785
rect -43175 -106793 -43131 -106785
rect -43075 -106793 -43031 -106785
rect -42975 -106793 -42931 -106785
rect -42875 -106793 -42831 -106785
rect -42775 -106793 -42731 -106785
rect -42675 -106793 -42631 -106785
rect -42575 -106793 -42531 -106785
rect -50031 -106837 -50023 -106793
rect -49931 -106837 -49923 -106793
rect -49831 -106837 -49823 -106793
rect -49731 -106837 -49723 -106793
rect -49631 -106837 -49623 -106793
rect -49531 -106837 -49523 -106793
rect -49431 -106837 -49423 -106793
rect -49331 -106837 -49323 -106793
rect -49231 -106837 -49223 -106793
rect -49131 -106837 -49123 -106793
rect -49031 -106837 -49023 -106793
rect -48931 -106837 -48923 -106793
rect -48831 -106837 -48823 -106793
rect -48731 -106837 -48723 -106793
rect -48631 -106837 -48623 -106793
rect -48531 -106837 -48523 -106793
rect -48031 -106837 -48023 -106793
rect -47931 -106837 -47923 -106793
rect -47831 -106837 -47823 -106793
rect -47731 -106837 -47723 -106793
rect -47631 -106837 -47623 -106793
rect -47531 -106837 -47523 -106793
rect -47431 -106837 -47423 -106793
rect -47331 -106837 -47323 -106793
rect -47231 -106837 -47223 -106793
rect -47131 -106837 -47123 -106793
rect -47031 -106837 -47023 -106793
rect -46931 -106837 -46923 -106793
rect -46831 -106837 -46823 -106793
rect -46731 -106837 -46723 -106793
rect -46631 -106837 -46623 -106793
rect -46531 -106837 -46523 -106793
rect -46031 -106837 -46023 -106793
rect -45931 -106837 -45923 -106793
rect -45831 -106837 -45823 -106793
rect -45731 -106837 -45723 -106793
rect -45631 -106837 -45623 -106793
rect -45531 -106837 -45523 -106793
rect -45431 -106837 -45423 -106793
rect -45331 -106837 -45323 -106793
rect -45231 -106837 -45223 -106793
rect -45131 -106837 -45123 -106793
rect -45031 -106837 -45023 -106793
rect -44931 -106837 -44923 -106793
rect -44831 -106837 -44823 -106793
rect -44731 -106837 -44723 -106793
rect -44631 -106837 -44623 -106793
rect -44531 -106837 -44523 -106793
rect -44031 -106837 -44023 -106793
rect -43931 -106837 -43923 -106793
rect -43831 -106837 -43823 -106793
rect -43731 -106837 -43723 -106793
rect -43631 -106837 -43623 -106793
rect -43531 -106837 -43523 -106793
rect -43431 -106837 -43423 -106793
rect -43331 -106837 -43323 -106793
rect -43231 -106837 -43223 -106793
rect -43131 -106837 -43123 -106793
rect -43031 -106837 -43023 -106793
rect -42931 -106837 -42923 -106793
rect -42831 -106837 -42823 -106793
rect -42731 -106837 -42723 -106793
rect -42631 -106837 -42623 -106793
rect -42531 -106837 -42523 -106793
rect -50075 -106893 -50031 -106885
rect -49975 -106893 -49931 -106885
rect -49875 -106893 -49831 -106885
rect -49775 -106893 -49731 -106885
rect -49675 -106893 -49631 -106885
rect -49575 -106893 -49531 -106885
rect -49475 -106893 -49431 -106885
rect -49375 -106893 -49331 -106885
rect -49275 -106893 -49231 -106885
rect -49175 -106893 -49131 -106885
rect -49075 -106893 -49031 -106885
rect -48975 -106893 -48931 -106885
rect -48875 -106893 -48831 -106885
rect -48775 -106893 -48731 -106885
rect -48675 -106893 -48631 -106885
rect -48575 -106893 -48531 -106885
rect -48075 -106893 -48031 -106885
rect -47975 -106893 -47931 -106885
rect -47875 -106893 -47831 -106885
rect -47775 -106893 -47731 -106885
rect -47675 -106893 -47631 -106885
rect -47575 -106893 -47531 -106885
rect -47475 -106893 -47431 -106885
rect -47375 -106893 -47331 -106885
rect -47275 -106893 -47231 -106885
rect -47175 -106893 -47131 -106885
rect -47075 -106893 -47031 -106885
rect -46975 -106893 -46931 -106885
rect -46875 -106893 -46831 -106885
rect -46775 -106893 -46731 -106885
rect -46675 -106893 -46631 -106885
rect -46575 -106893 -46531 -106885
rect -46075 -106893 -46031 -106885
rect -45975 -106893 -45931 -106885
rect -45875 -106893 -45831 -106885
rect -45775 -106893 -45731 -106885
rect -45675 -106893 -45631 -106885
rect -45575 -106893 -45531 -106885
rect -45475 -106893 -45431 -106885
rect -45375 -106893 -45331 -106885
rect -45275 -106893 -45231 -106885
rect -45175 -106893 -45131 -106885
rect -45075 -106893 -45031 -106885
rect -44975 -106893 -44931 -106885
rect -44875 -106893 -44831 -106885
rect -44775 -106893 -44731 -106885
rect -44675 -106893 -44631 -106885
rect -44575 -106893 -44531 -106885
rect -44075 -106893 -44031 -106885
rect -43975 -106893 -43931 -106885
rect -43875 -106893 -43831 -106885
rect -43775 -106893 -43731 -106885
rect -43675 -106893 -43631 -106885
rect -43575 -106893 -43531 -106885
rect -43475 -106893 -43431 -106885
rect -43375 -106893 -43331 -106885
rect -43275 -106893 -43231 -106885
rect -43175 -106893 -43131 -106885
rect -43075 -106893 -43031 -106885
rect -42975 -106893 -42931 -106885
rect -42875 -106893 -42831 -106885
rect -42775 -106893 -42731 -106885
rect -42675 -106893 -42631 -106885
rect -42575 -106893 -42531 -106885
rect -50031 -106937 -50023 -106893
rect -49931 -106937 -49923 -106893
rect -49831 -106937 -49823 -106893
rect -49731 -106937 -49723 -106893
rect -49631 -106937 -49623 -106893
rect -49531 -106937 -49523 -106893
rect -49431 -106937 -49423 -106893
rect -49331 -106937 -49323 -106893
rect -49231 -106937 -49223 -106893
rect -49131 -106937 -49123 -106893
rect -49031 -106937 -49023 -106893
rect -48931 -106937 -48923 -106893
rect -48831 -106937 -48823 -106893
rect -48731 -106937 -48723 -106893
rect -48631 -106937 -48623 -106893
rect -48531 -106937 -48523 -106893
rect -48031 -106937 -48023 -106893
rect -47931 -106937 -47923 -106893
rect -47831 -106937 -47823 -106893
rect -47731 -106937 -47723 -106893
rect -47631 -106937 -47623 -106893
rect -47531 -106937 -47523 -106893
rect -47431 -106937 -47423 -106893
rect -47331 -106937 -47323 -106893
rect -47231 -106937 -47223 -106893
rect -47131 -106937 -47123 -106893
rect -47031 -106937 -47023 -106893
rect -46931 -106937 -46923 -106893
rect -46831 -106937 -46823 -106893
rect -46731 -106937 -46723 -106893
rect -46631 -106937 -46623 -106893
rect -46531 -106937 -46523 -106893
rect -46031 -106937 -46023 -106893
rect -45931 -106937 -45923 -106893
rect -45831 -106937 -45823 -106893
rect -45731 -106937 -45723 -106893
rect -45631 -106937 -45623 -106893
rect -45531 -106937 -45523 -106893
rect -45431 -106937 -45423 -106893
rect -45331 -106937 -45323 -106893
rect -45231 -106937 -45223 -106893
rect -45131 -106937 -45123 -106893
rect -45031 -106937 -45023 -106893
rect -44931 -106937 -44923 -106893
rect -44831 -106937 -44823 -106893
rect -44731 -106937 -44723 -106893
rect -44631 -106937 -44623 -106893
rect -44531 -106937 -44523 -106893
rect -44031 -106937 -44023 -106893
rect -43931 -106937 -43923 -106893
rect -43831 -106937 -43823 -106893
rect -43731 -106937 -43723 -106893
rect -43631 -106937 -43623 -106893
rect -43531 -106937 -43523 -106893
rect -43431 -106937 -43423 -106893
rect -43331 -106937 -43323 -106893
rect -43231 -106937 -43223 -106893
rect -43131 -106937 -43123 -106893
rect -43031 -106937 -43023 -106893
rect -42931 -106937 -42923 -106893
rect -42831 -106937 -42823 -106893
rect -42731 -106937 -42723 -106893
rect -42631 -106937 -42623 -106893
rect -42531 -106937 -42523 -106893
rect -50075 -106993 -50031 -106985
rect -49975 -106993 -49931 -106985
rect -49875 -106993 -49831 -106985
rect -49775 -106993 -49731 -106985
rect -49675 -106993 -49631 -106985
rect -49575 -106993 -49531 -106985
rect -49475 -106993 -49431 -106985
rect -49375 -106993 -49331 -106985
rect -49275 -106993 -49231 -106985
rect -49175 -106993 -49131 -106985
rect -49075 -106993 -49031 -106985
rect -48975 -106993 -48931 -106985
rect -48875 -106993 -48831 -106985
rect -48775 -106993 -48731 -106985
rect -48675 -106993 -48631 -106985
rect -48575 -106993 -48531 -106985
rect -48075 -106993 -48031 -106985
rect -47975 -106993 -47931 -106985
rect -47875 -106993 -47831 -106985
rect -47775 -106993 -47731 -106985
rect -47675 -106993 -47631 -106985
rect -47575 -106993 -47531 -106985
rect -47475 -106993 -47431 -106985
rect -47375 -106993 -47331 -106985
rect -47275 -106993 -47231 -106985
rect -47175 -106993 -47131 -106985
rect -47075 -106993 -47031 -106985
rect -46975 -106993 -46931 -106985
rect -46875 -106993 -46831 -106985
rect -46775 -106993 -46731 -106985
rect -46675 -106993 -46631 -106985
rect -46575 -106993 -46531 -106985
rect -46075 -106993 -46031 -106985
rect -45975 -106993 -45931 -106985
rect -45875 -106993 -45831 -106985
rect -45775 -106993 -45731 -106985
rect -45675 -106993 -45631 -106985
rect -45575 -106993 -45531 -106985
rect -45475 -106993 -45431 -106985
rect -45375 -106993 -45331 -106985
rect -45275 -106993 -45231 -106985
rect -45175 -106993 -45131 -106985
rect -45075 -106993 -45031 -106985
rect -44975 -106993 -44931 -106985
rect -44875 -106993 -44831 -106985
rect -44775 -106993 -44731 -106985
rect -44675 -106993 -44631 -106985
rect -44575 -106993 -44531 -106985
rect -44075 -106993 -44031 -106985
rect -43975 -106993 -43931 -106985
rect -43875 -106993 -43831 -106985
rect -43775 -106993 -43731 -106985
rect -43675 -106993 -43631 -106985
rect -43575 -106993 -43531 -106985
rect -43475 -106993 -43431 -106985
rect -43375 -106993 -43331 -106985
rect -43275 -106993 -43231 -106985
rect -43175 -106993 -43131 -106985
rect -43075 -106993 -43031 -106985
rect -42975 -106993 -42931 -106985
rect -42875 -106993 -42831 -106985
rect -42775 -106993 -42731 -106985
rect -42675 -106993 -42631 -106985
rect -42575 -106993 -42531 -106985
rect -50031 -107037 -50023 -106993
rect -49931 -107037 -49923 -106993
rect -49831 -107037 -49823 -106993
rect -49731 -107037 -49723 -106993
rect -49631 -107037 -49623 -106993
rect -49531 -107037 -49523 -106993
rect -49431 -107037 -49423 -106993
rect -49331 -107037 -49323 -106993
rect -49231 -107037 -49223 -106993
rect -49131 -107037 -49123 -106993
rect -49031 -107037 -49023 -106993
rect -48931 -107037 -48923 -106993
rect -48831 -107037 -48823 -106993
rect -48731 -107037 -48723 -106993
rect -48631 -107037 -48623 -106993
rect -48531 -107037 -48523 -106993
rect -48031 -107037 -48023 -106993
rect -47931 -107037 -47923 -106993
rect -47831 -107037 -47823 -106993
rect -47731 -107037 -47723 -106993
rect -47631 -107037 -47623 -106993
rect -47531 -107037 -47523 -106993
rect -47431 -107037 -47423 -106993
rect -47331 -107037 -47323 -106993
rect -47231 -107037 -47223 -106993
rect -47131 -107037 -47123 -106993
rect -47031 -107037 -47023 -106993
rect -46931 -107037 -46923 -106993
rect -46831 -107037 -46823 -106993
rect -46731 -107037 -46723 -106993
rect -46631 -107037 -46623 -106993
rect -46531 -107037 -46523 -106993
rect -46031 -107037 -46023 -106993
rect -45931 -107037 -45923 -106993
rect -45831 -107037 -45823 -106993
rect -45731 -107037 -45723 -106993
rect -45631 -107037 -45623 -106993
rect -45531 -107037 -45523 -106993
rect -45431 -107037 -45423 -106993
rect -45331 -107037 -45323 -106993
rect -45231 -107037 -45223 -106993
rect -45131 -107037 -45123 -106993
rect -45031 -107037 -45023 -106993
rect -44931 -107037 -44923 -106993
rect -44831 -107037 -44823 -106993
rect -44731 -107037 -44723 -106993
rect -44631 -107037 -44623 -106993
rect -44531 -107037 -44523 -106993
rect -44031 -107037 -44023 -106993
rect -43931 -107037 -43923 -106993
rect -43831 -107037 -43823 -106993
rect -43731 -107037 -43723 -106993
rect -43631 -107037 -43623 -106993
rect -43531 -107037 -43523 -106993
rect -43431 -107037 -43423 -106993
rect -43331 -107037 -43323 -106993
rect -43231 -107037 -43223 -106993
rect -43131 -107037 -43123 -106993
rect -43031 -107037 -43023 -106993
rect -42931 -107037 -42923 -106993
rect -42831 -107037 -42823 -106993
rect -42731 -107037 -42723 -106993
rect -42631 -107037 -42623 -106993
rect -42531 -107037 -42523 -106993
rect -50075 -107093 -50031 -107085
rect -49975 -107093 -49931 -107085
rect -49875 -107093 -49831 -107085
rect -49775 -107093 -49731 -107085
rect -49675 -107093 -49631 -107085
rect -49575 -107093 -49531 -107085
rect -49475 -107093 -49431 -107085
rect -49375 -107093 -49331 -107085
rect -49275 -107093 -49231 -107085
rect -49175 -107093 -49131 -107085
rect -49075 -107093 -49031 -107085
rect -48975 -107093 -48931 -107085
rect -48875 -107093 -48831 -107085
rect -48775 -107093 -48731 -107085
rect -48675 -107093 -48631 -107085
rect -48575 -107093 -48531 -107085
rect -48075 -107093 -48031 -107085
rect -47975 -107093 -47931 -107085
rect -47875 -107093 -47831 -107085
rect -47775 -107093 -47731 -107085
rect -47675 -107093 -47631 -107085
rect -47575 -107093 -47531 -107085
rect -47475 -107093 -47431 -107085
rect -47375 -107093 -47331 -107085
rect -47275 -107093 -47231 -107085
rect -47175 -107093 -47131 -107085
rect -47075 -107093 -47031 -107085
rect -46975 -107093 -46931 -107085
rect -46875 -107093 -46831 -107085
rect -46775 -107093 -46731 -107085
rect -46675 -107093 -46631 -107085
rect -46575 -107093 -46531 -107085
rect -46075 -107093 -46031 -107085
rect -45975 -107093 -45931 -107085
rect -45875 -107093 -45831 -107085
rect -45775 -107093 -45731 -107085
rect -45675 -107093 -45631 -107085
rect -45575 -107093 -45531 -107085
rect -45475 -107093 -45431 -107085
rect -45375 -107093 -45331 -107085
rect -45275 -107093 -45231 -107085
rect -45175 -107093 -45131 -107085
rect -45075 -107093 -45031 -107085
rect -44975 -107093 -44931 -107085
rect -44875 -107093 -44831 -107085
rect -44775 -107093 -44731 -107085
rect -44675 -107093 -44631 -107085
rect -44575 -107093 -44531 -107085
rect -44075 -107093 -44031 -107085
rect -43975 -107093 -43931 -107085
rect -43875 -107093 -43831 -107085
rect -43775 -107093 -43731 -107085
rect -43675 -107093 -43631 -107085
rect -43575 -107093 -43531 -107085
rect -43475 -107093 -43431 -107085
rect -43375 -107093 -43331 -107085
rect -43275 -107093 -43231 -107085
rect -43175 -107093 -43131 -107085
rect -43075 -107093 -43031 -107085
rect -42975 -107093 -42931 -107085
rect -42875 -107093 -42831 -107085
rect -42775 -107093 -42731 -107085
rect -42675 -107093 -42631 -107085
rect -42575 -107093 -42531 -107085
rect -50031 -107137 -50023 -107093
rect -49931 -107137 -49923 -107093
rect -49831 -107137 -49823 -107093
rect -49731 -107137 -49723 -107093
rect -49631 -107137 -49623 -107093
rect -49531 -107137 -49523 -107093
rect -49431 -107137 -49423 -107093
rect -49331 -107137 -49323 -107093
rect -49231 -107137 -49223 -107093
rect -49131 -107137 -49123 -107093
rect -49031 -107137 -49023 -107093
rect -48931 -107137 -48923 -107093
rect -48831 -107137 -48823 -107093
rect -48731 -107137 -48723 -107093
rect -48631 -107137 -48623 -107093
rect -48531 -107137 -48523 -107093
rect -48031 -107137 -48023 -107093
rect -47931 -107137 -47923 -107093
rect -47831 -107137 -47823 -107093
rect -47731 -107137 -47723 -107093
rect -47631 -107137 -47623 -107093
rect -47531 -107137 -47523 -107093
rect -47431 -107137 -47423 -107093
rect -47331 -107137 -47323 -107093
rect -47231 -107137 -47223 -107093
rect -47131 -107137 -47123 -107093
rect -47031 -107137 -47023 -107093
rect -46931 -107137 -46923 -107093
rect -46831 -107137 -46823 -107093
rect -46731 -107137 -46723 -107093
rect -46631 -107137 -46623 -107093
rect -46531 -107137 -46523 -107093
rect -46031 -107137 -46023 -107093
rect -45931 -107137 -45923 -107093
rect -45831 -107137 -45823 -107093
rect -45731 -107137 -45723 -107093
rect -45631 -107137 -45623 -107093
rect -45531 -107137 -45523 -107093
rect -45431 -107137 -45423 -107093
rect -45331 -107137 -45323 -107093
rect -45231 -107137 -45223 -107093
rect -45131 -107137 -45123 -107093
rect -45031 -107137 -45023 -107093
rect -44931 -107137 -44923 -107093
rect -44831 -107137 -44823 -107093
rect -44731 -107137 -44723 -107093
rect -44631 -107137 -44623 -107093
rect -44531 -107137 -44523 -107093
rect -44031 -107137 -44023 -107093
rect -43931 -107137 -43923 -107093
rect -43831 -107137 -43823 -107093
rect -43731 -107137 -43723 -107093
rect -43631 -107137 -43623 -107093
rect -43531 -107137 -43523 -107093
rect -43431 -107137 -43423 -107093
rect -43331 -107137 -43323 -107093
rect -43231 -107137 -43223 -107093
rect -43131 -107137 -43123 -107093
rect -43031 -107137 -43023 -107093
rect -42931 -107137 -42923 -107093
rect -42831 -107137 -42823 -107093
rect -42731 -107137 -42723 -107093
rect -42631 -107137 -42623 -107093
rect -42531 -107137 -42523 -107093
rect -50075 -107193 -50031 -107185
rect -49975 -107193 -49931 -107185
rect -49875 -107193 -49831 -107185
rect -49775 -107193 -49731 -107185
rect -49675 -107193 -49631 -107185
rect -49575 -107193 -49531 -107185
rect -49475 -107193 -49431 -107185
rect -49375 -107193 -49331 -107185
rect -49275 -107193 -49231 -107185
rect -49175 -107193 -49131 -107185
rect -49075 -107193 -49031 -107185
rect -48975 -107193 -48931 -107185
rect -48875 -107193 -48831 -107185
rect -48775 -107193 -48731 -107185
rect -48675 -107193 -48631 -107185
rect -48575 -107193 -48531 -107185
rect -48075 -107193 -48031 -107185
rect -47975 -107193 -47931 -107185
rect -47875 -107193 -47831 -107185
rect -47775 -107193 -47731 -107185
rect -47675 -107193 -47631 -107185
rect -47575 -107193 -47531 -107185
rect -47475 -107193 -47431 -107185
rect -47375 -107193 -47331 -107185
rect -47275 -107193 -47231 -107185
rect -47175 -107193 -47131 -107185
rect -47075 -107193 -47031 -107185
rect -46975 -107193 -46931 -107185
rect -46875 -107193 -46831 -107185
rect -46775 -107193 -46731 -107185
rect -46675 -107193 -46631 -107185
rect -46575 -107193 -46531 -107185
rect -46075 -107193 -46031 -107185
rect -45975 -107193 -45931 -107185
rect -45875 -107193 -45831 -107185
rect -45775 -107193 -45731 -107185
rect -45675 -107193 -45631 -107185
rect -45575 -107193 -45531 -107185
rect -45475 -107193 -45431 -107185
rect -45375 -107193 -45331 -107185
rect -45275 -107193 -45231 -107185
rect -45175 -107193 -45131 -107185
rect -45075 -107193 -45031 -107185
rect -44975 -107193 -44931 -107185
rect -44875 -107193 -44831 -107185
rect -44775 -107193 -44731 -107185
rect -44675 -107193 -44631 -107185
rect -44575 -107193 -44531 -107185
rect -44075 -107193 -44031 -107185
rect -43975 -107193 -43931 -107185
rect -43875 -107193 -43831 -107185
rect -43775 -107193 -43731 -107185
rect -43675 -107193 -43631 -107185
rect -43575 -107193 -43531 -107185
rect -43475 -107193 -43431 -107185
rect -43375 -107193 -43331 -107185
rect -43275 -107193 -43231 -107185
rect -43175 -107193 -43131 -107185
rect -43075 -107193 -43031 -107185
rect -42975 -107193 -42931 -107185
rect -42875 -107193 -42831 -107185
rect -42775 -107193 -42731 -107185
rect -42675 -107193 -42631 -107185
rect -42575 -107193 -42531 -107185
rect -50031 -107237 -50023 -107193
rect -49931 -107237 -49923 -107193
rect -49831 -107237 -49823 -107193
rect -49731 -107237 -49723 -107193
rect -49631 -107237 -49623 -107193
rect -49531 -107237 -49523 -107193
rect -49431 -107237 -49423 -107193
rect -49331 -107237 -49323 -107193
rect -49231 -107237 -49223 -107193
rect -49131 -107237 -49123 -107193
rect -49031 -107237 -49023 -107193
rect -48931 -107237 -48923 -107193
rect -48831 -107237 -48823 -107193
rect -48731 -107237 -48723 -107193
rect -48631 -107237 -48623 -107193
rect -48531 -107237 -48523 -107193
rect -48031 -107237 -48023 -107193
rect -47931 -107237 -47923 -107193
rect -47831 -107237 -47823 -107193
rect -47731 -107237 -47723 -107193
rect -47631 -107237 -47623 -107193
rect -47531 -107237 -47523 -107193
rect -47431 -107237 -47423 -107193
rect -47331 -107237 -47323 -107193
rect -47231 -107237 -47223 -107193
rect -47131 -107237 -47123 -107193
rect -47031 -107237 -47023 -107193
rect -46931 -107237 -46923 -107193
rect -46831 -107237 -46823 -107193
rect -46731 -107237 -46723 -107193
rect -46631 -107237 -46623 -107193
rect -46531 -107237 -46523 -107193
rect -46031 -107237 -46023 -107193
rect -45931 -107237 -45923 -107193
rect -45831 -107237 -45823 -107193
rect -45731 -107237 -45723 -107193
rect -45631 -107237 -45623 -107193
rect -45531 -107237 -45523 -107193
rect -45431 -107237 -45423 -107193
rect -45331 -107237 -45323 -107193
rect -45231 -107237 -45223 -107193
rect -45131 -107237 -45123 -107193
rect -45031 -107237 -45023 -107193
rect -44931 -107237 -44923 -107193
rect -44831 -107237 -44823 -107193
rect -44731 -107237 -44723 -107193
rect -44631 -107237 -44623 -107193
rect -44531 -107237 -44523 -107193
rect -44031 -107237 -44023 -107193
rect -43931 -107237 -43923 -107193
rect -43831 -107237 -43823 -107193
rect -43731 -107237 -43723 -107193
rect -43631 -107237 -43623 -107193
rect -43531 -107237 -43523 -107193
rect -43431 -107237 -43423 -107193
rect -43331 -107237 -43323 -107193
rect -43231 -107237 -43223 -107193
rect -43131 -107237 -43123 -107193
rect -43031 -107237 -43023 -107193
rect -42931 -107237 -42923 -107193
rect -42831 -107237 -42823 -107193
rect -42731 -107237 -42723 -107193
rect -42631 -107237 -42623 -107193
rect -42531 -107237 -42523 -107193
rect -50075 -107293 -50031 -107285
rect -49975 -107293 -49931 -107285
rect -49875 -107293 -49831 -107285
rect -49775 -107293 -49731 -107285
rect -49675 -107293 -49631 -107285
rect -49575 -107293 -49531 -107285
rect -49475 -107293 -49431 -107285
rect -49375 -107293 -49331 -107285
rect -49275 -107293 -49231 -107285
rect -49175 -107293 -49131 -107285
rect -49075 -107293 -49031 -107285
rect -48975 -107293 -48931 -107285
rect -48875 -107293 -48831 -107285
rect -48775 -107293 -48731 -107285
rect -48675 -107293 -48631 -107285
rect -48575 -107293 -48531 -107285
rect -48075 -107293 -48031 -107285
rect -47975 -107293 -47931 -107285
rect -47875 -107293 -47831 -107285
rect -47775 -107293 -47731 -107285
rect -47675 -107293 -47631 -107285
rect -47575 -107293 -47531 -107285
rect -47475 -107293 -47431 -107285
rect -47375 -107293 -47331 -107285
rect -47275 -107293 -47231 -107285
rect -47175 -107293 -47131 -107285
rect -47075 -107293 -47031 -107285
rect -46975 -107293 -46931 -107285
rect -46875 -107293 -46831 -107285
rect -46775 -107293 -46731 -107285
rect -46675 -107293 -46631 -107285
rect -46575 -107293 -46531 -107285
rect -46075 -107293 -46031 -107285
rect -45975 -107293 -45931 -107285
rect -45875 -107293 -45831 -107285
rect -45775 -107293 -45731 -107285
rect -45675 -107293 -45631 -107285
rect -45575 -107293 -45531 -107285
rect -45475 -107293 -45431 -107285
rect -45375 -107293 -45331 -107285
rect -45275 -107293 -45231 -107285
rect -45175 -107293 -45131 -107285
rect -45075 -107293 -45031 -107285
rect -44975 -107293 -44931 -107285
rect -44875 -107293 -44831 -107285
rect -44775 -107293 -44731 -107285
rect -44675 -107293 -44631 -107285
rect -44575 -107293 -44531 -107285
rect -44075 -107293 -44031 -107285
rect -43975 -107293 -43931 -107285
rect -43875 -107293 -43831 -107285
rect -43775 -107293 -43731 -107285
rect -43675 -107293 -43631 -107285
rect -43575 -107293 -43531 -107285
rect -43475 -107293 -43431 -107285
rect -43375 -107293 -43331 -107285
rect -43275 -107293 -43231 -107285
rect -43175 -107293 -43131 -107285
rect -43075 -107293 -43031 -107285
rect -42975 -107293 -42931 -107285
rect -42875 -107293 -42831 -107285
rect -42775 -107293 -42731 -107285
rect -42675 -107293 -42631 -107285
rect -42575 -107293 -42531 -107285
rect -50031 -107337 -50023 -107293
rect -49931 -107337 -49923 -107293
rect -49831 -107337 -49823 -107293
rect -49731 -107337 -49723 -107293
rect -49631 -107337 -49623 -107293
rect -49531 -107337 -49523 -107293
rect -49431 -107337 -49423 -107293
rect -49331 -107337 -49323 -107293
rect -49231 -107337 -49223 -107293
rect -49131 -107337 -49123 -107293
rect -49031 -107337 -49023 -107293
rect -48931 -107337 -48923 -107293
rect -48831 -107337 -48823 -107293
rect -48731 -107337 -48723 -107293
rect -48631 -107337 -48623 -107293
rect -48531 -107337 -48523 -107293
rect -48031 -107337 -48023 -107293
rect -47931 -107337 -47923 -107293
rect -47831 -107337 -47823 -107293
rect -47731 -107337 -47723 -107293
rect -47631 -107337 -47623 -107293
rect -47531 -107337 -47523 -107293
rect -47431 -107337 -47423 -107293
rect -47331 -107337 -47323 -107293
rect -47231 -107337 -47223 -107293
rect -47131 -107337 -47123 -107293
rect -47031 -107337 -47023 -107293
rect -46931 -107337 -46923 -107293
rect -46831 -107337 -46823 -107293
rect -46731 -107337 -46723 -107293
rect -46631 -107337 -46623 -107293
rect -46531 -107337 -46523 -107293
rect -46031 -107337 -46023 -107293
rect -45931 -107337 -45923 -107293
rect -45831 -107337 -45823 -107293
rect -45731 -107337 -45723 -107293
rect -45631 -107337 -45623 -107293
rect -45531 -107337 -45523 -107293
rect -45431 -107337 -45423 -107293
rect -45331 -107337 -45323 -107293
rect -45231 -107337 -45223 -107293
rect -45131 -107337 -45123 -107293
rect -45031 -107337 -45023 -107293
rect -44931 -107337 -44923 -107293
rect -44831 -107337 -44823 -107293
rect -44731 -107337 -44723 -107293
rect -44631 -107337 -44623 -107293
rect -44531 -107337 -44523 -107293
rect -44031 -107337 -44023 -107293
rect -43931 -107337 -43923 -107293
rect -43831 -107337 -43823 -107293
rect -43731 -107337 -43723 -107293
rect -43631 -107337 -43623 -107293
rect -43531 -107337 -43523 -107293
rect -43431 -107337 -43423 -107293
rect -43331 -107337 -43323 -107293
rect -43231 -107337 -43223 -107293
rect -43131 -107337 -43123 -107293
rect -43031 -107337 -43023 -107293
rect -42931 -107337 -42923 -107293
rect -42831 -107337 -42823 -107293
rect -42731 -107337 -42723 -107293
rect -42631 -107337 -42623 -107293
rect -42531 -107337 -42523 -107293
rect -50075 -107393 -50031 -107385
rect -49975 -107393 -49931 -107385
rect -49875 -107393 -49831 -107385
rect -49775 -107393 -49731 -107385
rect -49675 -107393 -49631 -107385
rect -49575 -107393 -49531 -107385
rect -49475 -107393 -49431 -107385
rect -49375 -107393 -49331 -107385
rect -49275 -107393 -49231 -107385
rect -49175 -107393 -49131 -107385
rect -49075 -107393 -49031 -107385
rect -48975 -107393 -48931 -107385
rect -48875 -107393 -48831 -107385
rect -48775 -107393 -48731 -107385
rect -48675 -107393 -48631 -107385
rect -48575 -107393 -48531 -107385
rect -48075 -107393 -48031 -107385
rect -47975 -107393 -47931 -107385
rect -47875 -107393 -47831 -107385
rect -47775 -107393 -47731 -107385
rect -47675 -107393 -47631 -107385
rect -47575 -107393 -47531 -107385
rect -47475 -107393 -47431 -107385
rect -47375 -107393 -47331 -107385
rect -47275 -107393 -47231 -107385
rect -47175 -107393 -47131 -107385
rect -47075 -107393 -47031 -107385
rect -46975 -107393 -46931 -107385
rect -46875 -107393 -46831 -107385
rect -46775 -107393 -46731 -107385
rect -46675 -107393 -46631 -107385
rect -46575 -107393 -46531 -107385
rect -46075 -107393 -46031 -107385
rect -45975 -107393 -45931 -107385
rect -45875 -107393 -45831 -107385
rect -45775 -107393 -45731 -107385
rect -45675 -107393 -45631 -107385
rect -45575 -107393 -45531 -107385
rect -45475 -107393 -45431 -107385
rect -45375 -107393 -45331 -107385
rect -45275 -107393 -45231 -107385
rect -45175 -107393 -45131 -107385
rect -45075 -107393 -45031 -107385
rect -44975 -107393 -44931 -107385
rect -44875 -107393 -44831 -107385
rect -44775 -107393 -44731 -107385
rect -44675 -107393 -44631 -107385
rect -44575 -107393 -44531 -107385
rect -44075 -107393 -44031 -107385
rect -43975 -107393 -43931 -107385
rect -43875 -107393 -43831 -107385
rect -43775 -107393 -43731 -107385
rect -43675 -107393 -43631 -107385
rect -43575 -107393 -43531 -107385
rect -43475 -107393 -43431 -107385
rect -43375 -107393 -43331 -107385
rect -43275 -107393 -43231 -107385
rect -43175 -107393 -43131 -107385
rect -43075 -107393 -43031 -107385
rect -42975 -107393 -42931 -107385
rect -42875 -107393 -42831 -107385
rect -42775 -107393 -42731 -107385
rect -42675 -107393 -42631 -107385
rect -42575 -107393 -42531 -107385
rect -50031 -107437 -50023 -107393
rect -49931 -107437 -49923 -107393
rect -49831 -107437 -49823 -107393
rect -49731 -107437 -49723 -107393
rect -49631 -107437 -49623 -107393
rect -49531 -107437 -49523 -107393
rect -49431 -107437 -49423 -107393
rect -49331 -107437 -49323 -107393
rect -49231 -107437 -49223 -107393
rect -49131 -107437 -49123 -107393
rect -49031 -107437 -49023 -107393
rect -48931 -107437 -48923 -107393
rect -48831 -107437 -48823 -107393
rect -48731 -107437 -48723 -107393
rect -48631 -107437 -48623 -107393
rect -48531 -107437 -48523 -107393
rect -48031 -107437 -48023 -107393
rect -47931 -107437 -47923 -107393
rect -47831 -107437 -47823 -107393
rect -47731 -107437 -47723 -107393
rect -47631 -107437 -47623 -107393
rect -47531 -107437 -47523 -107393
rect -47431 -107437 -47423 -107393
rect -47331 -107437 -47323 -107393
rect -47231 -107437 -47223 -107393
rect -47131 -107437 -47123 -107393
rect -47031 -107437 -47023 -107393
rect -46931 -107437 -46923 -107393
rect -46831 -107437 -46823 -107393
rect -46731 -107437 -46723 -107393
rect -46631 -107437 -46623 -107393
rect -46531 -107437 -46523 -107393
rect -46031 -107437 -46023 -107393
rect -45931 -107437 -45923 -107393
rect -45831 -107437 -45823 -107393
rect -45731 -107437 -45723 -107393
rect -45631 -107437 -45623 -107393
rect -45531 -107437 -45523 -107393
rect -45431 -107437 -45423 -107393
rect -45331 -107437 -45323 -107393
rect -45231 -107437 -45223 -107393
rect -45131 -107437 -45123 -107393
rect -45031 -107437 -45023 -107393
rect -44931 -107437 -44923 -107393
rect -44831 -107437 -44823 -107393
rect -44731 -107437 -44723 -107393
rect -44631 -107437 -44623 -107393
rect -44531 -107437 -44523 -107393
rect -44031 -107437 -44023 -107393
rect -43931 -107437 -43923 -107393
rect -43831 -107437 -43823 -107393
rect -43731 -107437 -43723 -107393
rect -43631 -107437 -43623 -107393
rect -43531 -107437 -43523 -107393
rect -43431 -107437 -43423 -107393
rect -43331 -107437 -43323 -107393
rect -43231 -107437 -43223 -107393
rect -43131 -107437 -43123 -107393
rect -43031 -107437 -43023 -107393
rect -42931 -107437 -42923 -107393
rect -42831 -107437 -42823 -107393
rect -42731 -107437 -42723 -107393
rect -42631 -107437 -42623 -107393
rect -42531 -107437 -42523 -107393
rect -50075 -107493 -50031 -107485
rect -49975 -107493 -49931 -107485
rect -49875 -107493 -49831 -107485
rect -49775 -107493 -49731 -107485
rect -49675 -107493 -49631 -107485
rect -49575 -107493 -49531 -107485
rect -49475 -107493 -49431 -107485
rect -49375 -107493 -49331 -107485
rect -49275 -107493 -49231 -107485
rect -49175 -107493 -49131 -107485
rect -49075 -107493 -49031 -107485
rect -48975 -107493 -48931 -107485
rect -48875 -107493 -48831 -107485
rect -48775 -107493 -48731 -107485
rect -48675 -107493 -48631 -107485
rect -48575 -107493 -48531 -107485
rect -48075 -107493 -48031 -107485
rect -47975 -107493 -47931 -107485
rect -47875 -107493 -47831 -107485
rect -47775 -107493 -47731 -107485
rect -47675 -107493 -47631 -107485
rect -47575 -107493 -47531 -107485
rect -47475 -107493 -47431 -107485
rect -47375 -107493 -47331 -107485
rect -47275 -107493 -47231 -107485
rect -47175 -107493 -47131 -107485
rect -47075 -107493 -47031 -107485
rect -46975 -107493 -46931 -107485
rect -46875 -107493 -46831 -107485
rect -46775 -107493 -46731 -107485
rect -46675 -107493 -46631 -107485
rect -46575 -107493 -46531 -107485
rect -46075 -107493 -46031 -107485
rect -45975 -107493 -45931 -107485
rect -45875 -107493 -45831 -107485
rect -45775 -107493 -45731 -107485
rect -45675 -107493 -45631 -107485
rect -45575 -107493 -45531 -107485
rect -45475 -107493 -45431 -107485
rect -45375 -107493 -45331 -107485
rect -45275 -107493 -45231 -107485
rect -45175 -107493 -45131 -107485
rect -45075 -107493 -45031 -107485
rect -44975 -107493 -44931 -107485
rect -44875 -107493 -44831 -107485
rect -44775 -107493 -44731 -107485
rect -44675 -107493 -44631 -107485
rect -44575 -107493 -44531 -107485
rect -44075 -107493 -44031 -107485
rect -43975 -107493 -43931 -107485
rect -43875 -107493 -43831 -107485
rect -43775 -107493 -43731 -107485
rect -43675 -107493 -43631 -107485
rect -43575 -107493 -43531 -107485
rect -43475 -107493 -43431 -107485
rect -43375 -107493 -43331 -107485
rect -43275 -107493 -43231 -107485
rect -43175 -107493 -43131 -107485
rect -43075 -107493 -43031 -107485
rect -42975 -107493 -42931 -107485
rect -42875 -107493 -42831 -107485
rect -42775 -107493 -42731 -107485
rect -42675 -107493 -42631 -107485
rect -42575 -107493 -42531 -107485
rect -50031 -107537 -50023 -107493
rect -49931 -107537 -49923 -107493
rect -49831 -107537 -49823 -107493
rect -49731 -107537 -49723 -107493
rect -49631 -107537 -49623 -107493
rect -49531 -107537 -49523 -107493
rect -49431 -107537 -49423 -107493
rect -49331 -107537 -49323 -107493
rect -49231 -107537 -49223 -107493
rect -49131 -107537 -49123 -107493
rect -49031 -107537 -49023 -107493
rect -48931 -107537 -48923 -107493
rect -48831 -107537 -48823 -107493
rect -48731 -107537 -48723 -107493
rect -48631 -107537 -48623 -107493
rect -48531 -107537 -48523 -107493
rect -48031 -107537 -48023 -107493
rect -47931 -107537 -47923 -107493
rect -47831 -107537 -47823 -107493
rect -47731 -107537 -47723 -107493
rect -47631 -107537 -47623 -107493
rect -47531 -107537 -47523 -107493
rect -47431 -107537 -47423 -107493
rect -47331 -107537 -47323 -107493
rect -47231 -107537 -47223 -107493
rect -47131 -107537 -47123 -107493
rect -47031 -107537 -47023 -107493
rect -46931 -107537 -46923 -107493
rect -46831 -107537 -46823 -107493
rect -46731 -107537 -46723 -107493
rect -46631 -107537 -46623 -107493
rect -46531 -107537 -46523 -107493
rect -46031 -107537 -46023 -107493
rect -45931 -107537 -45923 -107493
rect -45831 -107537 -45823 -107493
rect -45731 -107537 -45723 -107493
rect -45631 -107537 -45623 -107493
rect -45531 -107537 -45523 -107493
rect -45431 -107537 -45423 -107493
rect -45331 -107537 -45323 -107493
rect -45231 -107537 -45223 -107493
rect -45131 -107537 -45123 -107493
rect -45031 -107537 -45023 -107493
rect -44931 -107537 -44923 -107493
rect -44831 -107537 -44823 -107493
rect -44731 -107537 -44723 -107493
rect -44631 -107537 -44623 -107493
rect -44531 -107537 -44523 -107493
rect -44031 -107537 -44023 -107493
rect -43931 -107537 -43923 -107493
rect -43831 -107537 -43823 -107493
rect -43731 -107537 -43723 -107493
rect -43631 -107537 -43623 -107493
rect -43531 -107537 -43523 -107493
rect -43431 -107537 -43423 -107493
rect -43331 -107537 -43323 -107493
rect -43231 -107537 -43223 -107493
rect -43131 -107537 -43123 -107493
rect -43031 -107537 -43023 -107493
rect -42931 -107537 -42923 -107493
rect -42831 -107537 -42823 -107493
rect -42731 -107537 -42723 -107493
rect -42631 -107537 -42623 -107493
rect -42531 -107537 -42523 -107493
rect -50075 -107593 -50031 -107585
rect -49975 -107593 -49931 -107585
rect -49875 -107593 -49831 -107585
rect -49775 -107593 -49731 -107585
rect -49675 -107593 -49631 -107585
rect -49575 -107593 -49531 -107585
rect -49475 -107593 -49431 -107585
rect -49375 -107593 -49331 -107585
rect -49275 -107593 -49231 -107585
rect -49175 -107593 -49131 -107585
rect -49075 -107593 -49031 -107585
rect -48975 -107593 -48931 -107585
rect -48875 -107593 -48831 -107585
rect -48775 -107593 -48731 -107585
rect -48675 -107593 -48631 -107585
rect -48575 -107593 -48531 -107585
rect -48075 -107593 -48031 -107585
rect -47975 -107593 -47931 -107585
rect -47875 -107593 -47831 -107585
rect -47775 -107593 -47731 -107585
rect -47675 -107593 -47631 -107585
rect -47575 -107593 -47531 -107585
rect -47475 -107593 -47431 -107585
rect -47375 -107593 -47331 -107585
rect -47275 -107593 -47231 -107585
rect -47175 -107593 -47131 -107585
rect -47075 -107593 -47031 -107585
rect -46975 -107593 -46931 -107585
rect -46875 -107593 -46831 -107585
rect -46775 -107593 -46731 -107585
rect -46675 -107593 -46631 -107585
rect -46575 -107593 -46531 -107585
rect -46075 -107593 -46031 -107585
rect -45975 -107593 -45931 -107585
rect -45875 -107593 -45831 -107585
rect -45775 -107593 -45731 -107585
rect -45675 -107593 -45631 -107585
rect -45575 -107593 -45531 -107585
rect -45475 -107593 -45431 -107585
rect -45375 -107593 -45331 -107585
rect -45275 -107593 -45231 -107585
rect -45175 -107593 -45131 -107585
rect -45075 -107593 -45031 -107585
rect -44975 -107593 -44931 -107585
rect -44875 -107593 -44831 -107585
rect -44775 -107593 -44731 -107585
rect -44675 -107593 -44631 -107585
rect -44575 -107593 -44531 -107585
rect -44075 -107593 -44031 -107585
rect -43975 -107593 -43931 -107585
rect -43875 -107593 -43831 -107585
rect -43775 -107593 -43731 -107585
rect -43675 -107593 -43631 -107585
rect -43575 -107593 -43531 -107585
rect -43475 -107593 -43431 -107585
rect -43375 -107593 -43331 -107585
rect -43275 -107593 -43231 -107585
rect -43175 -107593 -43131 -107585
rect -43075 -107593 -43031 -107585
rect -42975 -107593 -42931 -107585
rect -42875 -107593 -42831 -107585
rect -42775 -107593 -42731 -107585
rect -42675 -107593 -42631 -107585
rect -42575 -107593 -42531 -107585
rect -50031 -107637 -50023 -107593
rect -49931 -107637 -49923 -107593
rect -49831 -107637 -49823 -107593
rect -49731 -107637 -49723 -107593
rect -49631 -107637 -49623 -107593
rect -49531 -107637 -49523 -107593
rect -49431 -107637 -49423 -107593
rect -49331 -107637 -49323 -107593
rect -49231 -107637 -49223 -107593
rect -49131 -107637 -49123 -107593
rect -49031 -107637 -49023 -107593
rect -48931 -107637 -48923 -107593
rect -48831 -107637 -48823 -107593
rect -48731 -107637 -48723 -107593
rect -48631 -107637 -48623 -107593
rect -48531 -107637 -48523 -107593
rect -48031 -107637 -48023 -107593
rect -47931 -107637 -47923 -107593
rect -47831 -107637 -47823 -107593
rect -47731 -107637 -47723 -107593
rect -47631 -107637 -47623 -107593
rect -47531 -107637 -47523 -107593
rect -47431 -107637 -47423 -107593
rect -47331 -107637 -47323 -107593
rect -47231 -107637 -47223 -107593
rect -47131 -107637 -47123 -107593
rect -47031 -107637 -47023 -107593
rect -46931 -107637 -46923 -107593
rect -46831 -107637 -46823 -107593
rect -46731 -107637 -46723 -107593
rect -46631 -107637 -46623 -107593
rect -46531 -107637 -46523 -107593
rect -46031 -107637 -46023 -107593
rect -45931 -107637 -45923 -107593
rect -45831 -107637 -45823 -107593
rect -45731 -107637 -45723 -107593
rect -45631 -107637 -45623 -107593
rect -45531 -107637 -45523 -107593
rect -45431 -107637 -45423 -107593
rect -45331 -107637 -45323 -107593
rect -45231 -107637 -45223 -107593
rect -45131 -107637 -45123 -107593
rect -45031 -107637 -45023 -107593
rect -44931 -107637 -44923 -107593
rect -44831 -107637 -44823 -107593
rect -44731 -107637 -44723 -107593
rect -44631 -107637 -44623 -107593
rect -44531 -107637 -44523 -107593
rect -44031 -107637 -44023 -107593
rect -43931 -107637 -43923 -107593
rect -43831 -107637 -43823 -107593
rect -43731 -107637 -43723 -107593
rect -43631 -107637 -43623 -107593
rect -43531 -107637 -43523 -107593
rect -43431 -107637 -43423 -107593
rect -43331 -107637 -43323 -107593
rect -43231 -107637 -43223 -107593
rect -43131 -107637 -43123 -107593
rect -43031 -107637 -43023 -107593
rect -42931 -107637 -42923 -107593
rect -42831 -107637 -42823 -107593
rect -42731 -107637 -42723 -107593
rect -42631 -107637 -42623 -107593
rect -42531 -107637 -42523 -107593
rect -50075 -107693 -50031 -107685
rect -49975 -107693 -49931 -107685
rect -49875 -107693 -49831 -107685
rect -49775 -107693 -49731 -107685
rect -49675 -107693 -49631 -107685
rect -49575 -107693 -49531 -107685
rect -49475 -107693 -49431 -107685
rect -49375 -107693 -49331 -107685
rect -49275 -107693 -49231 -107685
rect -49175 -107693 -49131 -107685
rect -49075 -107693 -49031 -107685
rect -48975 -107693 -48931 -107685
rect -48875 -107693 -48831 -107685
rect -48775 -107693 -48731 -107685
rect -48675 -107693 -48631 -107685
rect -48575 -107693 -48531 -107685
rect -48075 -107693 -48031 -107685
rect -47975 -107693 -47931 -107685
rect -47875 -107693 -47831 -107685
rect -47775 -107693 -47731 -107685
rect -47675 -107693 -47631 -107685
rect -47575 -107693 -47531 -107685
rect -47475 -107693 -47431 -107685
rect -47375 -107693 -47331 -107685
rect -47275 -107693 -47231 -107685
rect -47175 -107693 -47131 -107685
rect -47075 -107693 -47031 -107685
rect -46975 -107693 -46931 -107685
rect -46875 -107693 -46831 -107685
rect -46775 -107693 -46731 -107685
rect -46675 -107693 -46631 -107685
rect -46575 -107693 -46531 -107685
rect -46075 -107693 -46031 -107685
rect -45975 -107693 -45931 -107685
rect -45875 -107693 -45831 -107685
rect -45775 -107693 -45731 -107685
rect -45675 -107693 -45631 -107685
rect -45575 -107693 -45531 -107685
rect -45475 -107693 -45431 -107685
rect -45375 -107693 -45331 -107685
rect -45275 -107693 -45231 -107685
rect -45175 -107693 -45131 -107685
rect -45075 -107693 -45031 -107685
rect -44975 -107693 -44931 -107685
rect -44875 -107693 -44831 -107685
rect -44775 -107693 -44731 -107685
rect -44675 -107693 -44631 -107685
rect -44575 -107693 -44531 -107685
rect -44075 -107693 -44031 -107685
rect -43975 -107693 -43931 -107685
rect -43875 -107693 -43831 -107685
rect -43775 -107693 -43731 -107685
rect -43675 -107693 -43631 -107685
rect -43575 -107693 -43531 -107685
rect -43475 -107693 -43431 -107685
rect -43375 -107693 -43331 -107685
rect -43275 -107693 -43231 -107685
rect -43175 -107693 -43131 -107685
rect -43075 -107693 -43031 -107685
rect -42975 -107693 -42931 -107685
rect -42875 -107693 -42831 -107685
rect -42775 -107693 -42731 -107685
rect -42675 -107693 -42631 -107685
rect -42575 -107693 -42531 -107685
rect -50031 -107737 -50023 -107693
rect -49931 -107737 -49923 -107693
rect -49831 -107737 -49823 -107693
rect -49731 -107737 -49723 -107693
rect -49631 -107737 -49623 -107693
rect -49531 -107737 -49523 -107693
rect -49431 -107737 -49423 -107693
rect -49331 -107737 -49323 -107693
rect -49231 -107737 -49223 -107693
rect -49131 -107737 -49123 -107693
rect -49031 -107737 -49023 -107693
rect -48931 -107737 -48923 -107693
rect -48831 -107737 -48823 -107693
rect -48731 -107737 -48723 -107693
rect -48631 -107737 -48623 -107693
rect -48531 -107737 -48523 -107693
rect -48031 -107737 -48023 -107693
rect -47931 -107737 -47923 -107693
rect -47831 -107737 -47823 -107693
rect -47731 -107737 -47723 -107693
rect -47631 -107737 -47623 -107693
rect -47531 -107737 -47523 -107693
rect -47431 -107737 -47423 -107693
rect -47331 -107737 -47323 -107693
rect -47231 -107737 -47223 -107693
rect -47131 -107737 -47123 -107693
rect -47031 -107737 -47023 -107693
rect -46931 -107737 -46923 -107693
rect -46831 -107737 -46823 -107693
rect -46731 -107737 -46723 -107693
rect -46631 -107737 -46623 -107693
rect -46531 -107737 -46523 -107693
rect -46031 -107737 -46023 -107693
rect -45931 -107737 -45923 -107693
rect -45831 -107737 -45823 -107693
rect -45731 -107737 -45723 -107693
rect -45631 -107737 -45623 -107693
rect -45531 -107737 -45523 -107693
rect -45431 -107737 -45423 -107693
rect -45331 -107737 -45323 -107693
rect -45231 -107737 -45223 -107693
rect -45131 -107737 -45123 -107693
rect -45031 -107737 -45023 -107693
rect -44931 -107737 -44923 -107693
rect -44831 -107737 -44823 -107693
rect -44731 -107737 -44723 -107693
rect -44631 -107737 -44623 -107693
rect -44531 -107737 -44523 -107693
rect -44031 -107737 -44023 -107693
rect -43931 -107737 -43923 -107693
rect -43831 -107737 -43823 -107693
rect -43731 -107737 -43723 -107693
rect -43631 -107737 -43623 -107693
rect -43531 -107737 -43523 -107693
rect -43431 -107737 -43423 -107693
rect -43331 -107737 -43323 -107693
rect -43231 -107737 -43223 -107693
rect -43131 -107737 -43123 -107693
rect -43031 -107737 -43023 -107693
rect -42931 -107737 -42923 -107693
rect -42831 -107737 -42823 -107693
rect -42731 -107737 -42723 -107693
rect -42631 -107737 -42623 -107693
rect -42531 -107737 -42523 -107693
rect -109180 -129119 -109178 -109119
rect -109114 -129119 -109112 -109119
rect -77180 -129119 -77178 -109119
rect -77114 -129119 -77112 -109119
rect -45180 -129119 -45178 -109119
rect -45114 -129119 -45112 -109119
rect -13180 -129119 -13178 -109119
rect -13114 -129119 -13112 -109119
rect 18820 -129119 18822 -109119
rect 18886 -129119 18888 -109119
rect 50820 -129119 50822 -109119
rect 50886 -129119 50888 -109119
rect 82820 -129119 82822 -109119
rect 82886 -129119 82888 -109119
rect 114820 -129119 114822 -109119
rect 114886 -129119 114888 -109119
rect 146820 -129119 146822 -109119
rect 146886 -129119 146888 -109119
rect -13354 -131251 -13310 -131243
rect -13254 -131251 -13210 -131243
rect -13154 -131251 -13110 -131243
rect -13054 -131251 -13010 -131243
rect -12954 -131251 -12910 -131243
rect -12854 -131251 -12810 -131243
rect -12754 -131251 -12710 -131243
rect -12654 -131251 -12610 -131243
rect -12554 -131251 -12510 -131243
rect -12454 -131251 -12410 -131243
rect -12354 -131251 -12310 -131243
rect -12254 -131251 -12210 -131243
rect -12154 -131251 -12110 -131243
rect -12054 -131251 -12010 -131243
rect -11954 -131251 -11910 -131243
rect -11854 -131251 -11810 -131243
rect -11354 -131251 -11310 -131243
rect -11254 -131251 -11210 -131243
rect -11154 -131251 -11110 -131243
rect -11054 -131251 -11010 -131243
rect -10954 -131251 -10910 -131243
rect -10854 -131251 -10810 -131243
rect -10754 -131251 -10710 -131243
rect -10654 -131251 -10610 -131243
rect -10554 -131251 -10510 -131243
rect -10454 -131251 -10410 -131243
rect -10354 -131251 -10310 -131243
rect -10254 -131251 -10210 -131243
rect -10154 -131251 -10110 -131243
rect -10054 -131251 -10010 -131243
rect -9954 -131251 -9910 -131243
rect -9854 -131251 -9810 -131243
rect -9354 -131251 -9310 -131243
rect -9254 -131251 -9210 -131243
rect -9154 -131251 -9110 -131243
rect -9054 -131251 -9010 -131243
rect -8954 -131251 -8910 -131243
rect -8854 -131251 -8810 -131243
rect -8754 -131251 -8710 -131243
rect -8654 -131251 -8610 -131243
rect -8554 -131251 -8510 -131243
rect -8454 -131251 -8410 -131243
rect -8354 -131251 -8310 -131243
rect -8254 -131251 -8210 -131243
rect -8154 -131251 -8110 -131243
rect -8054 -131251 -8010 -131243
rect -7954 -131251 -7910 -131243
rect -7854 -131251 -7810 -131243
rect -7354 -131251 -7310 -131243
rect -7254 -131251 -7210 -131243
rect -7154 -131251 -7110 -131243
rect -7054 -131251 -7010 -131243
rect -6954 -131251 -6910 -131243
rect -6854 -131251 -6810 -131243
rect -6754 -131251 -6710 -131243
rect -6654 -131251 -6610 -131243
rect -6554 -131251 -6510 -131243
rect -6454 -131251 -6410 -131243
rect -6354 -131251 -6310 -131243
rect -6254 -131251 -6210 -131243
rect -6154 -131251 -6110 -131243
rect -6054 -131251 -6010 -131243
rect -5954 -131251 -5910 -131243
rect -5854 -131251 -5810 -131243
rect -13310 -131295 -13302 -131251
rect -13210 -131295 -13202 -131251
rect -13110 -131295 -13102 -131251
rect -13010 -131295 -13002 -131251
rect -12910 -131295 -12902 -131251
rect -12810 -131295 -12802 -131251
rect -12710 -131295 -12702 -131251
rect -12610 -131295 -12602 -131251
rect -12510 -131295 -12502 -131251
rect -12410 -131295 -12402 -131251
rect -12310 -131295 -12302 -131251
rect -12210 -131295 -12202 -131251
rect -12110 -131295 -12102 -131251
rect -12010 -131295 -12002 -131251
rect -11910 -131295 -11902 -131251
rect -11810 -131295 -11802 -131251
rect -11310 -131295 -11302 -131251
rect -11210 -131295 -11202 -131251
rect -11110 -131295 -11102 -131251
rect -11010 -131295 -11002 -131251
rect -10910 -131295 -10902 -131251
rect -10810 -131295 -10802 -131251
rect -10710 -131295 -10702 -131251
rect -10610 -131295 -10602 -131251
rect -10510 -131295 -10502 -131251
rect -10410 -131295 -10402 -131251
rect -10310 -131295 -10302 -131251
rect -10210 -131295 -10202 -131251
rect -10110 -131295 -10102 -131251
rect -10010 -131295 -10002 -131251
rect -9910 -131295 -9902 -131251
rect -9810 -131295 -9802 -131251
rect -9310 -131295 -9302 -131251
rect -9210 -131295 -9202 -131251
rect -9110 -131295 -9102 -131251
rect -9010 -131295 -9002 -131251
rect -8910 -131295 -8902 -131251
rect -8810 -131295 -8802 -131251
rect -8710 -131295 -8702 -131251
rect -8610 -131295 -8602 -131251
rect -8510 -131295 -8502 -131251
rect -8410 -131295 -8402 -131251
rect -8310 -131295 -8302 -131251
rect -8210 -131295 -8202 -131251
rect -8110 -131295 -8102 -131251
rect -8010 -131295 -8002 -131251
rect -7910 -131295 -7902 -131251
rect -7810 -131295 -7802 -131251
rect -7310 -131295 -7302 -131251
rect -7210 -131295 -7202 -131251
rect -7110 -131295 -7102 -131251
rect -7010 -131295 -7002 -131251
rect -6910 -131295 -6902 -131251
rect -6810 -131295 -6802 -131251
rect -6710 -131295 -6702 -131251
rect -6610 -131295 -6602 -131251
rect -6510 -131295 -6502 -131251
rect -6410 -131295 -6402 -131251
rect -6310 -131295 -6302 -131251
rect -6210 -131295 -6202 -131251
rect -6110 -131295 -6102 -131251
rect -6010 -131295 -6002 -131251
rect -5910 -131295 -5902 -131251
rect -5810 -131295 -5802 -131251
rect -13354 -131351 -13310 -131343
rect -13254 -131351 -13210 -131343
rect -13154 -131351 -13110 -131343
rect -13054 -131351 -13010 -131343
rect -12954 -131351 -12910 -131343
rect -12854 -131351 -12810 -131343
rect -12754 -131351 -12710 -131343
rect -12654 -131351 -12610 -131343
rect -12554 -131351 -12510 -131343
rect -12454 -131351 -12410 -131343
rect -12354 -131351 -12310 -131343
rect -12254 -131351 -12210 -131343
rect -12154 -131351 -12110 -131343
rect -12054 -131351 -12010 -131343
rect -11954 -131351 -11910 -131343
rect -11854 -131351 -11810 -131343
rect -11354 -131351 -11310 -131343
rect -11254 -131351 -11210 -131343
rect -11154 -131351 -11110 -131343
rect -11054 -131351 -11010 -131343
rect -10954 -131351 -10910 -131343
rect -10854 -131351 -10810 -131343
rect -10754 -131351 -10710 -131343
rect -10654 -131351 -10610 -131343
rect -10554 -131351 -10510 -131343
rect -10454 -131351 -10410 -131343
rect -10354 -131351 -10310 -131343
rect -10254 -131351 -10210 -131343
rect -10154 -131351 -10110 -131343
rect -10054 -131351 -10010 -131343
rect -9954 -131351 -9910 -131343
rect -9854 -131351 -9810 -131343
rect -9354 -131351 -9310 -131343
rect -9254 -131351 -9210 -131343
rect -9154 -131351 -9110 -131343
rect -9054 -131351 -9010 -131343
rect -8954 -131351 -8910 -131343
rect -8854 -131351 -8810 -131343
rect -8754 -131351 -8710 -131343
rect -8654 -131351 -8610 -131343
rect -8554 -131351 -8510 -131343
rect -8454 -131351 -8410 -131343
rect -8354 -131351 -8310 -131343
rect -8254 -131351 -8210 -131343
rect -8154 -131351 -8110 -131343
rect -8054 -131351 -8010 -131343
rect -7954 -131351 -7910 -131343
rect -7854 -131351 -7810 -131343
rect -7354 -131351 -7310 -131343
rect -7254 -131351 -7210 -131343
rect -7154 -131351 -7110 -131343
rect -7054 -131351 -7010 -131343
rect -6954 -131351 -6910 -131343
rect -6854 -131351 -6810 -131343
rect -6754 -131351 -6710 -131343
rect -6654 -131351 -6610 -131343
rect -6554 -131351 -6510 -131343
rect -6454 -131351 -6410 -131343
rect -6354 -131351 -6310 -131343
rect -6254 -131351 -6210 -131343
rect -6154 -131351 -6110 -131343
rect -6054 -131351 -6010 -131343
rect -5954 -131351 -5910 -131343
rect -5854 -131351 -5810 -131343
rect -13310 -131395 -13302 -131351
rect -13210 -131395 -13202 -131351
rect -13110 -131395 -13102 -131351
rect -13010 -131395 -13002 -131351
rect -12910 -131395 -12902 -131351
rect -12810 -131395 -12802 -131351
rect -12710 -131395 -12702 -131351
rect -12610 -131395 -12602 -131351
rect -12510 -131395 -12502 -131351
rect -12410 -131395 -12402 -131351
rect -12310 -131395 -12302 -131351
rect -12210 -131395 -12202 -131351
rect -12110 -131395 -12102 -131351
rect -12010 -131395 -12002 -131351
rect -11910 -131395 -11902 -131351
rect -11810 -131395 -11802 -131351
rect -11310 -131395 -11302 -131351
rect -11210 -131395 -11202 -131351
rect -11110 -131395 -11102 -131351
rect -11010 -131395 -11002 -131351
rect -10910 -131395 -10902 -131351
rect -10810 -131395 -10802 -131351
rect -10710 -131395 -10702 -131351
rect -10610 -131395 -10602 -131351
rect -10510 -131395 -10502 -131351
rect -10410 -131395 -10402 -131351
rect -10310 -131395 -10302 -131351
rect -10210 -131395 -10202 -131351
rect -10110 -131395 -10102 -131351
rect -10010 -131395 -10002 -131351
rect -9910 -131395 -9902 -131351
rect -9810 -131395 -9802 -131351
rect -9310 -131395 -9302 -131351
rect -9210 -131395 -9202 -131351
rect -9110 -131395 -9102 -131351
rect -9010 -131395 -9002 -131351
rect -8910 -131395 -8902 -131351
rect -8810 -131395 -8802 -131351
rect -8710 -131395 -8702 -131351
rect -8610 -131395 -8602 -131351
rect -8510 -131395 -8502 -131351
rect -8410 -131395 -8402 -131351
rect -8310 -131395 -8302 -131351
rect -8210 -131395 -8202 -131351
rect -8110 -131395 -8102 -131351
rect -8010 -131395 -8002 -131351
rect -7910 -131395 -7902 -131351
rect -7810 -131395 -7802 -131351
rect -7310 -131395 -7302 -131351
rect -7210 -131395 -7202 -131351
rect -7110 -131395 -7102 -131351
rect -7010 -131395 -7002 -131351
rect -6910 -131395 -6902 -131351
rect -6810 -131395 -6802 -131351
rect -6710 -131395 -6702 -131351
rect -6610 -131395 -6602 -131351
rect -6510 -131395 -6502 -131351
rect -6410 -131395 -6402 -131351
rect -6310 -131395 -6302 -131351
rect -6210 -131395 -6202 -131351
rect -6110 -131395 -6102 -131351
rect -6010 -131395 -6002 -131351
rect -5910 -131395 -5902 -131351
rect -5810 -131395 -5802 -131351
rect 37387 -131385 37431 -131377
rect 37487 -131385 37531 -131377
rect 37587 -131385 37631 -131377
rect 37687 -131385 37731 -131377
rect 37787 -131385 37831 -131377
rect 37887 -131385 37931 -131377
rect 37987 -131385 38031 -131377
rect 38087 -131385 38131 -131377
rect 38187 -131385 38231 -131377
rect 38287 -131385 38331 -131377
rect 38387 -131385 38431 -131377
rect 38487 -131385 38531 -131377
rect 38587 -131385 38631 -131377
rect 38687 -131385 38731 -131377
rect 38787 -131385 38831 -131377
rect 38887 -131385 38931 -131377
rect 39387 -131385 39431 -131377
rect 39487 -131385 39531 -131377
rect 39587 -131385 39631 -131377
rect 39687 -131385 39731 -131377
rect 39787 -131385 39831 -131377
rect 39887 -131385 39931 -131377
rect 39987 -131385 40031 -131377
rect 40087 -131385 40131 -131377
rect 40187 -131385 40231 -131377
rect 40287 -131385 40331 -131377
rect 40387 -131385 40431 -131377
rect 40487 -131385 40531 -131377
rect 40587 -131385 40631 -131377
rect 40687 -131385 40731 -131377
rect 40787 -131385 40831 -131377
rect 40887 -131385 40931 -131377
rect 41387 -131385 41431 -131377
rect 41487 -131385 41531 -131377
rect 41587 -131385 41631 -131377
rect 41687 -131385 41731 -131377
rect 41787 -131385 41831 -131377
rect 41887 -131385 41931 -131377
rect 41987 -131385 42031 -131377
rect 42087 -131385 42131 -131377
rect 42187 -131385 42231 -131377
rect 42287 -131385 42331 -131377
rect 42387 -131385 42431 -131377
rect 42487 -131385 42531 -131377
rect 42587 -131385 42631 -131377
rect 42687 -131385 42731 -131377
rect 42787 -131385 42831 -131377
rect 42887 -131385 42931 -131377
rect 43387 -131385 43431 -131377
rect 43487 -131385 43531 -131377
rect 43587 -131385 43631 -131377
rect 43687 -131385 43731 -131377
rect 43787 -131385 43831 -131377
rect 43887 -131385 43931 -131377
rect 43987 -131385 44031 -131377
rect 44087 -131385 44131 -131377
rect 44187 -131385 44231 -131377
rect 44287 -131385 44331 -131377
rect 44387 -131385 44431 -131377
rect 44487 -131385 44531 -131377
rect 44587 -131385 44631 -131377
rect 44687 -131385 44731 -131377
rect 44787 -131385 44831 -131377
rect 44887 -131385 44931 -131377
rect 37431 -131429 37439 -131385
rect 37531 -131429 37539 -131385
rect 37631 -131429 37639 -131385
rect 37731 -131429 37739 -131385
rect 37831 -131429 37839 -131385
rect 37931 -131429 37939 -131385
rect 38031 -131429 38039 -131385
rect 38131 -131429 38139 -131385
rect 38231 -131429 38239 -131385
rect 38331 -131429 38339 -131385
rect 38431 -131429 38439 -131385
rect 38531 -131429 38539 -131385
rect 38631 -131429 38639 -131385
rect 38731 -131429 38739 -131385
rect 38831 -131429 38839 -131385
rect 38931 -131429 38939 -131385
rect 39431 -131429 39439 -131385
rect 39531 -131429 39539 -131385
rect 39631 -131429 39639 -131385
rect 39731 -131429 39739 -131385
rect 39831 -131429 39839 -131385
rect 39931 -131429 39939 -131385
rect 40031 -131429 40039 -131385
rect 40131 -131429 40139 -131385
rect 40231 -131429 40239 -131385
rect 40331 -131429 40339 -131385
rect 40431 -131429 40439 -131385
rect 40531 -131429 40539 -131385
rect 40631 -131429 40639 -131385
rect 40731 -131429 40739 -131385
rect 40831 -131429 40839 -131385
rect 40931 -131429 40939 -131385
rect 41431 -131429 41439 -131385
rect 41531 -131429 41539 -131385
rect 41631 -131429 41639 -131385
rect 41731 -131429 41739 -131385
rect 41831 -131429 41839 -131385
rect 41931 -131429 41939 -131385
rect 42031 -131429 42039 -131385
rect 42131 -131429 42139 -131385
rect 42231 -131429 42239 -131385
rect 42331 -131429 42339 -131385
rect 42431 -131429 42439 -131385
rect 42531 -131429 42539 -131385
rect 42631 -131429 42639 -131385
rect 42731 -131429 42739 -131385
rect 42831 -131429 42839 -131385
rect 42931 -131429 42939 -131385
rect 43431 -131429 43439 -131385
rect 43531 -131429 43539 -131385
rect 43631 -131429 43639 -131385
rect 43731 -131429 43739 -131385
rect 43831 -131429 43839 -131385
rect 43931 -131429 43939 -131385
rect 44031 -131429 44039 -131385
rect 44131 -131429 44139 -131385
rect 44231 -131429 44239 -131385
rect 44331 -131429 44339 -131385
rect 44431 -131429 44439 -131385
rect 44531 -131429 44539 -131385
rect 44631 -131429 44639 -131385
rect 44731 -131429 44739 -131385
rect 44831 -131429 44839 -131385
rect 44931 -131429 44939 -131385
rect -13354 -131451 -13310 -131443
rect -13254 -131451 -13210 -131443
rect -13154 -131451 -13110 -131443
rect -13054 -131451 -13010 -131443
rect -12954 -131451 -12910 -131443
rect -12854 -131451 -12810 -131443
rect -12754 -131451 -12710 -131443
rect -12654 -131451 -12610 -131443
rect -12554 -131451 -12510 -131443
rect -12454 -131451 -12410 -131443
rect -12354 -131451 -12310 -131443
rect -12254 -131451 -12210 -131443
rect -12154 -131451 -12110 -131443
rect -12054 -131451 -12010 -131443
rect -11954 -131451 -11910 -131443
rect -11854 -131451 -11810 -131443
rect -11354 -131451 -11310 -131443
rect -11254 -131451 -11210 -131443
rect -11154 -131451 -11110 -131443
rect -11054 -131451 -11010 -131443
rect -10954 -131451 -10910 -131443
rect -10854 -131451 -10810 -131443
rect -10754 -131451 -10710 -131443
rect -10654 -131451 -10610 -131443
rect -10554 -131451 -10510 -131443
rect -10454 -131451 -10410 -131443
rect -10354 -131451 -10310 -131443
rect -10254 -131451 -10210 -131443
rect -10154 -131451 -10110 -131443
rect -10054 -131451 -10010 -131443
rect -9954 -131451 -9910 -131443
rect -9854 -131451 -9810 -131443
rect -9354 -131451 -9310 -131443
rect -9254 -131451 -9210 -131443
rect -9154 -131451 -9110 -131443
rect -9054 -131451 -9010 -131443
rect -8954 -131451 -8910 -131443
rect -8854 -131451 -8810 -131443
rect -8754 -131451 -8710 -131443
rect -8654 -131451 -8610 -131443
rect -8554 -131451 -8510 -131443
rect -8454 -131451 -8410 -131443
rect -8354 -131451 -8310 -131443
rect -8254 -131451 -8210 -131443
rect -8154 -131451 -8110 -131443
rect -8054 -131451 -8010 -131443
rect -7954 -131451 -7910 -131443
rect -7854 -131451 -7810 -131443
rect -7354 -131451 -7310 -131443
rect -7254 -131451 -7210 -131443
rect -7154 -131451 -7110 -131443
rect -7054 -131451 -7010 -131443
rect -6954 -131451 -6910 -131443
rect -6854 -131451 -6810 -131443
rect -6754 -131451 -6710 -131443
rect -6654 -131451 -6610 -131443
rect -6554 -131451 -6510 -131443
rect -6454 -131451 -6410 -131443
rect -6354 -131451 -6310 -131443
rect -6254 -131451 -6210 -131443
rect -6154 -131451 -6110 -131443
rect -6054 -131451 -6010 -131443
rect -5954 -131451 -5910 -131443
rect -5854 -131451 -5810 -131443
rect -13310 -131495 -13302 -131451
rect -13210 -131495 -13202 -131451
rect -13110 -131495 -13102 -131451
rect -13010 -131495 -13002 -131451
rect -12910 -131495 -12902 -131451
rect -12810 -131495 -12802 -131451
rect -12710 -131495 -12702 -131451
rect -12610 -131495 -12602 -131451
rect -12510 -131495 -12502 -131451
rect -12410 -131495 -12402 -131451
rect -12310 -131495 -12302 -131451
rect -12210 -131495 -12202 -131451
rect -12110 -131495 -12102 -131451
rect -12010 -131495 -12002 -131451
rect -11910 -131495 -11902 -131451
rect -11810 -131495 -11802 -131451
rect -11310 -131495 -11302 -131451
rect -11210 -131495 -11202 -131451
rect -11110 -131495 -11102 -131451
rect -11010 -131495 -11002 -131451
rect -10910 -131495 -10902 -131451
rect -10810 -131495 -10802 -131451
rect -10710 -131495 -10702 -131451
rect -10610 -131495 -10602 -131451
rect -10510 -131495 -10502 -131451
rect -10410 -131495 -10402 -131451
rect -10310 -131495 -10302 -131451
rect -10210 -131495 -10202 -131451
rect -10110 -131495 -10102 -131451
rect -10010 -131495 -10002 -131451
rect -9910 -131495 -9902 -131451
rect -9810 -131495 -9802 -131451
rect -9310 -131495 -9302 -131451
rect -9210 -131495 -9202 -131451
rect -9110 -131495 -9102 -131451
rect -9010 -131495 -9002 -131451
rect -8910 -131495 -8902 -131451
rect -8810 -131495 -8802 -131451
rect -8710 -131495 -8702 -131451
rect -8610 -131495 -8602 -131451
rect -8510 -131495 -8502 -131451
rect -8410 -131495 -8402 -131451
rect -8310 -131495 -8302 -131451
rect -8210 -131495 -8202 -131451
rect -8110 -131495 -8102 -131451
rect -8010 -131495 -8002 -131451
rect -7910 -131495 -7902 -131451
rect -7810 -131495 -7802 -131451
rect -7310 -131495 -7302 -131451
rect -7210 -131495 -7202 -131451
rect -7110 -131495 -7102 -131451
rect -7010 -131495 -7002 -131451
rect -6910 -131495 -6902 -131451
rect -6810 -131495 -6802 -131451
rect -6710 -131495 -6702 -131451
rect -6610 -131495 -6602 -131451
rect -6510 -131495 -6502 -131451
rect -6410 -131495 -6402 -131451
rect -6310 -131495 -6302 -131451
rect -6210 -131495 -6202 -131451
rect -6110 -131495 -6102 -131451
rect -6010 -131495 -6002 -131451
rect -5910 -131495 -5902 -131451
rect -5810 -131495 -5802 -131451
rect 37387 -131485 37431 -131477
rect 37487 -131485 37531 -131477
rect 37587 -131485 37631 -131477
rect 37687 -131485 37731 -131477
rect 37787 -131485 37831 -131477
rect 37887 -131485 37931 -131477
rect 37987 -131485 38031 -131477
rect 38087 -131485 38131 -131477
rect 38187 -131485 38231 -131477
rect 38287 -131485 38331 -131477
rect 38387 -131485 38431 -131477
rect 38487 -131485 38531 -131477
rect 38587 -131485 38631 -131477
rect 38687 -131485 38731 -131477
rect 38787 -131485 38831 -131477
rect 38887 -131485 38931 -131477
rect 39387 -131485 39431 -131477
rect 39487 -131485 39531 -131477
rect 39587 -131485 39631 -131477
rect 39687 -131485 39731 -131477
rect 39787 -131485 39831 -131477
rect 39887 -131485 39931 -131477
rect 39987 -131485 40031 -131477
rect 40087 -131485 40131 -131477
rect 40187 -131485 40231 -131477
rect 40287 -131485 40331 -131477
rect 40387 -131485 40431 -131477
rect 40487 -131485 40531 -131477
rect 40587 -131485 40631 -131477
rect 40687 -131485 40731 -131477
rect 40787 -131485 40831 -131477
rect 40887 -131485 40931 -131477
rect 41387 -131485 41431 -131477
rect 41487 -131485 41531 -131477
rect 41587 -131485 41631 -131477
rect 41687 -131485 41731 -131477
rect 41787 -131485 41831 -131477
rect 41887 -131485 41931 -131477
rect 41987 -131485 42031 -131477
rect 42087 -131485 42131 -131477
rect 42187 -131485 42231 -131477
rect 42287 -131485 42331 -131477
rect 42387 -131485 42431 -131477
rect 42487 -131485 42531 -131477
rect 42587 -131485 42631 -131477
rect 42687 -131485 42731 -131477
rect 42787 -131485 42831 -131477
rect 42887 -131485 42931 -131477
rect 43387 -131485 43431 -131477
rect 43487 -131485 43531 -131477
rect 43587 -131485 43631 -131477
rect 43687 -131485 43731 -131477
rect 43787 -131485 43831 -131477
rect 43887 -131485 43931 -131477
rect 43987 -131485 44031 -131477
rect 44087 -131485 44131 -131477
rect 44187 -131485 44231 -131477
rect 44287 -131485 44331 -131477
rect 44387 -131485 44431 -131477
rect 44487 -131485 44531 -131477
rect 44587 -131485 44631 -131477
rect 44687 -131485 44731 -131477
rect 44787 -131485 44831 -131477
rect 44887 -131485 44931 -131477
rect 37431 -131529 37439 -131485
rect 37531 -131529 37539 -131485
rect 37631 -131529 37639 -131485
rect 37731 -131529 37739 -131485
rect 37831 -131529 37839 -131485
rect 37931 -131529 37939 -131485
rect 38031 -131529 38039 -131485
rect 38131 -131529 38139 -131485
rect 38231 -131529 38239 -131485
rect 38331 -131529 38339 -131485
rect 38431 -131529 38439 -131485
rect 38531 -131529 38539 -131485
rect 38631 -131529 38639 -131485
rect 38731 -131529 38739 -131485
rect 38831 -131529 38839 -131485
rect 38931 -131529 38939 -131485
rect 39431 -131529 39439 -131485
rect 39531 -131529 39539 -131485
rect 39631 -131529 39639 -131485
rect 39731 -131529 39739 -131485
rect 39831 -131529 39839 -131485
rect 39931 -131529 39939 -131485
rect 40031 -131529 40039 -131485
rect 40131 -131529 40139 -131485
rect 40231 -131529 40239 -131485
rect 40331 -131529 40339 -131485
rect 40431 -131529 40439 -131485
rect 40531 -131529 40539 -131485
rect 40631 -131529 40639 -131485
rect 40731 -131529 40739 -131485
rect 40831 -131529 40839 -131485
rect 40931 -131529 40939 -131485
rect 41431 -131529 41439 -131485
rect 41531 -131529 41539 -131485
rect 41631 -131529 41639 -131485
rect 41731 -131529 41739 -131485
rect 41831 -131529 41839 -131485
rect 41931 -131529 41939 -131485
rect 42031 -131529 42039 -131485
rect 42131 -131529 42139 -131485
rect 42231 -131529 42239 -131485
rect 42331 -131529 42339 -131485
rect 42431 -131529 42439 -131485
rect 42531 -131529 42539 -131485
rect 42631 -131529 42639 -131485
rect 42731 -131529 42739 -131485
rect 42831 -131529 42839 -131485
rect 42931 -131529 42939 -131485
rect 43431 -131529 43439 -131485
rect 43531 -131529 43539 -131485
rect 43631 -131529 43639 -131485
rect 43731 -131529 43739 -131485
rect 43831 -131529 43839 -131485
rect 43931 -131529 43939 -131485
rect 44031 -131529 44039 -131485
rect 44131 -131529 44139 -131485
rect 44231 -131529 44239 -131485
rect 44331 -131529 44339 -131485
rect 44431 -131529 44439 -131485
rect 44531 -131529 44539 -131485
rect 44631 -131529 44639 -131485
rect 44731 -131529 44739 -131485
rect 44831 -131529 44839 -131485
rect 44931 -131529 44939 -131485
rect -13354 -131551 -13310 -131543
rect -13254 -131551 -13210 -131543
rect -13154 -131551 -13110 -131543
rect -13054 -131551 -13010 -131543
rect -12954 -131551 -12910 -131543
rect -12854 -131551 -12810 -131543
rect -12754 -131551 -12710 -131543
rect -12654 -131551 -12610 -131543
rect -12554 -131551 -12510 -131543
rect -12454 -131551 -12410 -131543
rect -12354 -131551 -12310 -131543
rect -12254 -131551 -12210 -131543
rect -12154 -131551 -12110 -131543
rect -12054 -131551 -12010 -131543
rect -11954 -131551 -11910 -131543
rect -11854 -131551 -11810 -131543
rect -11354 -131551 -11310 -131543
rect -11254 -131551 -11210 -131543
rect -11154 -131551 -11110 -131543
rect -11054 -131551 -11010 -131543
rect -10954 -131551 -10910 -131543
rect -10854 -131551 -10810 -131543
rect -10754 -131551 -10710 -131543
rect -10654 -131551 -10610 -131543
rect -10554 -131551 -10510 -131543
rect -10454 -131551 -10410 -131543
rect -10354 -131551 -10310 -131543
rect -10254 -131551 -10210 -131543
rect -10154 -131551 -10110 -131543
rect -10054 -131551 -10010 -131543
rect -9954 -131551 -9910 -131543
rect -9854 -131551 -9810 -131543
rect -9354 -131551 -9310 -131543
rect -9254 -131551 -9210 -131543
rect -9154 -131551 -9110 -131543
rect -9054 -131551 -9010 -131543
rect -8954 -131551 -8910 -131543
rect -8854 -131551 -8810 -131543
rect -8754 -131551 -8710 -131543
rect -8654 -131551 -8610 -131543
rect -8554 -131551 -8510 -131543
rect -8454 -131551 -8410 -131543
rect -8354 -131551 -8310 -131543
rect -8254 -131551 -8210 -131543
rect -8154 -131551 -8110 -131543
rect -8054 -131551 -8010 -131543
rect -7954 -131551 -7910 -131543
rect -7854 -131551 -7810 -131543
rect -7354 -131551 -7310 -131543
rect -7254 -131551 -7210 -131543
rect -7154 -131551 -7110 -131543
rect -7054 -131551 -7010 -131543
rect -6954 -131551 -6910 -131543
rect -6854 -131551 -6810 -131543
rect -6754 -131551 -6710 -131543
rect -6654 -131551 -6610 -131543
rect -6554 -131551 -6510 -131543
rect -6454 -131551 -6410 -131543
rect -6354 -131551 -6310 -131543
rect -6254 -131551 -6210 -131543
rect -6154 -131551 -6110 -131543
rect -6054 -131551 -6010 -131543
rect -5954 -131551 -5910 -131543
rect -5854 -131551 -5810 -131543
rect -13310 -131595 -13302 -131551
rect -13210 -131595 -13202 -131551
rect -13110 -131595 -13102 -131551
rect -13010 -131595 -13002 -131551
rect -12910 -131595 -12902 -131551
rect -12810 -131595 -12802 -131551
rect -12710 -131595 -12702 -131551
rect -12610 -131595 -12602 -131551
rect -12510 -131595 -12502 -131551
rect -12410 -131595 -12402 -131551
rect -12310 -131595 -12302 -131551
rect -12210 -131595 -12202 -131551
rect -12110 -131595 -12102 -131551
rect -12010 -131595 -12002 -131551
rect -11910 -131595 -11902 -131551
rect -11810 -131595 -11802 -131551
rect -11310 -131595 -11302 -131551
rect -11210 -131595 -11202 -131551
rect -11110 -131595 -11102 -131551
rect -11010 -131595 -11002 -131551
rect -10910 -131595 -10902 -131551
rect -10810 -131595 -10802 -131551
rect -10710 -131595 -10702 -131551
rect -10610 -131595 -10602 -131551
rect -10510 -131595 -10502 -131551
rect -10410 -131595 -10402 -131551
rect -10310 -131595 -10302 -131551
rect -10210 -131595 -10202 -131551
rect -10110 -131595 -10102 -131551
rect -10010 -131595 -10002 -131551
rect -9910 -131595 -9902 -131551
rect -9810 -131595 -9802 -131551
rect -9310 -131595 -9302 -131551
rect -9210 -131595 -9202 -131551
rect -9110 -131595 -9102 -131551
rect -9010 -131595 -9002 -131551
rect -8910 -131595 -8902 -131551
rect -8810 -131595 -8802 -131551
rect -8710 -131595 -8702 -131551
rect -8610 -131595 -8602 -131551
rect -8510 -131595 -8502 -131551
rect -8410 -131595 -8402 -131551
rect -8310 -131595 -8302 -131551
rect -8210 -131595 -8202 -131551
rect -8110 -131595 -8102 -131551
rect -8010 -131595 -8002 -131551
rect -7910 -131595 -7902 -131551
rect -7810 -131595 -7802 -131551
rect -7310 -131595 -7302 -131551
rect -7210 -131595 -7202 -131551
rect -7110 -131595 -7102 -131551
rect -7010 -131595 -7002 -131551
rect -6910 -131595 -6902 -131551
rect -6810 -131595 -6802 -131551
rect -6710 -131595 -6702 -131551
rect -6610 -131595 -6602 -131551
rect -6510 -131595 -6502 -131551
rect -6410 -131595 -6402 -131551
rect -6310 -131595 -6302 -131551
rect -6210 -131595 -6202 -131551
rect -6110 -131595 -6102 -131551
rect -6010 -131595 -6002 -131551
rect -5910 -131595 -5902 -131551
rect -5810 -131595 -5802 -131551
rect 37387 -131585 37431 -131577
rect 37487 -131585 37531 -131577
rect 37587 -131585 37631 -131577
rect 37687 -131585 37731 -131577
rect 37787 -131585 37831 -131577
rect 37887 -131585 37931 -131577
rect 37987 -131585 38031 -131577
rect 38087 -131585 38131 -131577
rect 38187 -131585 38231 -131577
rect 38287 -131585 38331 -131577
rect 38387 -131585 38431 -131577
rect 38487 -131585 38531 -131577
rect 38587 -131585 38631 -131577
rect 38687 -131585 38731 -131577
rect 38787 -131585 38831 -131577
rect 38887 -131585 38931 -131577
rect 39387 -131585 39431 -131577
rect 39487 -131585 39531 -131577
rect 39587 -131585 39631 -131577
rect 39687 -131585 39731 -131577
rect 39787 -131585 39831 -131577
rect 39887 -131585 39931 -131577
rect 39987 -131585 40031 -131577
rect 40087 -131585 40131 -131577
rect 40187 -131585 40231 -131577
rect 40287 -131585 40331 -131577
rect 40387 -131585 40431 -131577
rect 40487 -131585 40531 -131577
rect 40587 -131585 40631 -131577
rect 40687 -131585 40731 -131577
rect 40787 -131585 40831 -131577
rect 40887 -131585 40931 -131577
rect 41387 -131585 41431 -131577
rect 41487 -131585 41531 -131577
rect 41587 -131585 41631 -131577
rect 41687 -131585 41731 -131577
rect 41787 -131585 41831 -131577
rect 41887 -131585 41931 -131577
rect 41987 -131585 42031 -131577
rect 42087 -131585 42131 -131577
rect 42187 -131585 42231 -131577
rect 42287 -131585 42331 -131577
rect 42387 -131585 42431 -131577
rect 42487 -131585 42531 -131577
rect 42587 -131585 42631 -131577
rect 42687 -131585 42731 -131577
rect 42787 -131585 42831 -131577
rect 42887 -131585 42931 -131577
rect 43387 -131585 43431 -131577
rect 43487 -131585 43531 -131577
rect 43587 -131585 43631 -131577
rect 43687 -131585 43731 -131577
rect 43787 -131585 43831 -131577
rect 43887 -131585 43931 -131577
rect 43987 -131585 44031 -131577
rect 44087 -131585 44131 -131577
rect 44187 -131585 44231 -131577
rect 44287 -131585 44331 -131577
rect 44387 -131585 44431 -131577
rect 44487 -131585 44531 -131577
rect 44587 -131585 44631 -131577
rect 44687 -131585 44731 -131577
rect 44787 -131585 44831 -131577
rect 44887 -131585 44931 -131577
rect 37431 -131629 37439 -131585
rect 37531 -131629 37539 -131585
rect 37631 -131629 37639 -131585
rect 37731 -131629 37739 -131585
rect 37831 -131629 37839 -131585
rect 37931 -131629 37939 -131585
rect 38031 -131629 38039 -131585
rect 38131 -131629 38139 -131585
rect 38231 -131629 38239 -131585
rect 38331 -131629 38339 -131585
rect 38431 -131629 38439 -131585
rect 38531 -131629 38539 -131585
rect 38631 -131629 38639 -131585
rect 38731 -131629 38739 -131585
rect 38831 -131629 38839 -131585
rect 38931 -131629 38939 -131585
rect 39431 -131629 39439 -131585
rect 39531 -131629 39539 -131585
rect 39631 -131629 39639 -131585
rect 39731 -131629 39739 -131585
rect 39831 -131629 39839 -131585
rect 39931 -131629 39939 -131585
rect 40031 -131629 40039 -131585
rect 40131 -131629 40139 -131585
rect 40231 -131629 40239 -131585
rect 40331 -131629 40339 -131585
rect 40431 -131629 40439 -131585
rect 40531 -131629 40539 -131585
rect 40631 -131629 40639 -131585
rect 40731 -131629 40739 -131585
rect 40831 -131629 40839 -131585
rect 40931 -131629 40939 -131585
rect 41431 -131629 41439 -131585
rect 41531 -131629 41539 -131585
rect 41631 -131629 41639 -131585
rect 41731 -131629 41739 -131585
rect 41831 -131629 41839 -131585
rect 41931 -131629 41939 -131585
rect 42031 -131629 42039 -131585
rect 42131 -131629 42139 -131585
rect 42231 -131629 42239 -131585
rect 42331 -131629 42339 -131585
rect 42431 -131629 42439 -131585
rect 42531 -131629 42539 -131585
rect 42631 -131629 42639 -131585
rect 42731 -131629 42739 -131585
rect 42831 -131629 42839 -131585
rect 42931 -131629 42939 -131585
rect 43431 -131629 43439 -131585
rect 43531 -131629 43539 -131585
rect 43631 -131629 43639 -131585
rect 43731 -131629 43739 -131585
rect 43831 -131629 43839 -131585
rect 43931 -131629 43939 -131585
rect 44031 -131629 44039 -131585
rect 44131 -131629 44139 -131585
rect 44231 -131629 44239 -131585
rect 44331 -131629 44339 -131585
rect 44431 -131629 44439 -131585
rect 44531 -131629 44539 -131585
rect 44631 -131629 44639 -131585
rect 44731 -131629 44739 -131585
rect 44831 -131629 44839 -131585
rect 44931 -131629 44939 -131585
rect -13354 -131651 -13310 -131643
rect -13254 -131651 -13210 -131643
rect -13154 -131651 -13110 -131643
rect -13054 -131651 -13010 -131643
rect -12954 -131651 -12910 -131643
rect -12854 -131651 -12810 -131643
rect -12754 -131651 -12710 -131643
rect -12654 -131651 -12610 -131643
rect -12554 -131651 -12510 -131643
rect -12454 -131651 -12410 -131643
rect -12354 -131651 -12310 -131643
rect -12254 -131651 -12210 -131643
rect -12154 -131651 -12110 -131643
rect -12054 -131651 -12010 -131643
rect -11954 -131651 -11910 -131643
rect -11854 -131651 -11810 -131643
rect -11354 -131651 -11310 -131643
rect -11254 -131651 -11210 -131643
rect -11154 -131651 -11110 -131643
rect -11054 -131651 -11010 -131643
rect -10954 -131651 -10910 -131643
rect -10854 -131651 -10810 -131643
rect -10754 -131651 -10710 -131643
rect -10654 -131651 -10610 -131643
rect -10554 -131651 -10510 -131643
rect -10454 -131651 -10410 -131643
rect -10354 -131651 -10310 -131643
rect -10254 -131651 -10210 -131643
rect -10154 -131651 -10110 -131643
rect -10054 -131651 -10010 -131643
rect -9954 -131651 -9910 -131643
rect -9854 -131651 -9810 -131643
rect -9354 -131651 -9310 -131643
rect -9254 -131651 -9210 -131643
rect -9154 -131651 -9110 -131643
rect -9054 -131651 -9010 -131643
rect -8954 -131651 -8910 -131643
rect -8854 -131651 -8810 -131643
rect -8754 -131651 -8710 -131643
rect -8654 -131651 -8610 -131643
rect -8554 -131651 -8510 -131643
rect -8454 -131651 -8410 -131643
rect -8354 -131651 -8310 -131643
rect -8254 -131651 -8210 -131643
rect -8154 -131651 -8110 -131643
rect -8054 -131651 -8010 -131643
rect -7954 -131651 -7910 -131643
rect -7854 -131651 -7810 -131643
rect -7354 -131651 -7310 -131643
rect -7254 -131651 -7210 -131643
rect -7154 -131651 -7110 -131643
rect -7054 -131651 -7010 -131643
rect -6954 -131651 -6910 -131643
rect -6854 -131651 -6810 -131643
rect -6754 -131651 -6710 -131643
rect -6654 -131651 -6610 -131643
rect -6554 -131651 -6510 -131643
rect -6454 -131651 -6410 -131643
rect -6354 -131651 -6310 -131643
rect -6254 -131651 -6210 -131643
rect -6154 -131651 -6110 -131643
rect -6054 -131651 -6010 -131643
rect -5954 -131651 -5910 -131643
rect -5854 -131651 -5810 -131643
rect -13310 -131695 -13302 -131651
rect -13210 -131695 -13202 -131651
rect -13110 -131695 -13102 -131651
rect -13010 -131695 -13002 -131651
rect -12910 -131695 -12902 -131651
rect -12810 -131695 -12802 -131651
rect -12710 -131695 -12702 -131651
rect -12610 -131695 -12602 -131651
rect -12510 -131695 -12502 -131651
rect -12410 -131695 -12402 -131651
rect -12310 -131695 -12302 -131651
rect -12210 -131695 -12202 -131651
rect -12110 -131695 -12102 -131651
rect -12010 -131695 -12002 -131651
rect -11910 -131695 -11902 -131651
rect -11810 -131695 -11802 -131651
rect -11310 -131695 -11302 -131651
rect -11210 -131695 -11202 -131651
rect -11110 -131695 -11102 -131651
rect -11010 -131695 -11002 -131651
rect -10910 -131695 -10902 -131651
rect -10810 -131695 -10802 -131651
rect -10710 -131695 -10702 -131651
rect -10610 -131695 -10602 -131651
rect -10510 -131695 -10502 -131651
rect -10410 -131695 -10402 -131651
rect -10310 -131695 -10302 -131651
rect -10210 -131695 -10202 -131651
rect -10110 -131695 -10102 -131651
rect -10010 -131695 -10002 -131651
rect -9910 -131695 -9902 -131651
rect -9810 -131695 -9802 -131651
rect -9310 -131695 -9302 -131651
rect -9210 -131695 -9202 -131651
rect -9110 -131695 -9102 -131651
rect -9010 -131695 -9002 -131651
rect -8910 -131695 -8902 -131651
rect -8810 -131695 -8802 -131651
rect -8710 -131695 -8702 -131651
rect -8610 -131695 -8602 -131651
rect -8510 -131695 -8502 -131651
rect -8410 -131695 -8402 -131651
rect -8310 -131695 -8302 -131651
rect -8210 -131695 -8202 -131651
rect -8110 -131695 -8102 -131651
rect -8010 -131695 -8002 -131651
rect -7910 -131695 -7902 -131651
rect -7810 -131695 -7802 -131651
rect -7310 -131695 -7302 -131651
rect -7210 -131695 -7202 -131651
rect -7110 -131695 -7102 -131651
rect -7010 -131695 -7002 -131651
rect -6910 -131695 -6902 -131651
rect -6810 -131695 -6802 -131651
rect -6710 -131695 -6702 -131651
rect -6610 -131695 -6602 -131651
rect -6510 -131695 -6502 -131651
rect -6410 -131695 -6402 -131651
rect -6310 -131695 -6302 -131651
rect -6210 -131695 -6202 -131651
rect -6110 -131695 -6102 -131651
rect -6010 -131695 -6002 -131651
rect -5910 -131695 -5902 -131651
rect -5810 -131695 -5802 -131651
rect 37387 -131685 37431 -131677
rect 37487 -131685 37531 -131677
rect 37587 -131685 37631 -131677
rect 37687 -131685 37731 -131677
rect 37787 -131685 37831 -131677
rect 37887 -131685 37931 -131677
rect 37987 -131685 38031 -131677
rect 38087 -131685 38131 -131677
rect 38187 -131685 38231 -131677
rect 38287 -131685 38331 -131677
rect 38387 -131685 38431 -131677
rect 38487 -131685 38531 -131677
rect 38587 -131685 38631 -131677
rect 38687 -131685 38731 -131677
rect 38787 -131685 38831 -131677
rect 38887 -131685 38931 -131677
rect 39387 -131685 39431 -131677
rect 39487 -131685 39531 -131677
rect 39587 -131685 39631 -131677
rect 39687 -131685 39731 -131677
rect 39787 -131685 39831 -131677
rect 39887 -131685 39931 -131677
rect 39987 -131685 40031 -131677
rect 40087 -131685 40131 -131677
rect 40187 -131685 40231 -131677
rect 40287 -131685 40331 -131677
rect 40387 -131685 40431 -131677
rect 40487 -131685 40531 -131677
rect 40587 -131685 40631 -131677
rect 40687 -131685 40731 -131677
rect 40787 -131685 40831 -131677
rect 40887 -131685 40931 -131677
rect 41387 -131685 41431 -131677
rect 41487 -131685 41531 -131677
rect 41587 -131685 41631 -131677
rect 41687 -131685 41731 -131677
rect 41787 -131685 41831 -131677
rect 41887 -131685 41931 -131677
rect 41987 -131685 42031 -131677
rect 42087 -131685 42131 -131677
rect 42187 -131685 42231 -131677
rect 42287 -131685 42331 -131677
rect 42387 -131685 42431 -131677
rect 42487 -131685 42531 -131677
rect 42587 -131685 42631 -131677
rect 42687 -131685 42731 -131677
rect 42787 -131685 42831 -131677
rect 42887 -131685 42931 -131677
rect 43387 -131685 43431 -131677
rect 43487 -131685 43531 -131677
rect 43587 -131685 43631 -131677
rect 43687 -131685 43731 -131677
rect 43787 -131685 43831 -131677
rect 43887 -131685 43931 -131677
rect 43987 -131685 44031 -131677
rect 44087 -131685 44131 -131677
rect 44187 -131685 44231 -131677
rect 44287 -131685 44331 -131677
rect 44387 -131685 44431 -131677
rect 44487 -131685 44531 -131677
rect 44587 -131685 44631 -131677
rect 44687 -131685 44731 -131677
rect 44787 -131685 44831 -131677
rect 44887 -131685 44931 -131677
rect 37431 -131729 37439 -131685
rect 37531 -131729 37539 -131685
rect 37631 -131729 37639 -131685
rect 37731 -131729 37739 -131685
rect 37831 -131729 37839 -131685
rect 37931 -131729 37939 -131685
rect 38031 -131729 38039 -131685
rect 38131 -131729 38139 -131685
rect 38231 -131729 38239 -131685
rect 38331 -131729 38339 -131685
rect 38431 -131729 38439 -131685
rect 38531 -131729 38539 -131685
rect 38631 -131729 38639 -131685
rect 38731 -131729 38739 -131685
rect 38831 -131729 38839 -131685
rect 38931 -131729 38939 -131685
rect 39431 -131729 39439 -131685
rect 39531 -131729 39539 -131685
rect 39631 -131729 39639 -131685
rect 39731 -131729 39739 -131685
rect 39831 -131729 39839 -131685
rect 39931 -131729 39939 -131685
rect 40031 -131729 40039 -131685
rect 40131 -131729 40139 -131685
rect 40231 -131729 40239 -131685
rect 40331 -131729 40339 -131685
rect 40431 -131729 40439 -131685
rect 40531 -131729 40539 -131685
rect 40631 -131729 40639 -131685
rect 40731 -131729 40739 -131685
rect 40831 -131729 40839 -131685
rect 40931 -131729 40939 -131685
rect 41431 -131729 41439 -131685
rect 41531 -131729 41539 -131685
rect 41631 -131729 41639 -131685
rect 41731 -131729 41739 -131685
rect 41831 -131729 41839 -131685
rect 41931 -131729 41939 -131685
rect 42031 -131729 42039 -131685
rect 42131 -131729 42139 -131685
rect 42231 -131729 42239 -131685
rect 42331 -131729 42339 -131685
rect 42431 -131729 42439 -131685
rect 42531 -131729 42539 -131685
rect 42631 -131729 42639 -131685
rect 42731 -131729 42739 -131685
rect 42831 -131729 42839 -131685
rect 42931 -131729 42939 -131685
rect 43431 -131729 43439 -131685
rect 43531 -131729 43539 -131685
rect 43631 -131729 43639 -131685
rect 43731 -131729 43739 -131685
rect 43831 -131729 43839 -131685
rect 43931 -131729 43939 -131685
rect 44031 -131729 44039 -131685
rect 44131 -131729 44139 -131685
rect 44231 -131729 44239 -131685
rect 44331 -131729 44339 -131685
rect 44431 -131729 44439 -131685
rect 44531 -131729 44539 -131685
rect 44631 -131729 44639 -131685
rect 44731 -131729 44739 -131685
rect 44831 -131729 44839 -131685
rect 44931 -131729 44939 -131685
rect -13354 -131751 -13310 -131743
rect -13254 -131751 -13210 -131743
rect -13154 -131751 -13110 -131743
rect -13054 -131751 -13010 -131743
rect -12954 -131751 -12910 -131743
rect -12854 -131751 -12810 -131743
rect -12754 -131751 -12710 -131743
rect -12654 -131751 -12610 -131743
rect -12554 -131751 -12510 -131743
rect -12454 -131751 -12410 -131743
rect -12354 -131751 -12310 -131743
rect -12254 -131751 -12210 -131743
rect -12154 -131751 -12110 -131743
rect -12054 -131751 -12010 -131743
rect -11954 -131751 -11910 -131743
rect -11854 -131751 -11810 -131743
rect -11354 -131751 -11310 -131743
rect -11254 -131751 -11210 -131743
rect -11154 -131751 -11110 -131743
rect -11054 -131751 -11010 -131743
rect -10954 -131751 -10910 -131743
rect -10854 -131751 -10810 -131743
rect -10754 -131751 -10710 -131743
rect -10654 -131751 -10610 -131743
rect -10554 -131751 -10510 -131743
rect -10454 -131751 -10410 -131743
rect -10354 -131751 -10310 -131743
rect -10254 -131751 -10210 -131743
rect -10154 -131751 -10110 -131743
rect -10054 -131751 -10010 -131743
rect -9954 -131751 -9910 -131743
rect -9854 -131751 -9810 -131743
rect -9354 -131751 -9310 -131743
rect -9254 -131751 -9210 -131743
rect -9154 -131751 -9110 -131743
rect -9054 -131751 -9010 -131743
rect -8954 -131751 -8910 -131743
rect -8854 -131751 -8810 -131743
rect -8754 -131751 -8710 -131743
rect -8654 -131751 -8610 -131743
rect -8554 -131751 -8510 -131743
rect -8454 -131751 -8410 -131743
rect -8354 -131751 -8310 -131743
rect -8254 -131751 -8210 -131743
rect -8154 -131751 -8110 -131743
rect -8054 -131751 -8010 -131743
rect -7954 -131751 -7910 -131743
rect -7854 -131751 -7810 -131743
rect -7354 -131751 -7310 -131743
rect -7254 -131751 -7210 -131743
rect -7154 -131751 -7110 -131743
rect -7054 -131751 -7010 -131743
rect -6954 -131751 -6910 -131743
rect -6854 -131751 -6810 -131743
rect -6754 -131751 -6710 -131743
rect -6654 -131751 -6610 -131743
rect -6554 -131751 -6510 -131743
rect -6454 -131751 -6410 -131743
rect -6354 -131751 -6310 -131743
rect -6254 -131751 -6210 -131743
rect -6154 -131751 -6110 -131743
rect -6054 -131751 -6010 -131743
rect -5954 -131751 -5910 -131743
rect -5854 -131751 -5810 -131743
rect -13310 -131795 -13302 -131751
rect -13210 -131795 -13202 -131751
rect -13110 -131795 -13102 -131751
rect -13010 -131795 -13002 -131751
rect -12910 -131795 -12902 -131751
rect -12810 -131795 -12802 -131751
rect -12710 -131795 -12702 -131751
rect -12610 -131795 -12602 -131751
rect -12510 -131795 -12502 -131751
rect -12410 -131795 -12402 -131751
rect -12310 -131795 -12302 -131751
rect -12210 -131795 -12202 -131751
rect -12110 -131795 -12102 -131751
rect -12010 -131795 -12002 -131751
rect -11910 -131795 -11902 -131751
rect -11810 -131795 -11802 -131751
rect -11310 -131795 -11302 -131751
rect -11210 -131795 -11202 -131751
rect -11110 -131795 -11102 -131751
rect -11010 -131795 -11002 -131751
rect -10910 -131795 -10902 -131751
rect -10810 -131795 -10802 -131751
rect -10710 -131795 -10702 -131751
rect -10610 -131795 -10602 -131751
rect -10510 -131795 -10502 -131751
rect -10410 -131795 -10402 -131751
rect -10310 -131795 -10302 -131751
rect -10210 -131795 -10202 -131751
rect -10110 -131795 -10102 -131751
rect -10010 -131795 -10002 -131751
rect -9910 -131795 -9902 -131751
rect -9810 -131795 -9802 -131751
rect -9310 -131795 -9302 -131751
rect -9210 -131795 -9202 -131751
rect -9110 -131795 -9102 -131751
rect -9010 -131795 -9002 -131751
rect -8910 -131795 -8902 -131751
rect -8810 -131795 -8802 -131751
rect -8710 -131795 -8702 -131751
rect -8610 -131795 -8602 -131751
rect -8510 -131795 -8502 -131751
rect -8410 -131795 -8402 -131751
rect -8310 -131795 -8302 -131751
rect -8210 -131795 -8202 -131751
rect -8110 -131795 -8102 -131751
rect -8010 -131795 -8002 -131751
rect -7910 -131795 -7902 -131751
rect -7810 -131795 -7802 -131751
rect -7310 -131795 -7302 -131751
rect -7210 -131795 -7202 -131751
rect -7110 -131795 -7102 -131751
rect -7010 -131795 -7002 -131751
rect -6910 -131795 -6902 -131751
rect -6810 -131795 -6802 -131751
rect -6710 -131795 -6702 -131751
rect -6610 -131795 -6602 -131751
rect -6510 -131795 -6502 -131751
rect -6410 -131795 -6402 -131751
rect -6310 -131795 -6302 -131751
rect -6210 -131795 -6202 -131751
rect -6110 -131795 -6102 -131751
rect -6010 -131795 -6002 -131751
rect -5910 -131795 -5902 -131751
rect -5810 -131795 -5802 -131751
rect 37387 -131785 37431 -131777
rect 37487 -131785 37531 -131777
rect 37587 -131785 37631 -131777
rect 37687 -131785 37731 -131777
rect 37787 -131785 37831 -131777
rect 37887 -131785 37931 -131777
rect 37987 -131785 38031 -131777
rect 38087 -131785 38131 -131777
rect 38187 -131785 38231 -131777
rect 38287 -131785 38331 -131777
rect 38387 -131785 38431 -131777
rect 38487 -131785 38531 -131777
rect 38587 -131785 38631 -131777
rect 38687 -131785 38731 -131777
rect 38787 -131785 38831 -131777
rect 38887 -131785 38931 -131777
rect 39387 -131785 39431 -131777
rect 39487 -131785 39531 -131777
rect 39587 -131785 39631 -131777
rect 39687 -131785 39731 -131777
rect 39787 -131785 39831 -131777
rect 39887 -131785 39931 -131777
rect 39987 -131785 40031 -131777
rect 40087 -131785 40131 -131777
rect 40187 -131785 40231 -131777
rect 40287 -131785 40331 -131777
rect 40387 -131785 40431 -131777
rect 40487 -131785 40531 -131777
rect 40587 -131785 40631 -131777
rect 40687 -131785 40731 -131777
rect 40787 -131785 40831 -131777
rect 40887 -131785 40931 -131777
rect 41387 -131785 41431 -131777
rect 41487 -131785 41531 -131777
rect 41587 -131785 41631 -131777
rect 41687 -131785 41731 -131777
rect 41787 -131785 41831 -131777
rect 41887 -131785 41931 -131777
rect 41987 -131785 42031 -131777
rect 42087 -131785 42131 -131777
rect 42187 -131785 42231 -131777
rect 42287 -131785 42331 -131777
rect 42387 -131785 42431 -131777
rect 42487 -131785 42531 -131777
rect 42587 -131785 42631 -131777
rect 42687 -131785 42731 -131777
rect 42787 -131785 42831 -131777
rect 42887 -131785 42931 -131777
rect 43387 -131785 43431 -131777
rect 43487 -131785 43531 -131777
rect 43587 -131785 43631 -131777
rect 43687 -131785 43731 -131777
rect 43787 -131785 43831 -131777
rect 43887 -131785 43931 -131777
rect 43987 -131785 44031 -131777
rect 44087 -131785 44131 -131777
rect 44187 -131785 44231 -131777
rect 44287 -131785 44331 -131777
rect 44387 -131785 44431 -131777
rect 44487 -131785 44531 -131777
rect 44587 -131785 44631 -131777
rect 44687 -131785 44731 -131777
rect 44787 -131785 44831 -131777
rect 44887 -131785 44931 -131777
rect 37431 -131829 37439 -131785
rect 37531 -131829 37539 -131785
rect 37631 -131829 37639 -131785
rect 37731 -131829 37739 -131785
rect 37831 -131829 37839 -131785
rect 37931 -131829 37939 -131785
rect 38031 -131829 38039 -131785
rect 38131 -131829 38139 -131785
rect 38231 -131829 38239 -131785
rect 38331 -131829 38339 -131785
rect 38431 -131829 38439 -131785
rect 38531 -131829 38539 -131785
rect 38631 -131829 38639 -131785
rect 38731 -131829 38739 -131785
rect 38831 -131829 38839 -131785
rect 38931 -131829 38939 -131785
rect 39431 -131829 39439 -131785
rect 39531 -131829 39539 -131785
rect 39631 -131829 39639 -131785
rect 39731 -131829 39739 -131785
rect 39831 -131829 39839 -131785
rect 39931 -131829 39939 -131785
rect 40031 -131829 40039 -131785
rect 40131 -131829 40139 -131785
rect 40231 -131829 40239 -131785
rect 40331 -131829 40339 -131785
rect 40431 -131829 40439 -131785
rect 40531 -131829 40539 -131785
rect 40631 -131829 40639 -131785
rect 40731 -131829 40739 -131785
rect 40831 -131829 40839 -131785
rect 40931 -131829 40939 -131785
rect 41431 -131829 41439 -131785
rect 41531 -131829 41539 -131785
rect 41631 -131829 41639 -131785
rect 41731 -131829 41739 -131785
rect 41831 -131829 41839 -131785
rect 41931 -131829 41939 -131785
rect 42031 -131829 42039 -131785
rect 42131 -131829 42139 -131785
rect 42231 -131829 42239 -131785
rect 42331 -131829 42339 -131785
rect 42431 -131829 42439 -131785
rect 42531 -131829 42539 -131785
rect 42631 -131829 42639 -131785
rect 42731 -131829 42739 -131785
rect 42831 -131829 42839 -131785
rect 42931 -131829 42939 -131785
rect 43431 -131829 43439 -131785
rect 43531 -131829 43539 -131785
rect 43631 -131829 43639 -131785
rect 43731 -131829 43739 -131785
rect 43831 -131829 43839 -131785
rect 43931 -131829 43939 -131785
rect 44031 -131829 44039 -131785
rect 44131 -131829 44139 -131785
rect 44231 -131829 44239 -131785
rect 44331 -131829 44339 -131785
rect 44431 -131829 44439 -131785
rect 44531 -131829 44539 -131785
rect 44631 -131829 44639 -131785
rect 44731 -131829 44739 -131785
rect 44831 -131829 44839 -131785
rect 44931 -131829 44939 -131785
rect -13354 -131851 -13310 -131843
rect -13254 -131851 -13210 -131843
rect -13154 -131851 -13110 -131843
rect -13054 -131851 -13010 -131843
rect -12954 -131851 -12910 -131843
rect -12854 -131851 -12810 -131843
rect -12754 -131851 -12710 -131843
rect -12654 -131851 -12610 -131843
rect -12554 -131851 -12510 -131843
rect -12454 -131851 -12410 -131843
rect -12354 -131851 -12310 -131843
rect -12254 -131851 -12210 -131843
rect -12154 -131851 -12110 -131843
rect -12054 -131851 -12010 -131843
rect -11954 -131851 -11910 -131843
rect -11854 -131851 -11810 -131843
rect -11354 -131851 -11310 -131843
rect -11254 -131851 -11210 -131843
rect -11154 -131851 -11110 -131843
rect -11054 -131851 -11010 -131843
rect -10954 -131851 -10910 -131843
rect -10854 -131851 -10810 -131843
rect -10754 -131851 -10710 -131843
rect -10654 -131851 -10610 -131843
rect -10554 -131851 -10510 -131843
rect -10454 -131851 -10410 -131843
rect -10354 -131851 -10310 -131843
rect -10254 -131851 -10210 -131843
rect -10154 -131851 -10110 -131843
rect -10054 -131851 -10010 -131843
rect -9954 -131851 -9910 -131843
rect -9854 -131851 -9810 -131843
rect -9354 -131851 -9310 -131843
rect -9254 -131851 -9210 -131843
rect -9154 -131851 -9110 -131843
rect -9054 -131851 -9010 -131843
rect -8954 -131851 -8910 -131843
rect -8854 -131851 -8810 -131843
rect -8754 -131851 -8710 -131843
rect -8654 -131851 -8610 -131843
rect -8554 -131851 -8510 -131843
rect -8454 -131851 -8410 -131843
rect -8354 -131851 -8310 -131843
rect -8254 -131851 -8210 -131843
rect -8154 -131851 -8110 -131843
rect -8054 -131851 -8010 -131843
rect -7954 -131851 -7910 -131843
rect -7854 -131851 -7810 -131843
rect -7354 -131851 -7310 -131843
rect -7254 -131851 -7210 -131843
rect -7154 -131851 -7110 -131843
rect -7054 -131851 -7010 -131843
rect -6954 -131851 -6910 -131843
rect -6854 -131851 -6810 -131843
rect -6754 -131851 -6710 -131843
rect -6654 -131851 -6610 -131843
rect -6554 -131851 -6510 -131843
rect -6454 -131851 -6410 -131843
rect -6354 -131851 -6310 -131843
rect -6254 -131851 -6210 -131843
rect -6154 -131851 -6110 -131843
rect -6054 -131851 -6010 -131843
rect -5954 -131851 -5910 -131843
rect -5854 -131851 -5810 -131843
rect -13310 -131895 -13302 -131851
rect -13210 -131895 -13202 -131851
rect -13110 -131895 -13102 -131851
rect -13010 -131895 -13002 -131851
rect -12910 -131895 -12902 -131851
rect -12810 -131895 -12802 -131851
rect -12710 -131895 -12702 -131851
rect -12610 -131895 -12602 -131851
rect -12510 -131895 -12502 -131851
rect -12410 -131895 -12402 -131851
rect -12310 -131895 -12302 -131851
rect -12210 -131895 -12202 -131851
rect -12110 -131895 -12102 -131851
rect -12010 -131895 -12002 -131851
rect -11910 -131895 -11902 -131851
rect -11810 -131895 -11802 -131851
rect -11310 -131895 -11302 -131851
rect -11210 -131895 -11202 -131851
rect -11110 -131895 -11102 -131851
rect -11010 -131895 -11002 -131851
rect -10910 -131895 -10902 -131851
rect -10810 -131895 -10802 -131851
rect -10710 -131895 -10702 -131851
rect -10610 -131895 -10602 -131851
rect -10510 -131895 -10502 -131851
rect -10410 -131895 -10402 -131851
rect -10310 -131895 -10302 -131851
rect -10210 -131895 -10202 -131851
rect -10110 -131895 -10102 -131851
rect -10010 -131895 -10002 -131851
rect -9910 -131895 -9902 -131851
rect -9810 -131895 -9802 -131851
rect -9310 -131895 -9302 -131851
rect -9210 -131895 -9202 -131851
rect -9110 -131895 -9102 -131851
rect -9010 -131895 -9002 -131851
rect -8910 -131895 -8902 -131851
rect -8810 -131895 -8802 -131851
rect -8710 -131895 -8702 -131851
rect -8610 -131895 -8602 -131851
rect -8510 -131895 -8502 -131851
rect -8410 -131895 -8402 -131851
rect -8310 -131895 -8302 -131851
rect -8210 -131895 -8202 -131851
rect -8110 -131895 -8102 -131851
rect -8010 -131895 -8002 -131851
rect -7910 -131895 -7902 -131851
rect -7810 -131895 -7802 -131851
rect -7310 -131895 -7302 -131851
rect -7210 -131895 -7202 -131851
rect -7110 -131895 -7102 -131851
rect -7010 -131895 -7002 -131851
rect -6910 -131895 -6902 -131851
rect -6810 -131895 -6802 -131851
rect -6710 -131895 -6702 -131851
rect -6610 -131895 -6602 -131851
rect -6510 -131895 -6502 -131851
rect -6410 -131895 -6402 -131851
rect -6310 -131895 -6302 -131851
rect -6210 -131895 -6202 -131851
rect -6110 -131895 -6102 -131851
rect -6010 -131895 -6002 -131851
rect -5910 -131895 -5902 -131851
rect -5810 -131895 -5802 -131851
rect 37387 -131885 37431 -131877
rect 37487 -131885 37531 -131877
rect 37587 -131885 37631 -131877
rect 37687 -131885 37731 -131877
rect 37787 -131885 37831 -131877
rect 37887 -131885 37931 -131877
rect 37987 -131885 38031 -131877
rect 38087 -131885 38131 -131877
rect 38187 -131885 38231 -131877
rect 38287 -131885 38331 -131877
rect 38387 -131885 38431 -131877
rect 38487 -131885 38531 -131877
rect 38587 -131885 38631 -131877
rect 38687 -131885 38731 -131877
rect 38787 -131885 38831 -131877
rect 38887 -131885 38931 -131877
rect 39387 -131885 39431 -131877
rect 39487 -131885 39531 -131877
rect 39587 -131885 39631 -131877
rect 39687 -131885 39731 -131877
rect 39787 -131885 39831 -131877
rect 39887 -131885 39931 -131877
rect 39987 -131885 40031 -131877
rect 40087 -131885 40131 -131877
rect 40187 -131885 40231 -131877
rect 40287 -131885 40331 -131877
rect 40387 -131885 40431 -131877
rect 40487 -131885 40531 -131877
rect 40587 -131885 40631 -131877
rect 40687 -131885 40731 -131877
rect 40787 -131885 40831 -131877
rect 40887 -131885 40931 -131877
rect 41387 -131885 41431 -131877
rect 41487 -131885 41531 -131877
rect 41587 -131885 41631 -131877
rect 41687 -131885 41731 -131877
rect 41787 -131885 41831 -131877
rect 41887 -131885 41931 -131877
rect 41987 -131885 42031 -131877
rect 42087 -131885 42131 -131877
rect 42187 -131885 42231 -131877
rect 42287 -131885 42331 -131877
rect 42387 -131885 42431 -131877
rect 42487 -131885 42531 -131877
rect 42587 -131885 42631 -131877
rect 42687 -131885 42731 -131877
rect 42787 -131885 42831 -131877
rect 42887 -131885 42931 -131877
rect 43387 -131885 43431 -131877
rect 43487 -131885 43531 -131877
rect 43587 -131885 43631 -131877
rect 43687 -131885 43731 -131877
rect 43787 -131885 43831 -131877
rect 43887 -131885 43931 -131877
rect 43987 -131885 44031 -131877
rect 44087 -131885 44131 -131877
rect 44187 -131885 44231 -131877
rect 44287 -131885 44331 -131877
rect 44387 -131885 44431 -131877
rect 44487 -131885 44531 -131877
rect 44587 -131885 44631 -131877
rect 44687 -131885 44731 -131877
rect 44787 -131885 44831 -131877
rect 44887 -131885 44931 -131877
rect 37431 -131929 37439 -131885
rect 37531 -131929 37539 -131885
rect 37631 -131929 37639 -131885
rect 37731 -131929 37739 -131885
rect 37831 -131929 37839 -131885
rect 37931 -131929 37939 -131885
rect 38031 -131929 38039 -131885
rect 38131 -131929 38139 -131885
rect 38231 -131929 38239 -131885
rect 38331 -131929 38339 -131885
rect 38431 -131929 38439 -131885
rect 38531 -131929 38539 -131885
rect 38631 -131929 38639 -131885
rect 38731 -131929 38739 -131885
rect 38831 -131929 38839 -131885
rect 38931 -131929 38939 -131885
rect 39431 -131929 39439 -131885
rect 39531 -131929 39539 -131885
rect 39631 -131929 39639 -131885
rect 39731 -131929 39739 -131885
rect 39831 -131929 39839 -131885
rect 39931 -131929 39939 -131885
rect 40031 -131929 40039 -131885
rect 40131 -131929 40139 -131885
rect 40231 -131929 40239 -131885
rect 40331 -131929 40339 -131885
rect 40431 -131929 40439 -131885
rect 40531 -131929 40539 -131885
rect 40631 -131929 40639 -131885
rect 40731 -131929 40739 -131885
rect 40831 -131929 40839 -131885
rect 40931 -131929 40939 -131885
rect 41431 -131929 41439 -131885
rect 41531 -131929 41539 -131885
rect 41631 -131929 41639 -131885
rect 41731 -131929 41739 -131885
rect 41831 -131929 41839 -131885
rect 41931 -131929 41939 -131885
rect 42031 -131929 42039 -131885
rect 42131 -131929 42139 -131885
rect 42231 -131929 42239 -131885
rect 42331 -131929 42339 -131885
rect 42431 -131929 42439 -131885
rect 42531 -131929 42539 -131885
rect 42631 -131929 42639 -131885
rect 42731 -131929 42739 -131885
rect 42831 -131929 42839 -131885
rect 42931 -131929 42939 -131885
rect 43431 -131929 43439 -131885
rect 43531 -131929 43539 -131885
rect 43631 -131929 43639 -131885
rect 43731 -131929 43739 -131885
rect 43831 -131929 43839 -131885
rect 43931 -131929 43939 -131885
rect 44031 -131929 44039 -131885
rect 44131 -131929 44139 -131885
rect 44231 -131929 44239 -131885
rect 44331 -131929 44339 -131885
rect 44431 -131929 44439 -131885
rect 44531 -131929 44539 -131885
rect 44631 -131929 44639 -131885
rect 44731 -131929 44739 -131885
rect 44831 -131929 44839 -131885
rect 44931 -131929 44939 -131885
rect -13354 -131951 -13310 -131943
rect -13254 -131951 -13210 -131943
rect -13154 -131951 -13110 -131943
rect -13054 -131951 -13010 -131943
rect -12954 -131951 -12910 -131943
rect -12854 -131951 -12810 -131943
rect -12754 -131951 -12710 -131943
rect -12654 -131951 -12610 -131943
rect -12554 -131951 -12510 -131943
rect -12454 -131951 -12410 -131943
rect -12354 -131951 -12310 -131943
rect -12254 -131951 -12210 -131943
rect -12154 -131951 -12110 -131943
rect -12054 -131951 -12010 -131943
rect -11954 -131951 -11910 -131943
rect -11854 -131951 -11810 -131943
rect -11354 -131951 -11310 -131943
rect -11254 -131951 -11210 -131943
rect -11154 -131951 -11110 -131943
rect -11054 -131951 -11010 -131943
rect -10954 -131951 -10910 -131943
rect -10854 -131951 -10810 -131943
rect -10754 -131951 -10710 -131943
rect -10654 -131951 -10610 -131943
rect -10554 -131951 -10510 -131943
rect -10454 -131951 -10410 -131943
rect -10354 -131951 -10310 -131943
rect -10254 -131951 -10210 -131943
rect -10154 -131951 -10110 -131943
rect -10054 -131951 -10010 -131943
rect -9954 -131951 -9910 -131943
rect -9854 -131951 -9810 -131943
rect -9354 -131951 -9310 -131943
rect -9254 -131951 -9210 -131943
rect -9154 -131951 -9110 -131943
rect -9054 -131951 -9010 -131943
rect -8954 -131951 -8910 -131943
rect -8854 -131951 -8810 -131943
rect -8754 -131951 -8710 -131943
rect -8654 -131951 -8610 -131943
rect -8554 -131951 -8510 -131943
rect -8454 -131951 -8410 -131943
rect -8354 -131951 -8310 -131943
rect -8254 -131951 -8210 -131943
rect -8154 -131951 -8110 -131943
rect -8054 -131951 -8010 -131943
rect -7954 -131951 -7910 -131943
rect -7854 -131951 -7810 -131943
rect -7354 -131951 -7310 -131943
rect -7254 -131951 -7210 -131943
rect -7154 -131951 -7110 -131943
rect -7054 -131951 -7010 -131943
rect -6954 -131951 -6910 -131943
rect -6854 -131951 -6810 -131943
rect -6754 -131951 -6710 -131943
rect -6654 -131951 -6610 -131943
rect -6554 -131951 -6510 -131943
rect -6454 -131951 -6410 -131943
rect -6354 -131951 -6310 -131943
rect -6254 -131951 -6210 -131943
rect -6154 -131951 -6110 -131943
rect -6054 -131951 -6010 -131943
rect -5954 -131951 -5910 -131943
rect -5854 -131951 -5810 -131943
rect -13310 -131995 -13302 -131951
rect -13210 -131995 -13202 -131951
rect -13110 -131995 -13102 -131951
rect -13010 -131995 -13002 -131951
rect -12910 -131995 -12902 -131951
rect -12810 -131995 -12802 -131951
rect -12710 -131995 -12702 -131951
rect -12610 -131995 -12602 -131951
rect -12510 -131995 -12502 -131951
rect -12410 -131995 -12402 -131951
rect -12310 -131995 -12302 -131951
rect -12210 -131995 -12202 -131951
rect -12110 -131995 -12102 -131951
rect -12010 -131995 -12002 -131951
rect -11910 -131995 -11902 -131951
rect -11810 -131995 -11802 -131951
rect -11310 -131995 -11302 -131951
rect -11210 -131995 -11202 -131951
rect -11110 -131995 -11102 -131951
rect -11010 -131995 -11002 -131951
rect -10910 -131995 -10902 -131951
rect -10810 -131995 -10802 -131951
rect -10710 -131995 -10702 -131951
rect -10610 -131995 -10602 -131951
rect -10510 -131995 -10502 -131951
rect -10410 -131995 -10402 -131951
rect -10310 -131995 -10302 -131951
rect -10210 -131995 -10202 -131951
rect -10110 -131995 -10102 -131951
rect -10010 -131995 -10002 -131951
rect -9910 -131995 -9902 -131951
rect -9810 -131995 -9802 -131951
rect -9310 -131995 -9302 -131951
rect -9210 -131995 -9202 -131951
rect -9110 -131995 -9102 -131951
rect -9010 -131995 -9002 -131951
rect -8910 -131995 -8902 -131951
rect -8810 -131995 -8802 -131951
rect -8710 -131995 -8702 -131951
rect -8610 -131995 -8602 -131951
rect -8510 -131995 -8502 -131951
rect -8410 -131995 -8402 -131951
rect -8310 -131995 -8302 -131951
rect -8210 -131995 -8202 -131951
rect -8110 -131995 -8102 -131951
rect -8010 -131995 -8002 -131951
rect -7910 -131995 -7902 -131951
rect -7810 -131995 -7802 -131951
rect -7310 -131995 -7302 -131951
rect -7210 -131995 -7202 -131951
rect -7110 -131995 -7102 -131951
rect -7010 -131995 -7002 -131951
rect -6910 -131995 -6902 -131951
rect -6810 -131995 -6802 -131951
rect -6710 -131995 -6702 -131951
rect -6610 -131995 -6602 -131951
rect -6510 -131995 -6502 -131951
rect -6410 -131995 -6402 -131951
rect -6310 -131995 -6302 -131951
rect -6210 -131995 -6202 -131951
rect -6110 -131995 -6102 -131951
rect -6010 -131995 -6002 -131951
rect -5910 -131995 -5902 -131951
rect -5810 -131995 -5802 -131951
rect 37387 -131985 37431 -131977
rect 37487 -131985 37531 -131977
rect 37587 -131985 37631 -131977
rect 37687 -131985 37731 -131977
rect 37787 -131985 37831 -131977
rect 37887 -131985 37931 -131977
rect 37987 -131985 38031 -131977
rect 38087 -131985 38131 -131977
rect 38187 -131985 38231 -131977
rect 38287 -131985 38331 -131977
rect 38387 -131985 38431 -131977
rect 38487 -131985 38531 -131977
rect 38587 -131985 38631 -131977
rect 38687 -131985 38731 -131977
rect 38787 -131985 38831 -131977
rect 38887 -131985 38931 -131977
rect 39387 -131985 39431 -131977
rect 39487 -131985 39531 -131977
rect 39587 -131985 39631 -131977
rect 39687 -131985 39731 -131977
rect 39787 -131985 39831 -131977
rect 39887 -131985 39931 -131977
rect 39987 -131985 40031 -131977
rect 40087 -131985 40131 -131977
rect 40187 -131985 40231 -131977
rect 40287 -131985 40331 -131977
rect 40387 -131985 40431 -131977
rect 40487 -131985 40531 -131977
rect 40587 -131985 40631 -131977
rect 40687 -131985 40731 -131977
rect 40787 -131985 40831 -131977
rect 40887 -131985 40931 -131977
rect 41387 -131985 41431 -131977
rect 41487 -131985 41531 -131977
rect 41587 -131985 41631 -131977
rect 41687 -131985 41731 -131977
rect 41787 -131985 41831 -131977
rect 41887 -131985 41931 -131977
rect 41987 -131985 42031 -131977
rect 42087 -131985 42131 -131977
rect 42187 -131985 42231 -131977
rect 42287 -131985 42331 -131977
rect 42387 -131985 42431 -131977
rect 42487 -131985 42531 -131977
rect 42587 -131985 42631 -131977
rect 42687 -131985 42731 -131977
rect 42787 -131985 42831 -131977
rect 42887 -131985 42931 -131977
rect 43387 -131985 43431 -131977
rect 43487 -131985 43531 -131977
rect 43587 -131985 43631 -131977
rect 43687 -131985 43731 -131977
rect 43787 -131985 43831 -131977
rect 43887 -131985 43931 -131977
rect 43987 -131985 44031 -131977
rect 44087 -131985 44131 -131977
rect 44187 -131985 44231 -131977
rect 44287 -131985 44331 -131977
rect 44387 -131985 44431 -131977
rect 44487 -131985 44531 -131977
rect 44587 -131985 44631 -131977
rect 44687 -131985 44731 -131977
rect 44787 -131985 44831 -131977
rect 44887 -131985 44931 -131977
rect 37431 -132029 37439 -131985
rect 37531 -132029 37539 -131985
rect 37631 -132029 37639 -131985
rect 37731 -132029 37739 -131985
rect 37831 -132029 37839 -131985
rect 37931 -132029 37939 -131985
rect 38031 -132029 38039 -131985
rect 38131 -132029 38139 -131985
rect 38231 -132029 38239 -131985
rect 38331 -132029 38339 -131985
rect 38431 -132029 38439 -131985
rect 38531 -132029 38539 -131985
rect 38631 -132029 38639 -131985
rect 38731 -132029 38739 -131985
rect 38831 -132029 38839 -131985
rect 38931 -132029 38939 -131985
rect 39431 -132029 39439 -131985
rect 39531 -132029 39539 -131985
rect 39631 -132029 39639 -131985
rect 39731 -132029 39739 -131985
rect 39831 -132029 39839 -131985
rect 39931 -132029 39939 -131985
rect 40031 -132029 40039 -131985
rect 40131 -132029 40139 -131985
rect 40231 -132029 40239 -131985
rect 40331 -132029 40339 -131985
rect 40431 -132029 40439 -131985
rect 40531 -132029 40539 -131985
rect 40631 -132029 40639 -131985
rect 40731 -132029 40739 -131985
rect 40831 -132029 40839 -131985
rect 40931 -132029 40939 -131985
rect 41431 -132029 41439 -131985
rect 41531 -132029 41539 -131985
rect 41631 -132029 41639 -131985
rect 41731 -132029 41739 -131985
rect 41831 -132029 41839 -131985
rect 41931 -132029 41939 -131985
rect 42031 -132029 42039 -131985
rect 42131 -132029 42139 -131985
rect 42231 -132029 42239 -131985
rect 42331 -132029 42339 -131985
rect 42431 -132029 42439 -131985
rect 42531 -132029 42539 -131985
rect 42631 -132029 42639 -131985
rect 42731 -132029 42739 -131985
rect 42831 -132029 42839 -131985
rect 42931 -132029 42939 -131985
rect 43431 -132029 43439 -131985
rect 43531 -132029 43539 -131985
rect 43631 -132029 43639 -131985
rect 43731 -132029 43739 -131985
rect 43831 -132029 43839 -131985
rect 43931 -132029 43939 -131985
rect 44031 -132029 44039 -131985
rect 44131 -132029 44139 -131985
rect 44231 -132029 44239 -131985
rect 44331 -132029 44339 -131985
rect 44431 -132029 44439 -131985
rect 44531 -132029 44539 -131985
rect 44631 -132029 44639 -131985
rect 44731 -132029 44739 -131985
rect 44831 -132029 44839 -131985
rect 44931 -132029 44939 -131985
rect -13354 -132051 -13310 -132043
rect -13254 -132051 -13210 -132043
rect -13154 -132051 -13110 -132043
rect -13054 -132051 -13010 -132043
rect -12954 -132051 -12910 -132043
rect -12854 -132051 -12810 -132043
rect -12754 -132051 -12710 -132043
rect -12654 -132051 -12610 -132043
rect -12554 -132051 -12510 -132043
rect -12454 -132051 -12410 -132043
rect -12354 -132051 -12310 -132043
rect -12254 -132051 -12210 -132043
rect -12154 -132051 -12110 -132043
rect -12054 -132051 -12010 -132043
rect -11954 -132051 -11910 -132043
rect -11854 -132051 -11810 -132043
rect -11354 -132051 -11310 -132043
rect -11254 -132051 -11210 -132043
rect -11154 -132051 -11110 -132043
rect -11054 -132051 -11010 -132043
rect -10954 -132051 -10910 -132043
rect -10854 -132051 -10810 -132043
rect -10754 -132051 -10710 -132043
rect -10654 -132051 -10610 -132043
rect -10554 -132051 -10510 -132043
rect -10454 -132051 -10410 -132043
rect -10354 -132051 -10310 -132043
rect -10254 -132051 -10210 -132043
rect -10154 -132051 -10110 -132043
rect -10054 -132051 -10010 -132043
rect -9954 -132051 -9910 -132043
rect -9854 -132051 -9810 -132043
rect -9354 -132051 -9310 -132043
rect -9254 -132051 -9210 -132043
rect -9154 -132051 -9110 -132043
rect -9054 -132051 -9010 -132043
rect -8954 -132051 -8910 -132043
rect -8854 -132051 -8810 -132043
rect -8754 -132051 -8710 -132043
rect -8654 -132051 -8610 -132043
rect -8554 -132051 -8510 -132043
rect -8454 -132051 -8410 -132043
rect -8354 -132051 -8310 -132043
rect -8254 -132051 -8210 -132043
rect -8154 -132051 -8110 -132043
rect -8054 -132051 -8010 -132043
rect -7954 -132051 -7910 -132043
rect -7854 -132051 -7810 -132043
rect -7354 -132051 -7310 -132043
rect -7254 -132051 -7210 -132043
rect -7154 -132051 -7110 -132043
rect -7054 -132051 -7010 -132043
rect -6954 -132051 -6910 -132043
rect -6854 -132051 -6810 -132043
rect -6754 -132051 -6710 -132043
rect -6654 -132051 -6610 -132043
rect -6554 -132051 -6510 -132043
rect -6454 -132051 -6410 -132043
rect -6354 -132051 -6310 -132043
rect -6254 -132051 -6210 -132043
rect -6154 -132051 -6110 -132043
rect -6054 -132051 -6010 -132043
rect -5954 -132051 -5910 -132043
rect -5854 -132051 -5810 -132043
rect -13310 -132095 -13302 -132051
rect -13210 -132095 -13202 -132051
rect -13110 -132095 -13102 -132051
rect -13010 -132095 -13002 -132051
rect -12910 -132095 -12902 -132051
rect -12810 -132095 -12802 -132051
rect -12710 -132095 -12702 -132051
rect -12610 -132095 -12602 -132051
rect -12510 -132095 -12502 -132051
rect -12410 -132095 -12402 -132051
rect -12310 -132095 -12302 -132051
rect -12210 -132095 -12202 -132051
rect -12110 -132095 -12102 -132051
rect -12010 -132095 -12002 -132051
rect -11910 -132095 -11902 -132051
rect -11810 -132095 -11802 -132051
rect -11310 -132095 -11302 -132051
rect -11210 -132095 -11202 -132051
rect -11110 -132095 -11102 -132051
rect -11010 -132095 -11002 -132051
rect -10910 -132095 -10902 -132051
rect -10810 -132095 -10802 -132051
rect -10710 -132095 -10702 -132051
rect -10610 -132095 -10602 -132051
rect -10510 -132095 -10502 -132051
rect -10410 -132095 -10402 -132051
rect -10310 -132095 -10302 -132051
rect -10210 -132095 -10202 -132051
rect -10110 -132095 -10102 -132051
rect -10010 -132095 -10002 -132051
rect -9910 -132095 -9902 -132051
rect -9810 -132095 -9802 -132051
rect -9310 -132095 -9302 -132051
rect -9210 -132095 -9202 -132051
rect -9110 -132095 -9102 -132051
rect -9010 -132095 -9002 -132051
rect -8910 -132095 -8902 -132051
rect -8810 -132095 -8802 -132051
rect -8710 -132095 -8702 -132051
rect -8610 -132095 -8602 -132051
rect -8510 -132095 -8502 -132051
rect -8410 -132095 -8402 -132051
rect -8310 -132095 -8302 -132051
rect -8210 -132095 -8202 -132051
rect -8110 -132095 -8102 -132051
rect -8010 -132095 -8002 -132051
rect -7910 -132095 -7902 -132051
rect -7810 -132095 -7802 -132051
rect -7310 -132095 -7302 -132051
rect -7210 -132095 -7202 -132051
rect -7110 -132095 -7102 -132051
rect -7010 -132095 -7002 -132051
rect -6910 -132095 -6902 -132051
rect -6810 -132095 -6802 -132051
rect -6710 -132095 -6702 -132051
rect -6610 -132095 -6602 -132051
rect -6510 -132095 -6502 -132051
rect -6410 -132095 -6402 -132051
rect -6310 -132095 -6302 -132051
rect -6210 -132095 -6202 -132051
rect -6110 -132095 -6102 -132051
rect -6010 -132095 -6002 -132051
rect -5910 -132095 -5902 -132051
rect -5810 -132095 -5802 -132051
rect 37387 -132085 37431 -132077
rect 37487 -132085 37531 -132077
rect 37587 -132085 37631 -132077
rect 37687 -132085 37731 -132077
rect 37787 -132085 37831 -132077
rect 37887 -132085 37931 -132077
rect 37987 -132085 38031 -132077
rect 38087 -132085 38131 -132077
rect 38187 -132085 38231 -132077
rect 38287 -132085 38331 -132077
rect 38387 -132085 38431 -132077
rect 38487 -132085 38531 -132077
rect 38587 -132085 38631 -132077
rect 38687 -132085 38731 -132077
rect 38787 -132085 38831 -132077
rect 38887 -132085 38931 -132077
rect 39387 -132085 39431 -132077
rect 39487 -132085 39531 -132077
rect 39587 -132085 39631 -132077
rect 39687 -132085 39731 -132077
rect 39787 -132085 39831 -132077
rect 39887 -132085 39931 -132077
rect 39987 -132085 40031 -132077
rect 40087 -132085 40131 -132077
rect 40187 -132085 40231 -132077
rect 40287 -132085 40331 -132077
rect 40387 -132085 40431 -132077
rect 40487 -132085 40531 -132077
rect 40587 -132085 40631 -132077
rect 40687 -132085 40731 -132077
rect 40787 -132085 40831 -132077
rect 40887 -132085 40931 -132077
rect 41387 -132085 41431 -132077
rect 41487 -132085 41531 -132077
rect 41587 -132085 41631 -132077
rect 41687 -132085 41731 -132077
rect 41787 -132085 41831 -132077
rect 41887 -132085 41931 -132077
rect 41987 -132085 42031 -132077
rect 42087 -132085 42131 -132077
rect 42187 -132085 42231 -132077
rect 42287 -132085 42331 -132077
rect 42387 -132085 42431 -132077
rect 42487 -132085 42531 -132077
rect 42587 -132085 42631 -132077
rect 42687 -132085 42731 -132077
rect 42787 -132085 42831 -132077
rect 42887 -132085 42931 -132077
rect 43387 -132085 43431 -132077
rect 43487 -132085 43531 -132077
rect 43587 -132085 43631 -132077
rect 43687 -132085 43731 -132077
rect 43787 -132085 43831 -132077
rect 43887 -132085 43931 -132077
rect 43987 -132085 44031 -132077
rect 44087 -132085 44131 -132077
rect 44187 -132085 44231 -132077
rect 44287 -132085 44331 -132077
rect 44387 -132085 44431 -132077
rect 44487 -132085 44531 -132077
rect 44587 -132085 44631 -132077
rect 44687 -132085 44731 -132077
rect 44787 -132085 44831 -132077
rect 44887 -132085 44931 -132077
rect 37431 -132129 37439 -132085
rect 37531 -132129 37539 -132085
rect 37631 -132129 37639 -132085
rect 37731 -132129 37739 -132085
rect 37831 -132129 37839 -132085
rect 37931 -132129 37939 -132085
rect 38031 -132129 38039 -132085
rect 38131 -132129 38139 -132085
rect 38231 -132129 38239 -132085
rect 38331 -132129 38339 -132085
rect 38431 -132129 38439 -132085
rect 38531 -132129 38539 -132085
rect 38631 -132129 38639 -132085
rect 38731 -132129 38739 -132085
rect 38831 -132129 38839 -132085
rect 38931 -132129 38939 -132085
rect 39431 -132129 39439 -132085
rect 39531 -132129 39539 -132085
rect 39631 -132129 39639 -132085
rect 39731 -132129 39739 -132085
rect 39831 -132129 39839 -132085
rect 39931 -132129 39939 -132085
rect 40031 -132129 40039 -132085
rect 40131 -132129 40139 -132085
rect 40231 -132129 40239 -132085
rect 40331 -132129 40339 -132085
rect 40431 -132129 40439 -132085
rect 40531 -132129 40539 -132085
rect 40631 -132129 40639 -132085
rect 40731 -132129 40739 -132085
rect 40831 -132129 40839 -132085
rect 40931 -132129 40939 -132085
rect 41431 -132129 41439 -132085
rect 41531 -132129 41539 -132085
rect 41631 -132129 41639 -132085
rect 41731 -132129 41739 -132085
rect 41831 -132129 41839 -132085
rect 41931 -132129 41939 -132085
rect 42031 -132129 42039 -132085
rect 42131 -132129 42139 -132085
rect 42231 -132129 42239 -132085
rect 42331 -132129 42339 -132085
rect 42431 -132129 42439 -132085
rect 42531 -132129 42539 -132085
rect 42631 -132129 42639 -132085
rect 42731 -132129 42739 -132085
rect 42831 -132129 42839 -132085
rect 42931 -132129 42939 -132085
rect 43431 -132129 43439 -132085
rect 43531 -132129 43539 -132085
rect 43631 -132129 43639 -132085
rect 43731 -132129 43739 -132085
rect 43831 -132129 43839 -132085
rect 43931 -132129 43939 -132085
rect 44031 -132129 44039 -132085
rect 44131 -132129 44139 -132085
rect 44231 -132129 44239 -132085
rect 44331 -132129 44339 -132085
rect 44431 -132129 44439 -132085
rect 44531 -132129 44539 -132085
rect 44631 -132129 44639 -132085
rect 44731 -132129 44739 -132085
rect 44831 -132129 44839 -132085
rect 44931 -132129 44939 -132085
rect -13354 -132151 -13310 -132143
rect -13254 -132151 -13210 -132143
rect -13154 -132151 -13110 -132143
rect -13054 -132151 -13010 -132143
rect -12954 -132151 -12910 -132143
rect -12854 -132151 -12810 -132143
rect -12754 -132151 -12710 -132143
rect -12654 -132151 -12610 -132143
rect -12554 -132151 -12510 -132143
rect -12454 -132151 -12410 -132143
rect -12354 -132151 -12310 -132143
rect -12254 -132151 -12210 -132143
rect -12154 -132151 -12110 -132143
rect -12054 -132151 -12010 -132143
rect -11954 -132151 -11910 -132143
rect -11854 -132151 -11810 -132143
rect -11354 -132151 -11310 -132143
rect -11254 -132151 -11210 -132143
rect -11154 -132151 -11110 -132143
rect -11054 -132151 -11010 -132143
rect -10954 -132151 -10910 -132143
rect -10854 -132151 -10810 -132143
rect -10754 -132151 -10710 -132143
rect -10654 -132151 -10610 -132143
rect -10554 -132151 -10510 -132143
rect -10454 -132151 -10410 -132143
rect -10354 -132151 -10310 -132143
rect -10254 -132151 -10210 -132143
rect -10154 -132151 -10110 -132143
rect -10054 -132151 -10010 -132143
rect -9954 -132151 -9910 -132143
rect -9854 -132151 -9810 -132143
rect -9354 -132151 -9310 -132143
rect -9254 -132151 -9210 -132143
rect -9154 -132151 -9110 -132143
rect -9054 -132151 -9010 -132143
rect -8954 -132151 -8910 -132143
rect -8854 -132151 -8810 -132143
rect -8754 -132151 -8710 -132143
rect -8654 -132151 -8610 -132143
rect -8554 -132151 -8510 -132143
rect -8454 -132151 -8410 -132143
rect -8354 -132151 -8310 -132143
rect -8254 -132151 -8210 -132143
rect -8154 -132151 -8110 -132143
rect -8054 -132151 -8010 -132143
rect -7954 -132151 -7910 -132143
rect -7854 -132151 -7810 -132143
rect -7354 -132151 -7310 -132143
rect -7254 -132151 -7210 -132143
rect -7154 -132151 -7110 -132143
rect -7054 -132151 -7010 -132143
rect -6954 -132151 -6910 -132143
rect -6854 -132151 -6810 -132143
rect -6754 -132151 -6710 -132143
rect -6654 -132151 -6610 -132143
rect -6554 -132151 -6510 -132143
rect -6454 -132151 -6410 -132143
rect -6354 -132151 -6310 -132143
rect -6254 -132151 -6210 -132143
rect -6154 -132151 -6110 -132143
rect -6054 -132151 -6010 -132143
rect -5954 -132151 -5910 -132143
rect -5854 -132151 -5810 -132143
rect -13310 -132195 -13302 -132151
rect -13210 -132195 -13202 -132151
rect -13110 -132195 -13102 -132151
rect -13010 -132195 -13002 -132151
rect -12910 -132195 -12902 -132151
rect -12810 -132195 -12802 -132151
rect -12710 -132195 -12702 -132151
rect -12610 -132195 -12602 -132151
rect -12510 -132195 -12502 -132151
rect -12410 -132195 -12402 -132151
rect -12310 -132195 -12302 -132151
rect -12210 -132195 -12202 -132151
rect -12110 -132195 -12102 -132151
rect -12010 -132195 -12002 -132151
rect -11910 -132195 -11902 -132151
rect -11810 -132195 -11802 -132151
rect -11310 -132195 -11302 -132151
rect -11210 -132195 -11202 -132151
rect -11110 -132195 -11102 -132151
rect -11010 -132195 -11002 -132151
rect -10910 -132195 -10902 -132151
rect -10810 -132195 -10802 -132151
rect -10710 -132195 -10702 -132151
rect -10610 -132195 -10602 -132151
rect -10510 -132195 -10502 -132151
rect -10410 -132195 -10402 -132151
rect -10310 -132195 -10302 -132151
rect -10210 -132195 -10202 -132151
rect -10110 -132195 -10102 -132151
rect -10010 -132195 -10002 -132151
rect -9910 -132195 -9902 -132151
rect -9810 -132195 -9802 -132151
rect -9310 -132195 -9302 -132151
rect -9210 -132195 -9202 -132151
rect -9110 -132195 -9102 -132151
rect -9010 -132195 -9002 -132151
rect -8910 -132195 -8902 -132151
rect -8810 -132195 -8802 -132151
rect -8710 -132195 -8702 -132151
rect -8610 -132195 -8602 -132151
rect -8510 -132195 -8502 -132151
rect -8410 -132195 -8402 -132151
rect -8310 -132195 -8302 -132151
rect -8210 -132195 -8202 -132151
rect -8110 -132195 -8102 -132151
rect -8010 -132195 -8002 -132151
rect -7910 -132195 -7902 -132151
rect -7810 -132195 -7802 -132151
rect -7310 -132195 -7302 -132151
rect -7210 -132195 -7202 -132151
rect -7110 -132195 -7102 -132151
rect -7010 -132195 -7002 -132151
rect -6910 -132195 -6902 -132151
rect -6810 -132195 -6802 -132151
rect -6710 -132195 -6702 -132151
rect -6610 -132195 -6602 -132151
rect -6510 -132195 -6502 -132151
rect -6410 -132195 -6402 -132151
rect -6310 -132195 -6302 -132151
rect -6210 -132195 -6202 -132151
rect -6110 -132195 -6102 -132151
rect -6010 -132195 -6002 -132151
rect -5910 -132195 -5902 -132151
rect -5810 -132195 -5802 -132151
rect 37387 -132185 37431 -132177
rect 37487 -132185 37531 -132177
rect 37587 -132185 37631 -132177
rect 37687 -132185 37731 -132177
rect 37787 -132185 37831 -132177
rect 37887 -132185 37931 -132177
rect 37987 -132185 38031 -132177
rect 38087 -132185 38131 -132177
rect 38187 -132185 38231 -132177
rect 38287 -132185 38331 -132177
rect 38387 -132185 38431 -132177
rect 38487 -132185 38531 -132177
rect 38587 -132185 38631 -132177
rect 38687 -132185 38731 -132177
rect 38787 -132185 38831 -132177
rect 38887 -132185 38931 -132177
rect 39387 -132185 39431 -132177
rect 39487 -132185 39531 -132177
rect 39587 -132185 39631 -132177
rect 39687 -132185 39731 -132177
rect 39787 -132185 39831 -132177
rect 39887 -132185 39931 -132177
rect 39987 -132185 40031 -132177
rect 40087 -132185 40131 -132177
rect 40187 -132185 40231 -132177
rect 40287 -132185 40331 -132177
rect 40387 -132185 40431 -132177
rect 40487 -132185 40531 -132177
rect 40587 -132185 40631 -132177
rect 40687 -132185 40731 -132177
rect 40787 -132185 40831 -132177
rect 40887 -132185 40931 -132177
rect 41387 -132185 41431 -132177
rect 41487 -132185 41531 -132177
rect 41587 -132185 41631 -132177
rect 41687 -132185 41731 -132177
rect 41787 -132185 41831 -132177
rect 41887 -132185 41931 -132177
rect 41987 -132185 42031 -132177
rect 42087 -132185 42131 -132177
rect 42187 -132185 42231 -132177
rect 42287 -132185 42331 -132177
rect 42387 -132185 42431 -132177
rect 42487 -132185 42531 -132177
rect 42587 -132185 42631 -132177
rect 42687 -132185 42731 -132177
rect 42787 -132185 42831 -132177
rect 42887 -132185 42931 -132177
rect 43387 -132185 43431 -132177
rect 43487 -132185 43531 -132177
rect 43587 -132185 43631 -132177
rect 43687 -132185 43731 -132177
rect 43787 -132185 43831 -132177
rect 43887 -132185 43931 -132177
rect 43987 -132185 44031 -132177
rect 44087 -132185 44131 -132177
rect 44187 -132185 44231 -132177
rect 44287 -132185 44331 -132177
rect 44387 -132185 44431 -132177
rect 44487 -132185 44531 -132177
rect 44587 -132185 44631 -132177
rect 44687 -132185 44731 -132177
rect 44787 -132185 44831 -132177
rect 44887 -132185 44931 -132177
rect 37431 -132229 37439 -132185
rect 37531 -132229 37539 -132185
rect 37631 -132229 37639 -132185
rect 37731 -132229 37739 -132185
rect 37831 -132229 37839 -132185
rect 37931 -132229 37939 -132185
rect 38031 -132229 38039 -132185
rect 38131 -132229 38139 -132185
rect 38231 -132229 38239 -132185
rect 38331 -132229 38339 -132185
rect 38431 -132229 38439 -132185
rect 38531 -132229 38539 -132185
rect 38631 -132229 38639 -132185
rect 38731 -132229 38739 -132185
rect 38831 -132229 38839 -132185
rect 38931 -132229 38939 -132185
rect 39431 -132229 39439 -132185
rect 39531 -132229 39539 -132185
rect 39631 -132229 39639 -132185
rect 39731 -132229 39739 -132185
rect 39831 -132229 39839 -132185
rect 39931 -132229 39939 -132185
rect 40031 -132229 40039 -132185
rect 40131 -132229 40139 -132185
rect 40231 -132229 40239 -132185
rect 40331 -132229 40339 -132185
rect 40431 -132229 40439 -132185
rect 40531 -132229 40539 -132185
rect 40631 -132229 40639 -132185
rect 40731 -132229 40739 -132185
rect 40831 -132229 40839 -132185
rect 40931 -132229 40939 -132185
rect 41431 -132229 41439 -132185
rect 41531 -132229 41539 -132185
rect 41631 -132229 41639 -132185
rect 41731 -132229 41739 -132185
rect 41831 -132229 41839 -132185
rect 41931 -132229 41939 -132185
rect 42031 -132229 42039 -132185
rect 42131 -132229 42139 -132185
rect 42231 -132229 42239 -132185
rect 42331 -132229 42339 -132185
rect 42431 -132229 42439 -132185
rect 42531 -132229 42539 -132185
rect 42631 -132229 42639 -132185
rect 42731 -132229 42739 -132185
rect 42831 -132229 42839 -132185
rect 42931 -132229 42939 -132185
rect 43431 -132229 43439 -132185
rect 43531 -132229 43539 -132185
rect 43631 -132229 43639 -132185
rect 43731 -132229 43739 -132185
rect 43831 -132229 43839 -132185
rect 43931 -132229 43939 -132185
rect 44031 -132229 44039 -132185
rect 44131 -132229 44139 -132185
rect 44231 -132229 44239 -132185
rect 44331 -132229 44339 -132185
rect 44431 -132229 44439 -132185
rect 44531 -132229 44539 -132185
rect 44631 -132229 44639 -132185
rect 44731 -132229 44739 -132185
rect 44831 -132229 44839 -132185
rect 44931 -132229 44939 -132185
rect -13354 -132251 -13310 -132243
rect -13254 -132251 -13210 -132243
rect -13154 -132251 -13110 -132243
rect -13054 -132251 -13010 -132243
rect -12954 -132251 -12910 -132243
rect -12854 -132251 -12810 -132243
rect -12754 -132251 -12710 -132243
rect -12654 -132251 -12610 -132243
rect -12554 -132251 -12510 -132243
rect -12454 -132251 -12410 -132243
rect -12354 -132251 -12310 -132243
rect -12254 -132251 -12210 -132243
rect -12154 -132251 -12110 -132243
rect -12054 -132251 -12010 -132243
rect -11954 -132251 -11910 -132243
rect -11854 -132251 -11810 -132243
rect -11354 -132251 -11310 -132243
rect -11254 -132251 -11210 -132243
rect -11154 -132251 -11110 -132243
rect -11054 -132251 -11010 -132243
rect -10954 -132251 -10910 -132243
rect -10854 -132251 -10810 -132243
rect -10754 -132251 -10710 -132243
rect -10654 -132251 -10610 -132243
rect -10554 -132251 -10510 -132243
rect -10454 -132251 -10410 -132243
rect -10354 -132251 -10310 -132243
rect -10254 -132251 -10210 -132243
rect -10154 -132251 -10110 -132243
rect -10054 -132251 -10010 -132243
rect -9954 -132251 -9910 -132243
rect -9854 -132251 -9810 -132243
rect -9354 -132251 -9310 -132243
rect -9254 -132251 -9210 -132243
rect -9154 -132251 -9110 -132243
rect -9054 -132251 -9010 -132243
rect -8954 -132251 -8910 -132243
rect -8854 -132251 -8810 -132243
rect -8754 -132251 -8710 -132243
rect -8654 -132251 -8610 -132243
rect -8554 -132251 -8510 -132243
rect -8454 -132251 -8410 -132243
rect -8354 -132251 -8310 -132243
rect -8254 -132251 -8210 -132243
rect -8154 -132251 -8110 -132243
rect -8054 -132251 -8010 -132243
rect -7954 -132251 -7910 -132243
rect -7854 -132251 -7810 -132243
rect -7354 -132251 -7310 -132243
rect -7254 -132251 -7210 -132243
rect -7154 -132251 -7110 -132243
rect -7054 -132251 -7010 -132243
rect -6954 -132251 -6910 -132243
rect -6854 -132251 -6810 -132243
rect -6754 -132251 -6710 -132243
rect -6654 -132251 -6610 -132243
rect -6554 -132251 -6510 -132243
rect -6454 -132251 -6410 -132243
rect -6354 -132251 -6310 -132243
rect -6254 -132251 -6210 -132243
rect -6154 -132251 -6110 -132243
rect -6054 -132251 -6010 -132243
rect -5954 -132251 -5910 -132243
rect -5854 -132251 -5810 -132243
rect -13310 -132295 -13302 -132251
rect -13210 -132295 -13202 -132251
rect -13110 -132295 -13102 -132251
rect -13010 -132295 -13002 -132251
rect -12910 -132295 -12902 -132251
rect -12810 -132295 -12802 -132251
rect -12710 -132295 -12702 -132251
rect -12610 -132295 -12602 -132251
rect -12510 -132295 -12502 -132251
rect -12410 -132295 -12402 -132251
rect -12310 -132295 -12302 -132251
rect -12210 -132295 -12202 -132251
rect -12110 -132295 -12102 -132251
rect -12010 -132295 -12002 -132251
rect -11910 -132295 -11902 -132251
rect -11810 -132295 -11802 -132251
rect -11310 -132295 -11302 -132251
rect -11210 -132295 -11202 -132251
rect -11110 -132295 -11102 -132251
rect -11010 -132295 -11002 -132251
rect -10910 -132295 -10902 -132251
rect -10810 -132295 -10802 -132251
rect -10710 -132295 -10702 -132251
rect -10610 -132295 -10602 -132251
rect -10510 -132295 -10502 -132251
rect -10410 -132295 -10402 -132251
rect -10310 -132295 -10302 -132251
rect -10210 -132295 -10202 -132251
rect -10110 -132295 -10102 -132251
rect -10010 -132295 -10002 -132251
rect -9910 -132295 -9902 -132251
rect -9810 -132295 -9802 -132251
rect -9310 -132295 -9302 -132251
rect -9210 -132295 -9202 -132251
rect -9110 -132295 -9102 -132251
rect -9010 -132295 -9002 -132251
rect -8910 -132295 -8902 -132251
rect -8810 -132295 -8802 -132251
rect -8710 -132295 -8702 -132251
rect -8610 -132295 -8602 -132251
rect -8510 -132295 -8502 -132251
rect -8410 -132295 -8402 -132251
rect -8310 -132295 -8302 -132251
rect -8210 -132295 -8202 -132251
rect -8110 -132295 -8102 -132251
rect -8010 -132295 -8002 -132251
rect -7910 -132295 -7902 -132251
rect -7810 -132295 -7802 -132251
rect -7310 -132295 -7302 -132251
rect -7210 -132295 -7202 -132251
rect -7110 -132295 -7102 -132251
rect -7010 -132295 -7002 -132251
rect -6910 -132295 -6902 -132251
rect -6810 -132295 -6802 -132251
rect -6710 -132295 -6702 -132251
rect -6610 -132295 -6602 -132251
rect -6510 -132295 -6502 -132251
rect -6410 -132295 -6402 -132251
rect -6310 -132295 -6302 -132251
rect -6210 -132295 -6202 -132251
rect -6110 -132295 -6102 -132251
rect -6010 -132295 -6002 -132251
rect -5910 -132295 -5902 -132251
rect -5810 -132295 -5802 -132251
rect 37387 -132285 37431 -132277
rect 37487 -132285 37531 -132277
rect 37587 -132285 37631 -132277
rect 37687 -132285 37731 -132277
rect 37787 -132285 37831 -132277
rect 37887 -132285 37931 -132277
rect 37987 -132285 38031 -132277
rect 38087 -132285 38131 -132277
rect 38187 -132285 38231 -132277
rect 38287 -132285 38331 -132277
rect 38387 -132285 38431 -132277
rect 38487 -132285 38531 -132277
rect 38587 -132285 38631 -132277
rect 38687 -132285 38731 -132277
rect 38787 -132285 38831 -132277
rect 38887 -132285 38931 -132277
rect 39387 -132285 39431 -132277
rect 39487 -132285 39531 -132277
rect 39587 -132285 39631 -132277
rect 39687 -132285 39731 -132277
rect 39787 -132285 39831 -132277
rect 39887 -132285 39931 -132277
rect 39987 -132285 40031 -132277
rect 40087 -132285 40131 -132277
rect 40187 -132285 40231 -132277
rect 40287 -132285 40331 -132277
rect 40387 -132285 40431 -132277
rect 40487 -132285 40531 -132277
rect 40587 -132285 40631 -132277
rect 40687 -132285 40731 -132277
rect 40787 -132285 40831 -132277
rect 40887 -132285 40931 -132277
rect 41387 -132285 41431 -132277
rect 41487 -132285 41531 -132277
rect 41587 -132285 41631 -132277
rect 41687 -132285 41731 -132277
rect 41787 -132285 41831 -132277
rect 41887 -132285 41931 -132277
rect 41987 -132285 42031 -132277
rect 42087 -132285 42131 -132277
rect 42187 -132285 42231 -132277
rect 42287 -132285 42331 -132277
rect 42387 -132285 42431 -132277
rect 42487 -132285 42531 -132277
rect 42587 -132285 42631 -132277
rect 42687 -132285 42731 -132277
rect 42787 -132285 42831 -132277
rect 42887 -132285 42931 -132277
rect 43387 -132285 43431 -132277
rect 43487 -132285 43531 -132277
rect 43587 -132285 43631 -132277
rect 43687 -132285 43731 -132277
rect 43787 -132285 43831 -132277
rect 43887 -132285 43931 -132277
rect 43987 -132285 44031 -132277
rect 44087 -132285 44131 -132277
rect 44187 -132285 44231 -132277
rect 44287 -132285 44331 -132277
rect 44387 -132285 44431 -132277
rect 44487 -132285 44531 -132277
rect 44587 -132285 44631 -132277
rect 44687 -132285 44731 -132277
rect 44787 -132285 44831 -132277
rect 44887 -132285 44931 -132277
rect 37431 -132329 37439 -132285
rect 37531 -132329 37539 -132285
rect 37631 -132329 37639 -132285
rect 37731 -132329 37739 -132285
rect 37831 -132329 37839 -132285
rect 37931 -132329 37939 -132285
rect 38031 -132329 38039 -132285
rect 38131 -132329 38139 -132285
rect 38231 -132329 38239 -132285
rect 38331 -132329 38339 -132285
rect 38431 -132329 38439 -132285
rect 38531 -132329 38539 -132285
rect 38631 -132329 38639 -132285
rect 38731 -132329 38739 -132285
rect 38831 -132329 38839 -132285
rect 38931 -132329 38939 -132285
rect 39431 -132329 39439 -132285
rect 39531 -132329 39539 -132285
rect 39631 -132329 39639 -132285
rect 39731 -132329 39739 -132285
rect 39831 -132329 39839 -132285
rect 39931 -132329 39939 -132285
rect 40031 -132329 40039 -132285
rect 40131 -132329 40139 -132285
rect 40231 -132329 40239 -132285
rect 40331 -132329 40339 -132285
rect 40431 -132329 40439 -132285
rect 40531 -132329 40539 -132285
rect 40631 -132329 40639 -132285
rect 40731 -132329 40739 -132285
rect 40831 -132329 40839 -132285
rect 40931 -132329 40939 -132285
rect 41431 -132329 41439 -132285
rect 41531 -132329 41539 -132285
rect 41631 -132329 41639 -132285
rect 41731 -132329 41739 -132285
rect 41831 -132329 41839 -132285
rect 41931 -132329 41939 -132285
rect 42031 -132329 42039 -132285
rect 42131 -132329 42139 -132285
rect 42231 -132329 42239 -132285
rect 42331 -132329 42339 -132285
rect 42431 -132329 42439 -132285
rect 42531 -132329 42539 -132285
rect 42631 -132329 42639 -132285
rect 42731 -132329 42739 -132285
rect 42831 -132329 42839 -132285
rect 42931 -132329 42939 -132285
rect 43431 -132329 43439 -132285
rect 43531 -132329 43539 -132285
rect 43631 -132329 43639 -132285
rect 43731 -132329 43739 -132285
rect 43831 -132329 43839 -132285
rect 43931 -132329 43939 -132285
rect 44031 -132329 44039 -132285
rect 44131 -132329 44139 -132285
rect 44231 -132329 44239 -132285
rect 44331 -132329 44339 -132285
rect 44431 -132329 44439 -132285
rect 44531 -132329 44539 -132285
rect 44631 -132329 44639 -132285
rect 44731 -132329 44739 -132285
rect 44831 -132329 44839 -132285
rect 44931 -132329 44939 -132285
rect -13354 -132351 -13310 -132343
rect -13254 -132351 -13210 -132343
rect -13154 -132351 -13110 -132343
rect -13054 -132351 -13010 -132343
rect -12954 -132351 -12910 -132343
rect -12854 -132351 -12810 -132343
rect -12754 -132351 -12710 -132343
rect -12654 -132351 -12610 -132343
rect -12554 -132351 -12510 -132343
rect -12454 -132351 -12410 -132343
rect -12354 -132351 -12310 -132343
rect -12254 -132351 -12210 -132343
rect -12154 -132351 -12110 -132343
rect -12054 -132351 -12010 -132343
rect -11954 -132351 -11910 -132343
rect -11854 -132351 -11810 -132343
rect -11354 -132351 -11310 -132343
rect -11254 -132351 -11210 -132343
rect -11154 -132351 -11110 -132343
rect -11054 -132351 -11010 -132343
rect -10954 -132351 -10910 -132343
rect -10854 -132351 -10810 -132343
rect -10754 -132351 -10710 -132343
rect -10654 -132351 -10610 -132343
rect -10554 -132351 -10510 -132343
rect -10454 -132351 -10410 -132343
rect -10354 -132351 -10310 -132343
rect -10254 -132351 -10210 -132343
rect -10154 -132351 -10110 -132343
rect -10054 -132351 -10010 -132343
rect -9954 -132351 -9910 -132343
rect -9854 -132351 -9810 -132343
rect -9354 -132351 -9310 -132343
rect -9254 -132351 -9210 -132343
rect -9154 -132351 -9110 -132343
rect -9054 -132351 -9010 -132343
rect -8954 -132351 -8910 -132343
rect -8854 -132351 -8810 -132343
rect -8754 -132351 -8710 -132343
rect -8654 -132351 -8610 -132343
rect -8554 -132351 -8510 -132343
rect -8454 -132351 -8410 -132343
rect -8354 -132351 -8310 -132343
rect -8254 -132351 -8210 -132343
rect -8154 -132351 -8110 -132343
rect -8054 -132351 -8010 -132343
rect -7954 -132351 -7910 -132343
rect -7854 -132351 -7810 -132343
rect -7354 -132351 -7310 -132343
rect -7254 -132351 -7210 -132343
rect -7154 -132351 -7110 -132343
rect -7054 -132351 -7010 -132343
rect -6954 -132351 -6910 -132343
rect -6854 -132351 -6810 -132343
rect -6754 -132351 -6710 -132343
rect -6654 -132351 -6610 -132343
rect -6554 -132351 -6510 -132343
rect -6454 -132351 -6410 -132343
rect -6354 -132351 -6310 -132343
rect -6254 -132351 -6210 -132343
rect -6154 -132351 -6110 -132343
rect -6054 -132351 -6010 -132343
rect -5954 -132351 -5910 -132343
rect -5854 -132351 -5810 -132343
rect -13310 -132395 -13302 -132351
rect -13210 -132395 -13202 -132351
rect -13110 -132395 -13102 -132351
rect -13010 -132395 -13002 -132351
rect -12910 -132395 -12902 -132351
rect -12810 -132395 -12802 -132351
rect -12710 -132395 -12702 -132351
rect -12610 -132395 -12602 -132351
rect -12510 -132395 -12502 -132351
rect -12410 -132395 -12402 -132351
rect -12310 -132395 -12302 -132351
rect -12210 -132395 -12202 -132351
rect -12110 -132395 -12102 -132351
rect -12010 -132395 -12002 -132351
rect -11910 -132395 -11902 -132351
rect -11810 -132395 -11802 -132351
rect -11310 -132395 -11302 -132351
rect -11210 -132395 -11202 -132351
rect -11110 -132395 -11102 -132351
rect -11010 -132395 -11002 -132351
rect -10910 -132395 -10902 -132351
rect -10810 -132395 -10802 -132351
rect -10710 -132395 -10702 -132351
rect -10610 -132395 -10602 -132351
rect -10510 -132395 -10502 -132351
rect -10410 -132395 -10402 -132351
rect -10310 -132395 -10302 -132351
rect -10210 -132395 -10202 -132351
rect -10110 -132395 -10102 -132351
rect -10010 -132395 -10002 -132351
rect -9910 -132395 -9902 -132351
rect -9810 -132395 -9802 -132351
rect -9310 -132395 -9302 -132351
rect -9210 -132395 -9202 -132351
rect -9110 -132395 -9102 -132351
rect -9010 -132395 -9002 -132351
rect -8910 -132395 -8902 -132351
rect -8810 -132395 -8802 -132351
rect -8710 -132395 -8702 -132351
rect -8610 -132395 -8602 -132351
rect -8510 -132395 -8502 -132351
rect -8410 -132395 -8402 -132351
rect -8310 -132395 -8302 -132351
rect -8210 -132395 -8202 -132351
rect -8110 -132395 -8102 -132351
rect -8010 -132395 -8002 -132351
rect -7910 -132395 -7902 -132351
rect -7810 -132395 -7802 -132351
rect -7310 -132395 -7302 -132351
rect -7210 -132395 -7202 -132351
rect -7110 -132395 -7102 -132351
rect -7010 -132395 -7002 -132351
rect -6910 -132395 -6902 -132351
rect -6810 -132395 -6802 -132351
rect -6710 -132395 -6702 -132351
rect -6610 -132395 -6602 -132351
rect -6510 -132395 -6502 -132351
rect -6410 -132395 -6402 -132351
rect -6310 -132395 -6302 -132351
rect -6210 -132395 -6202 -132351
rect -6110 -132395 -6102 -132351
rect -6010 -132395 -6002 -132351
rect -5910 -132395 -5902 -132351
rect -5810 -132395 -5802 -132351
rect 37387 -132385 37431 -132377
rect 37487 -132385 37531 -132377
rect 37587 -132385 37631 -132377
rect 37687 -132385 37731 -132377
rect 37787 -132385 37831 -132377
rect 37887 -132385 37931 -132377
rect 37987 -132385 38031 -132377
rect 38087 -132385 38131 -132377
rect 38187 -132385 38231 -132377
rect 38287 -132385 38331 -132377
rect 38387 -132385 38431 -132377
rect 38487 -132385 38531 -132377
rect 38587 -132385 38631 -132377
rect 38687 -132385 38731 -132377
rect 38787 -132385 38831 -132377
rect 38887 -132385 38931 -132377
rect 39387 -132385 39431 -132377
rect 39487 -132385 39531 -132377
rect 39587 -132385 39631 -132377
rect 39687 -132385 39731 -132377
rect 39787 -132385 39831 -132377
rect 39887 -132385 39931 -132377
rect 39987 -132385 40031 -132377
rect 40087 -132385 40131 -132377
rect 40187 -132385 40231 -132377
rect 40287 -132385 40331 -132377
rect 40387 -132385 40431 -132377
rect 40487 -132385 40531 -132377
rect 40587 -132385 40631 -132377
rect 40687 -132385 40731 -132377
rect 40787 -132385 40831 -132377
rect 40887 -132385 40931 -132377
rect 41387 -132385 41431 -132377
rect 41487 -132385 41531 -132377
rect 41587 -132385 41631 -132377
rect 41687 -132385 41731 -132377
rect 41787 -132385 41831 -132377
rect 41887 -132385 41931 -132377
rect 41987 -132385 42031 -132377
rect 42087 -132385 42131 -132377
rect 42187 -132385 42231 -132377
rect 42287 -132385 42331 -132377
rect 42387 -132385 42431 -132377
rect 42487 -132385 42531 -132377
rect 42587 -132385 42631 -132377
rect 42687 -132385 42731 -132377
rect 42787 -132385 42831 -132377
rect 42887 -132385 42931 -132377
rect 43387 -132385 43431 -132377
rect 43487 -132385 43531 -132377
rect 43587 -132385 43631 -132377
rect 43687 -132385 43731 -132377
rect 43787 -132385 43831 -132377
rect 43887 -132385 43931 -132377
rect 43987 -132385 44031 -132377
rect 44087 -132385 44131 -132377
rect 44187 -132385 44231 -132377
rect 44287 -132385 44331 -132377
rect 44387 -132385 44431 -132377
rect 44487 -132385 44531 -132377
rect 44587 -132385 44631 -132377
rect 44687 -132385 44731 -132377
rect 44787 -132385 44831 -132377
rect 44887 -132385 44931 -132377
rect 37431 -132429 37439 -132385
rect 37531 -132429 37539 -132385
rect 37631 -132429 37639 -132385
rect 37731 -132429 37739 -132385
rect 37831 -132429 37839 -132385
rect 37931 -132429 37939 -132385
rect 38031 -132429 38039 -132385
rect 38131 -132429 38139 -132385
rect 38231 -132429 38239 -132385
rect 38331 -132429 38339 -132385
rect 38431 -132429 38439 -132385
rect 38531 -132429 38539 -132385
rect 38631 -132429 38639 -132385
rect 38731 -132429 38739 -132385
rect 38831 -132429 38839 -132385
rect 38931 -132429 38939 -132385
rect 39431 -132429 39439 -132385
rect 39531 -132429 39539 -132385
rect 39631 -132429 39639 -132385
rect 39731 -132429 39739 -132385
rect 39831 -132429 39839 -132385
rect 39931 -132429 39939 -132385
rect 40031 -132429 40039 -132385
rect 40131 -132429 40139 -132385
rect 40231 -132429 40239 -132385
rect 40331 -132429 40339 -132385
rect 40431 -132429 40439 -132385
rect 40531 -132429 40539 -132385
rect 40631 -132429 40639 -132385
rect 40731 -132429 40739 -132385
rect 40831 -132429 40839 -132385
rect 40931 -132429 40939 -132385
rect 41431 -132429 41439 -132385
rect 41531 -132429 41539 -132385
rect 41631 -132429 41639 -132385
rect 41731 -132429 41739 -132385
rect 41831 -132429 41839 -132385
rect 41931 -132429 41939 -132385
rect 42031 -132429 42039 -132385
rect 42131 -132429 42139 -132385
rect 42231 -132429 42239 -132385
rect 42331 -132429 42339 -132385
rect 42431 -132429 42439 -132385
rect 42531 -132429 42539 -132385
rect 42631 -132429 42639 -132385
rect 42731 -132429 42739 -132385
rect 42831 -132429 42839 -132385
rect 42931 -132429 42939 -132385
rect 43431 -132429 43439 -132385
rect 43531 -132429 43539 -132385
rect 43631 -132429 43639 -132385
rect 43731 -132429 43739 -132385
rect 43831 -132429 43839 -132385
rect 43931 -132429 43939 -132385
rect 44031 -132429 44039 -132385
rect 44131 -132429 44139 -132385
rect 44231 -132429 44239 -132385
rect 44331 -132429 44339 -132385
rect 44431 -132429 44439 -132385
rect 44531 -132429 44539 -132385
rect 44631 -132429 44639 -132385
rect 44731 -132429 44739 -132385
rect 44831 -132429 44839 -132385
rect 44931 -132429 44939 -132385
rect -13354 -132451 -13310 -132443
rect -13254 -132451 -13210 -132443
rect -13154 -132451 -13110 -132443
rect -13054 -132451 -13010 -132443
rect -12954 -132451 -12910 -132443
rect -12854 -132451 -12810 -132443
rect -12754 -132451 -12710 -132443
rect -12654 -132451 -12610 -132443
rect -12554 -132451 -12510 -132443
rect -12454 -132451 -12410 -132443
rect -12354 -132451 -12310 -132443
rect -12254 -132451 -12210 -132443
rect -12154 -132451 -12110 -132443
rect -12054 -132451 -12010 -132443
rect -11954 -132451 -11910 -132443
rect -11854 -132451 -11810 -132443
rect -11354 -132451 -11310 -132443
rect -11254 -132451 -11210 -132443
rect -11154 -132451 -11110 -132443
rect -11054 -132451 -11010 -132443
rect -10954 -132451 -10910 -132443
rect -10854 -132451 -10810 -132443
rect -10754 -132451 -10710 -132443
rect -10654 -132451 -10610 -132443
rect -10554 -132451 -10510 -132443
rect -10454 -132451 -10410 -132443
rect -10354 -132451 -10310 -132443
rect -10254 -132451 -10210 -132443
rect -10154 -132451 -10110 -132443
rect -10054 -132451 -10010 -132443
rect -9954 -132451 -9910 -132443
rect -9854 -132451 -9810 -132443
rect -9354 -132451 -9310 -132443
rect -9254 -132451 -9210 -132443
rect -9154 -132451 -9110 -132443
rect -9054 -132451 -9010 -132443
rect -8954 -132451 -8910 -132443
rect -8854 -132451 -8810 -132443
rect -8754 -132451 -8710 -132443
rect -8654 -132451 -8610 -132443
rect -8554 -132451 -8510 -132443
rect -8454 -132451 -8410 -132443
rect -8354 -132451 -8310 -132443
rect -8254 -132451 -8210 -132443
rect -8154 -132451 -8110 -132443
rect -8054 -132451 -8010 -132443
rect -7954 -132451 -7910 -132443
rect -7854 -132451 -7810 -132443
rect -7354 -132451 -7310 -132443
rect -7254 -132451 -7210 -132443
rect -7154 -132451 -7110 -132443
rect -7054 -132451 -7010 -132443
rect -6954 -132451 -6910 -132443
rect -6854 -132451 -6810 -132443
rect -6754 -132451 -6710 -132443
rect -6654 -132451 -6610 -132443
rect -6554 -132451 -6510 -132443
rect -6454 -132451 -6410 -132443
rect -6354 -132451 -6310 -132443
rect -6254 -132451 -6210 -132443
rect -6154 -132451 -6110 -132443
rect -6054 -132451 -6010 -132443
rect -5954 -132451 -5910 -132443
rect -5854 -132451 -5810 -132443
rect -13310 -132495 -13302 -132451
rect -13210 -132495 -13202 -132451
rect -13110 -132495 -13102 -132451
rect -13010 -132495 -13002 -132451
rect -12910 -132495 -12902 -132451
rect -12810 -132495 -12802 -132451
rect -12710 -132495 -12702 -132451
rect -12610 -132495 -12602 -132451
rect -12510 -132495 -12502 -132451
rect -12410 -132495 -12402 -132451
rect -12310 -132495 -12302 -132451
rect -12210 -132495 -12202 -132451
rect -12110 -132495 -12102 -132451
rect -12010 -132495 -12002 -132451
rect -11910 -132495 -11902 -132451
rect -11810 -132495 -11802 -132451
rect -11310 -132495 -11302 -132451
rect -11210 -132495 -11202 -132451
rect -11110 -132495 -11102 -132451
rect -11010 -132495 -11002 -132451
rect -10910 -132495 -10902 -132451
rect -10810 -132495 -10802 -132451
rect -10710 -132495 -10702 -132451
rect -10610 -132495 -10602 -132451
rect -10510 -132495 -10502 -132451
rect -10410 -132495 -10402 -132451
rect -10310 -132495 -10302 -132451
rect -10210 -132495 -10202 -132451
rect -10110 -132495 -10102 -132451
rect -10010 -132495 -10002 -132451
rect -9910 -132495 -9902 -132451
rect -9810 -132495 -9802 -132451
rect -9310 -132495 -9302 -132451
rect -9210 -132495 -9202 -132451
rect -9110 -132495 -9102 -132451
rect -9010 -132495 -9002 -132451
rect -8910 -132495 -8902 -132451
rect -8810 -132495 -8802 -132451
rect -8710 -132495 -8702 -132451
rect -8610 -132495 -8602 -132451
rect -8510 -132495 -8502 -132451
rect -8410 -132495 -8402 -132451
rect -8310 -132495 -8302 -132451
rect -8210 -132495 -8202 -132451
rect -8110 -132495 -8102 -132451
rect -8010 -132495 -8002 -132451
rect -7910 -132495 -7902 -132451
rect -7810 -132495 -7802 -132451
rect -7310 -132495 -7302 -132451
rect -7210 -132495 -7202 -132451
rect -7110 -132495 -7102 -132451
rect -7010 -132495 -7002 -132451
rect -6910 -132495 -6902 -132451
rect -6810 -132495 -6802 -132451
rect -6710 -132495 -6702 -132451
rect -6610 -132495 -6602 -132451
rect -6510 -132495 -6502 -132451
rect -6410 -132495 -6402 -132451
rect -6310 -132495 -6302 -132451
rect -6210 -132495 -6202 -132451
rect -6110 -132495 -6102 -132451
rect -6010 -132495 -6002 -132451
rect -5910 -132495 -5902 -132451
rect -5810 -132495 -5802 -132451
rect 37387 -132485 37431 -132477
rect 37487 -132485 37531 -132477
rect 37587 -132485 37631 -132477
rect 37687 -132485 37731 -132477
rect 37787 -132485 37831 -132477
rect 37887 -132485 37931 -132477
rect 37987 -132485 38031 -132477
rect 38087 -132485 38131 -132477
rect 38187 -132485 38231 -132477
rect 38287 -132485 38331 -132477
rect 38387 -132485 38431 -132477
rect 38487 -132485 38531 -132477
rect 38587 -132485 38631 -132477
rect 38687 -132485 38731 -132477
rect 38787 -132485 38831 -132477
rect 38887 -132485 38931 -132477
rect 39387 -132485 39431 -132477
rect 39487 -132485 39531 -132477
rect 39587 -132485 39631 -132477
rect 39687 -132485 39731 -132477
rect 39787 -132485 39831 -132477
rect 39887 -132485 39931 -132477
rect 39987 -132485 40031 -132477
rect 40087 -132485 40131 -132477
rect 40187 -132485 40231 -132477
rect 40287 -132485 40331 -132477
rect 40387 -132485 40431 -132477
rect 40487 -132485 40531 -132477
rect 40587 -132485 40631 -132477
rect 40687 -132485 40731 -132477
rect 40787 -132485 40831 -132477
rect 40887 -132485 40931 -132477
rect 41387 -132485 41431 -132477
rect 41487 -132485 41531 -132477
rect 41587 -132485 41631 -132477
rect 41687 -132485 41731 -132477
rect 41787 -132485 41831 -132477
rect 41887 -132485 41931 -132477
rect 41987 -132485 42031 -132477
rect 42087 -132485 42131 -132477
rect 42187 -132485 42231 -132477
rect 42287 -132485 42331 -132477
rect 42387 -132485 42431 -132477
rect 42487 -132485 42531 -132477
rect 42587 -132485 42631 -132477
rect 42687 -132485 42731 -132477
rect 42787 -132485 42831 -132477
rect 42887 -132485 42931 -132477
rect 43387 -132485 43431 -132477
rect 43487 -132485 43531 -132477
rect 43587 -132485 43631 -132477
rect 43687 -132485 43731 -132477
rect 43787 -132485 43831 -132477
rect 43887 -132485 43931 -132477
rect 43987 -132485 44031 -132477
rect 44087 -132485 44131 -132477
rect 44187 -132485 44231 -132477
rect 44287 -132485 44331 -132477
rect 44387 -132485 44431 -132477
rect 44487 -132485 44531 -132477
rect 44587 -132485 44631 -132477
rect 44687 -132485 44731 -132477
rect 44787 -132485 44831 -132477
rect 44887 -132485 44931 -132477
rect 37431 -132529 37439 -132485
rect 37531 -132529 37539 -132485
rect 37631 -132529 37639 -132485
rect 37731 -132529 37739 -132485
rect 37831 -132529 37839 -132485
rect 37931 -132529 37939 -132485
rect 38031 -132529 38039 -132485
rect 38131 -132529 38139 -132485
rect 38231 -132529 38239 -132485
rect 38331 -132529 38339 -132485
rect 38431 -132529 38439 -132485
rect 38531 -132529 38539 -132485
rect 38631 -132529 38639 -132485
rect 38731 -132529 38739 -132485
rect 38831 -132529 38839 -132485
rect 38931 -132529 38939 -132485
rect 39431 -132529 39439 -132485
rect 39531 -132529 39539 -132485
rect 39631 -132529 39639 -132485
rect 39731 -132529 39739 -132485
rect 39831 -132529 39839 -132485
rect 39931 -132529 39939 -132485
rect 40031 -132529 40039 -132485
rect 40131 -132529 40139 -132485
rect 40231 -132529 40239 -132485
rect 40331 -132529 40339 -132485
rect 40431 -132529 40439 -132485
rect 40531 -132529 40539 -132485
rect 40631 -132529 40639 -132485
rect 40731 -132529 40739 -132485
rect 40831 -132529 40839 -132485
rect 40931 -132529 40939 -132485
rect 41431 -132529 41439 -132485
rect 41531 -132529 41539 -132485
rect 41631 -132529 41639 -132485
rect 41731 -132529 41739 -132485
rect 41831 -132529 41839 -132485
rect 41931 -132529 41939 -132485
rect 42031 -132529 42039 -132485
rect 42131 -132529 42139 -132485
rect 42231 -132529 42239 -132485
rect 42331 -132529 42339 -132485
rect 42431 -132529 42439 -132485
rect 42531 -132529 42539 -132485
rect 42631 -132529 42639 -132485
rect 42731 -132529 42739 -132485
rect 42831 -132529 42839 -132485
rect 42931 -132529 42939 -132485
rect 43431 -132529 43439 -132485
rect 43531 -132529 43539 -132485
rect 43631 -132529 43639 -132485
rect 43731 -132529 43739 -132485
rect 43831 -132529 43839 -132485
rect 43931 -132529 43939 -132485
rect 44031 -132529 44039 -132485
rect 44131 -132529 44139 -132485
rect 44231 -132529 44239 -132485
rect 44331 -132529 44339 -132485
rect 44431 -132529 44439 -132485
rect 44531 -132529 44539 -132485
rect 44631 -132529 44639 -132485
rect 44731 -132529 44739 -132485
rect 44831 -132529 44839 -132485
rect 44931 -132529 44939 -132485
rect -13354 -132551 -13310 -132543
rect -13254 -132551 -13210 -132543
rect -13154 -132551 -13110 -132543
rect -13054 -132551 -13010 -132543
rect -12954 -132551 -12910 -132543
rect -12854 -132551 -12810 -132543
rect -12754 -132551 -12710 -132543
rect -12654 -132551 -12610 -132543
rect -12554 -132551 -12510 -132543
rect -12454 -132551 -12410 -132543
rect -12354 -132551 -12310 -132543
rect -12254 -132551 -12210 -132543
rect -12154 -132551 -12110 -132543
rect -12054 -132551 -12010 -132543
rect -11954 -132551 -11910 -132543
rect -11854 -132551 -11810 -132543
rect -11354 -132551 -11310 -132543
rect -11254 -132551 -11210 -132543
rect -11154 -132551 -11110 -132543
rect -11054 -132551 -11010 -132543
rect -10954 -132551 -10910 -132543
rect -10854 -132551 -10810 -132543
rect -10754 -132551 -10710 -132543
rect -10654 -132551 -10610 -132543
rect -10554 -132551 -10510 -132543
rect -10454 -132551 -10410 -132543
rect -10354 -132551 -10310 -132543
rect -10254 -132551 -10210 -132543
rect -10154 -132551 -10110 -132543
rect -10054 -132551 -10010 -132543
rect -9954 -132551 -9910 -132543
rect -9854 -132551 -9810 -132543
rect -9354 -132551 -9310 -132543
rect -9254 -132551 -9210 -132543
rect -9154 -132551 -9110 -132543
rect -9054 -132551 -9010 -132543
rect -8954 -132551 -8910 -132543
rect -8854 -132551 -8810 -132543
rect -8754 -132551 -8710 -132543
rect -8654 -132551 -8610 -132543
rect -8554 -132551 -8510 -132543
rect -8454 -132551 -8410 -132543
rect -8354 -132551 -8310 -132543
rect -8254 -132551 -8210 -132543
rect -8154 -132551 -8110 -132543
rect -8054 -132551 -8010 -132543
rect -7954 -132551 -7910 -132543
rect -7854 -132551 -7810 -132543
rect -7354 -132551 -7310 -132543
rect -7254 -132551 -7210 -132543
rect -7154 -132551 -7110 -132543
rect -7054 -132551 -7010 -132543
rect -6954 -132551 -6910 -132543
rect -6854 -132551 -6810 -132543
rect -6754 -132551 -6710 -132543
rect -6654 -132551 -6610 -132543
rect -6554 -132551 -6510 -132543
rect -6454 -132551 -6410 -132543
rect -6354 -132551 -6310 -132543
rect -6254 -132551 -6210 -132543
rect -6154 -132551 -6110 -132543
rect -6054 -132551 -6010 -132543
rect -5954 -132551 -5910 -132543
rect -5854 -132551 -5810 -132543
rect -13310 -132595 -13302 -132551
rect -13210 -132595 -13202 -132551
rect -13110 -132595 -13102 -132551
rect -13010 -132595 -13002 -132551
rect -12910 -132595 -12902 -132551
rect -12810 -132595 -12802 -132551
rect -12710 -132595 -12702 -132551
rect -12610 -132595 -12602 -132551
rect -12510 -132595 -12502 -132551
rect -12410 -132595 -12402 -132551
rect -12310 -132595 -12302 -132551
rect -12210 -132595 -12202 -132551
rect -12110 -132595 -12102 -132551
rect -12010 -132595 -12002 -132551
rect -11910 -132595 -11902 -132551
rect -11810 -132595 -11802 -132551
rect -11310 -132595 -11302 -132551
rect -11210 -132595 -11202 -132551
rect -11110 -132595 -11102 -132551
rect -11010 -132595 -11002 -132551
rect -10910 -132595 -10902 -132551
rect -10810 -132595 -10802 -132551
rect -10710 -132595 -10702 -132551
rect -10610 -132595 -10602 -132551
rect -10510 -132595 -10502 -132551
rect -10410 -132595 -10402 -132551
rect -10310 -132595 -10302 -132551
rect -10210 -132595 -10202 -132551
rect -10110 -132595 -10102 -132551
rect -10010 -132595 -10002 -132551
rect -9910 -132595 -9902 -132551
rect -9810 -132595 -9802 -132551
rect -9310 -132595 -9302 -132551
rect -9210 -132595 -9202 -132551
rect -9110 -132595 -9102 -132551
rect -9010 -132595 -9002 -132551
rect -8910 -132595 -8902 -132551
rect -8810 -132595 -8802 -132551
rect -8710 -132595 -8702 -132551
rect -8610 -132595 -8602 -132551
rect -8510 -132595 -8502 -132551
rect -8410 -132595 -8402 -132551
rect -8310 -132595 -8302 -132551
rect -8210 -132595 -8202 -132551
rect -8110 -132595 -8102 -132551
rect -8010 -132595 -8002 -132551
rect -7910 -132595 -7902 -132551
rect -7810 -132595 -7802 -132551
rect -7310 -132595 -7302 -132551
rect -7210 -132595 -7202 -132551
rect -7110 -132595 -7102 -132551
rect -7010 -132595 -7002 -132551
rect -6910 -132595 -6902 -132551
rect -6810 -132595 -6802 -132551
rect -6710 -132595 -6702 -132551
rect -6610 -132595 -6602 -132551
rect -6510 -132595 -6502 -132551
rect -6410 -132595 -6402 -132551
rect -6310 -132595 -6302 -132551
rect -6210 -132595 -6202 -132551
rect -6110 -132595 -6102 -132551
rect -6010 -132595 -6002 -132551
rect -5910 -132595 -5902 -132551
rect -5810 -132595 -5802 -132551
rect 37387 -132585 37431 -132577
rect 37487 -132585 37531 -132577
rect 37587 -132585 37631 -132577
rect 37687 -132585 37731 -132577
rect 37787 -132585 37831 -132577
rect 37887 -132585 37931 -132577
rect 37987 -132585 38031 -132577
rect 38087 -132585 38131 -132577
rect 38187 -132585 38231 -132577
rect 38287 -132585 38331 -132577
rect 38387 -132585 38431 -132577
rect 38487 -132585 38531 -132577
rect 38587 -132585 38631 -132577
rect 38687 -132585 38731 -132577
rect 38787 -132585 38831 -132577
rect 38887 -132585 38931 -132577
rect 39387 -132585 39431 -132577
rect 39487 -132585 39531 -132577
rect 39587 -132585 39631 -132577
rect 39687 -132585 39731 -132577
rect 39787 -132585 39831 -132577
rect 39887 -132585 39931 -132577
rect 39987 -132585 40031 -132577
rect 40087 -132585 40131 -132577
rect 40187 -132585 40231 -132577
rect 40287 -132585 40331 -132577
rect 40387 -132585 40431 -132577
rect 40487 -132585 40531 -132577
rect 40587 -132585 40631 -132577
rect 40687 -132585 40731 -132577
rect 40787 -132585 40831 -132577
rect 40887 -132585 40931 -132577
rect 41387 -132585 41431 -132577
rect 41487 -132585 41531 -132577
rect 41587 -132585 41631 -132577
rect 41687 -132585 41731 -132577
rect 41787 -132585 41831 -132577
rect 41887 -132585 41931 -132577
rect 41987 -132585 42031 -132577
rect 42087 -132585 42131 -132577
rect 42187 -132585 42231 -132577
rect 42287 -132585 42331 -132577
rect 42387 -132585 42431 -132577
rect 42487 -132585 42531 -132577
rect 42587 -132585 42631 -132577
rect 42687 -132585 42731 -132577
rect 42787 -132585 42831 -132577
rect 42887 -132585 42931 -132577
rect 43387 -132585 43431 -132577
rect 43487 -132585 43531 -132577
rect 43587 -132585 43631 -132577
rect 43687 -132585 43731 -132577
rect 43787 -132585 43831 -132577
rect 43887 -132585 43931 -132577
rect 43987 -132585 44031 -132577
rect 44087 -132585 44131 -132577
rect 44187 -132585 44231 -132577
rect 44287 -132585 44331 -132577
rect 44387 -132585 44431 -132577
rect 44487 -132585 44531 -132577
rect 44587 -132585 44631 -132577
rect 44687 -132585 44731 -132577
rect 44787 -132585 44831 -132577
rect 44887 -132585 44931 -132577
rect 37431 -132629 37439 -132585
rect 37531 -132629 37539 -132585
rect 37631 -132629 37639 -132585
rect 37731 -132629 37739 -132585
rect 37831 -132629 37839 -132585
rect 37931 -132629 37939 -132585
rect 38031 -132629 38039 -132585
rect 38131 -132629 38139 -132585
rect 38231 -132629 38239 -132585
rect 38331 -132629 38339 -132585
rect 38431 -132629 38439 -132585
rect 38531 -132629 38539 -132585
rect 38631 -132629 38639 -132585
rect 38731 -132629 38739 -132585
rect 38831 -132629 38839 -132585
rect 38931 -132629 38939 -132585
rect 39431 -132629 39439 -132585
rect 39531 -132629 39539 -132585
rect 39631 -132629 39639 -132585
rect 39731 -132629 39739 -132585
rect 39831 -132629 39839 -132585
rect 39931 -132629 39939 -132585
rect 40031 -132629 40039 -132585
rect 40131 -132629 40139 -132585
rect 40231 -132629 40239 -132585
rect 40331 -132629 40339 -132585
rect 40431 -132629 40439 -132585
rect 40531 -132629 40539 -132585
rect 40631 -132629 40639 -132585
rect 40731 -132629 40739 -132585
rect 40831 -132629 40839 -132585
rect 40931 -132629 40939 -132585
rect 41431 -132629 41439 -132585
rect 41531 -132629 41539 -132585
rect 41631 -132629 41639 -132585
rect 41731 -132629 41739 -132585
rect 41831 -132629 41839 -132585
rect 41931 -132629 41939 -132585
rect 42031 -132629 42039 -132585
rect 42131 -132629 42139 -132585
rect 42231 -132629 42239 -132585
rect 42331 -132629 42339 -132585
rect 42431 -132629 42439 -132585
rect 42531 -132629 42539 -132585
rect 42631 -132629 42639 -132585
rect 42731 -132629 42739 -132585
rect 42831 -132629 42839 -132585
rect 42931 -132629 42939 -132585
rect 43431 -132629 43439 -132585
rect 43531 -132629 43539 -132585
rect 43631 -132629 43639 -132585
rect 43731 -132629 43739 -132585
rect 43831 -132629 43839 -132585
rect 43931 -132629 43939 -132585
rect 44031 -132629 44039 -132585
rect 44131 -132629 44139 -132585
rect 44231 -132629 44239 -132585
rect 44331 -132629 44339 -132585
rect 44431 -132629 44439 -132585
rect 44531 -132629 44539 -132585
rect 44631 -132629 44639 -132585
rect 44731 -132629 44739 -132585
rect 44831 -132629 44839 -132585
rect 44931 -132629 44939 -132585
rect -13354 -132651 -13310 -132643
rect -13254 -132651 -13210 -132643
rect -13154 -132651 -13110 -132643
rect -13054 -132651 -13010 -132643
rect -12954 -132651 -12910 -132643
rect -12854 -132651 -12810 -132643
rect -12754 -132651 -12710 -132643
rect -12654 -132651 -12610 -132643
rect -12554 -132651 -12510 -132643
rect -12454 -132651 -12410 -132643
rect -12354 -132651 -12310 -132643
rect -12254 -132651 -12210 -132643
rect -12154 -132651 -12110 -132643
rect -12054 -132651 -12010 -132643
rect -11954 -132651 -11910 -132643
rect -11854 -132651 -11810 -132643
rect -11354 -132651 -11310 -132643
rect -11254 -132651 -11210 -132643
rect -11154 -132651 -11110 -132643
rect -11054 -132651 -11010 -132643
rect -10954 -132651 -10910 -132643
rect -10854 -132651 -10810 -132643
rect -10754 -132651 -10710 -132643
rect -10654 -132651 -10610 -132643
rect -10554 -132651 -10510 -132643
rect -10454 -132651 -10410 -132643
rect -10354 -132651 -10310 -132643
rect -10254 -132651 -10210 -132643
rect -10154 -132651 -10110 -132643
rect -10054 -132651 -10010 -132643
rect -9954 -132651 -9910 -132643
rect -9854 -132651 -9810 -132643
rect -9354 -132651 -9310 -132643
rect -9254 -132651 -9210 -132643
rect -9154 -132651 -9110 -132643
rect -9054 -132651 -9010 -132643
rect -8954 -132651 -8910 -132643
rect -8854 -132651 -8810 -132643
rect -8754 -132651 -8710 -132643
rect -8654 -132651 -8610 -132643
rect -8554 -132651 -8510 -132643
rect -8454 -132651 -8410 -132643
rect -8354 -132651 -8310 -132643
rect -8254 -132651 -8210 -132643
rect -8154 -132651 -8110 -132643
rect -8054 -132651 -8010 -132643
rect -7954 -132651 -7910 -132643
rect -7854 -132651 -7810 -132643
rect -7354 -132651 -7310 -132643
rect -7254 -132651 -7210 -132643
rect -7154 -132651 -7110 -132643
rect -7054 -132651 -7010 -132643
rect -6954 -132651 -6910 -132643
rect -6854 -132651 -6810 -132643
rect -6754 -132651 -6710 -132643
rect -6654 -132651 -6610 -132643
rect -6554 -132651 -6510 -132643
rect -6454 -132651 -6410 -132643
rect -6354 -132651 -6310 -132643
rect -6254 -132651 -6210 -132643
rect -6154 -132651 -6110 -132643
rect -6054 -132651 -6010 -132643
rect -5954 -132651 -5910 -132643
rect -5854 -132651 -5810 -132643
rect -13310 -132695 -13302 -132651
rect -13210 -132695 -13202 -132651
rect -13110 -132695 -13102 -132651
rect -13010 -132695 -13002 -132651
rect -12910 -132695 -12902 -132651
rect -12810 -132695 -12802 -132651
rect -12710 -132695 -12702 -132651
rect -12610 -132695 -12602 -132651
rect -12510 -132695 -12502 -132651
rect -12410 -132695 -12402 -132651
rect -12310 -132695 -12302 -132651
rect -12210 -132695 -12202 -132651
rect -12110 -132695 -12102 -132651
rect -12010 -132695 -12002 -132651
rect -11910 -132695 -11902 -132651
rect -11810 -132695 -11802 -132651
rect -11310 -132695 -11302 -132651
rect -11210 -132695 -11202 -132651
rect -11110 -132695 -11102 -132651
rect -11010 -132695 -11002 -132651
rect -10910 -132695 -10902 -132651
rect -10810 -132695 -10802 -132651
rect -10710 -132695 -10702 -132651
rect -10610 -132695 -10602 -132651
rect -10510 -132695 -10502 -132651
rect -10410 -132695 -10402 -132651
rect -10310 -132695 -10302 -132651
rect -10210 -132695 -10202 -132651
rect -10110 -132695 -10102 -132651
rect -10010 -132695 -10002 -132651
rect -9910 -132695 -9902 -132651
rect -9810 -132695 -9802 -132651
rect -9310 -132695 -9302 -132651
rect -9210 -132695 -9202 -132651
rect -9110 -132695 -9102 -132651
rect -9010 -132695 -9002 -132651
rect -8910 -132695 -8902 -132651
rect -8810 -132695 -8802 -132651
rect -8710 -132695 -8702 -132651
rect -8610 -132695 -8602 -132651
rect -8510 -132695 -8502 -132651
rect -8410 -132695 -8402 -132651
rect -8310 -132695 -8302 -132651
rect -8210 -132695 -8202 -132651
rect -8110 -132695 -8102 -132651
rect -8010 -132695 -8002 -132651
rect -7910 -132695 -7902 -132651
rect -7810 -132695 -7802 -132651
rect -7310 -132695 -7302 -132651
rect -7210 -132695 -7202 -132651
rect -7110 -132695 -7102 -132651
rect -7010 -132695 -7002 -132651
rect -6910 -132695 -6902 -132651
rect -6810 -132695 -6802 -132651
rect -6710 -132695 -6702 -132651
rect -6610 -132695 -6602 -132651
rect -6510 -132695 -6502 -132651
rect -6410 -132695 -6402 -132651
rect -6310 -132695 -6302 -132651
rect -6210 -132695 -6202 -132651
rect -6110 -132695 -6102 -132651
rect -6010 -132695 -6002 -132651
rect -5910 -132695 -5902 -132651
rect -5810 -132695 -5802 -132651
rect 37387 -132685 37431 -132677
rect 37487 -132685 37531 -132677
rect 37587 -132685 37631 -132677
rect 37687 -132685 37731 -132677
rect 37787 -132685 37831 -132677
rect 37887 -132685 37931 -132677
rect 37987 -132685 38031 -132677
rect 38087 -132685 38131 -132677
rect 38187 -132685 38231 -132677
rect 38287 -132685 38331 -132677
rect 38387 -132685 38431 -132677
rect 38487 -132685 38531 -132677
rect 38587 -132685 38631 -132677
rect 38687 -132685 38731 -132677
rect 38787 -132685 38831 -132677
rect 38887 -132685 38931 -132677
rect 39387 -132685 39431 -132677
rect 39487 -132685 39531 -132677
rect 39587 -132685 39631 -132677
rect 39687 -132685 39731 -132677
rect 39787 -132685 39831 -132677
rect 39887 -132685 39931 -132677
rect 39987 -132685 40031 -132677
rect 40087 -132685 40131 -132677
rect 40187 -132685 40231 -132677
rect 40287 -132685 40331 -132677
rect 40387 -132685 40431 -132677
rect 40487 -132685 40531 -132677
rect 40587 -132685 40631 -132677
rect 40687 -132685 40731 -132677
rect 40787 -132685 40831 -132677
rect 40887 -132685 40931 -132677
rect 41387 -132685 41431 -132677
rect 41487 -132685 41531 -132677
rect 41587 -132685 41631 -132677
rect 41687 -132685 41731 -132677
rect 41787 -132685 41831 -132677
rect 41887 -132685 41931 -132677
rect 41987 -132685 42031 -132677
rect 42087 -132685 42131 -132677
rect 42187 -132685 42231 -132677
rect 42287 -132685 42331 -132677
rect 42387 -132685 42431 -132677
rect 42487 -132685 42531 -132677
rect 42587 -132685 42631 -132677
rect 42687 -132685 42731 -132677
rect 42787 -132685 42831 -132677
rect 42887 -132685 42931 -132677
rect 43387 -132685 43431 -132677
rect 43487 -132685 43531 -132677
rect 43587 -132685 43631 -132677
rect 43687 -132685 43731 -132677
rect 43787 -132685 43831 -132677
rect 43887 -132685 43931 -132677
rect 43987 -132685 44031 -132677
rect 44087 -132685 44131 -132677
rect 44187 -132685 44231 -132677
rect 44287 -132685 44331 -132677
rect 44387 -132685 44431 -132677
rect 44487 -132685 44531 -132677
rect 44587 -132685 44631 -132677
rect 44687 -132685 44731 -132677
rect 44787 -132685 44831 -132677
rect 44887 -132685 44931 -132677
rect 37431 -132729 37439 -132685
rect 37531 -132729 37539 -132685
rect 37631 -132729 37639 -132685
rect 37731 -132729 37739 -132685
rect 37831 -132729 37839 -132685
rect 37931 -132729 37939 -132685
rect 38031 -132729 38039 -132685
rect 38131 -132729 38139 -132685
rect 38231 -132729 38239 -132685
rect 38331 -132729 38339 -132685
rect 38431 -132729 38439 -132685
rect 38531 -132729 38539 -132685
rect 38631 -132729 38639 -132685
rect 38731 -132729 38739 -132685
rect 38831 -132729 38839 -132685
rect 38931 -132729 38939 -132685
rect 39431 -132729 39439 -132685
rect 39531 -132729 39539 -132685
rect 39631 -132729 39639 -132685
rect 39731 -132729 39739 -132685
rect 39831 -132729 39839 -132685
rect 39931 -132729 39939 -132685
rect 40031 -132729 40039 -132685
rect 40131 -132729 40139 -132685
rect 40231 -132729 40239 -132685
rect 40331 -132729 40339 -132685
rect 40431 -132729 40439 -132685
rect 40531 -132729 40539 -132685
rect 40631 -132729 40639 -132685
rect 40731 -132729 40739 -132685
rect 40831 -132729 40839 -132685
rect 40931 -132729 40939 -132685
rect 41431 -132729 41439 -132685
rect 41531 -132729 41539 -132685
rect 41631 -132729 41639 -132685
rect 41731 -132729 41739 -132685
rect 41831 -132729 41839 -132685
rect 41931 -132729 41939 -132685
rect 42031 -132729 42039 -132685
rect 42131 -132729 42139 -132685
rect 42231 -132729 42239 -132685
rect 42331 -132729 42339 -132685
rect 42431 -132729 42439 -132685
rect 42531 -132729 42539 -132685
rect 42631 -132729 42639 -132685
rect 42731 -132729 42739 -132685
rect 42831 -132729 42839 -132685
rect 42931 -132729 42939 -132685
rect 43431 -132729 43439 -132685
rect 43531 -132729 43539 -132685
rect 43631 -132729 43639 -132685
rect 43731 -132729 43739 -132685
rect 43831 -132729 43839 -132685
rect 43931 -132729 43939 -132685
rect 44031 -132729 44039 -132685
rect 44131 -132729 44139 -132685
rect 44231 -132729 44239 -132685
rect 44331 -132729 44339 -132685
rect 44431 -132729 44439 -132685
rect 44531 -132729 44539 -132685
rect 44631 -132729 44639 -132685
rect 44731 -132729 44739 -132685
rect 44831 -132729 44839 -132685
rect 44931 -132729 44939 -132685
rect -13354 -132751 -13310 -132743
rect -13254 -132751 -13210 -132743
rect -13154 -132751 -13110 -132743
rect -13054 -132751 -13010 -132743
rect -12954 -132751 -12910 -132743
rect -12854 -132751 -12810 -132743
rect -12754 -132751 -12710 -132743
rect -12654 -132751 -12610 -132743
rect -12554 -132751 -12510 -132743
rect -12454 -132751 -12410 -132743
rect -12354 -132751 -12310 -132743
rect -12254 -132751 -12210 -132743
rect -12154 -132751 -12110 -132743
rect -12054 -132751 -12010 -132743
rect -11954 -132751 -11910 -132743
rect -11854 -132751 -11810 -132743
rect -11354 -132751 -11310 -132743
rect -11254 -132751 -11210 -132743
rect -11154 -132751 -11110 -132743
rect -11054 -132751 -11010 -132743
rect -10954 -132751 -10910 -132743
rect -10854 -132751 -10810 -132743
rect -10754 -132751 -10710 -132743
rect -10654 -132751 -10610 -132743
rect -10554 -132751 -10510 -132743
rect -10454 -132751 -10410 -132743
rect -10354 -132751 -10310 -132743
rect -10254 -132751 -10210 -132743
rect -10154 -132751 -10110 -132743
rect -10054 -132751 -10010 -132743
rect -9954 -132751 -9910 -132743
rect -9854 -132751 -9810 -132743
rect -9354 -132751 -9310 -132743
rect -9254 -132751 -9210 -132743
rect -9154 -132751 -9110 -132743
rect -9054 -132751 -9010 -132743
rect -8954 -132751 -8910 -132743
rect -8854 -132751 -8810 -132743
rect -8754 -132751 -8710 -132743
rect -8654 -132751 -8610 -132743
rect -8554 -132751 -8510 -132743
rect -8454 -132751 -8410 -132743
rect -8354 -132751 -8310 -132743
rect -8254 -132751 -8210 -132743
rect -8154 -132751 -8110 -132743
rect -8054 -132751 -8010 -132743
rect -7954 -132751 -7910 -132743
rect -7854 -132751 -7810 -132743
rect -7354 -132751 -7310 -132743
rect -7254 -132751 -7210 -132743
rect -7154 -132751 -7110 -132743
rect -7054 -132751 -7010 -132743
rect -6954 -132751 -6910 -132743
rect -6854 -132751 -6810 -132743
rect -6754 -132751 -6710 -132743
rect -6654 -132751 -6610 -132743
rect -6554 -132751 -6510 -132743
rect -6454 -132751 -6410 -132743
rect -6354 -132751 -6310 -132743
rect -6254 -132751 -6210 -132743
rect -6154 -132751 -6110 -132743
rect -6054 -132751 -6010 -132743
rect -5954 -132751 -5910 -132743
rect -5854 -132751 -5810 -132743
rect -13310 -132795 -13302 -132751
rect -13210 -132795 -13202 -132751
rect -13110 -132795 -13102 -132751
rect -13010 -132795 -13002 -132751
rect -12910 -132795 -12902 -132751
rect -12810 -132795 -12802 -132751
rect -12710 -132795 -12702 -132751
rect -12610 -132795 -12602 -132751
rect -12510 -132795 -12502 -132751
rect -12410 -132795 -12402 -132751
rect -12310 -132795 -12302 -132751
rect -12210 -132795 -12202 -132751
rect -12110 -132795 -12102 -132751
rect -12010 -132795 -12002 -132751
rect -11910 -132795 -11902 -132751
rect -11810 -132795 -11802 -132751
rect -11310 -132795 -11302 -132751
rect -11210 -132795 -11202 -132751
rect -11110 -132795 -11102 -132751
rect -11010 -132795 -11002 -132751
rect -10910 -132795 -10902 -132751
rect -10810 -132795 -10802 -132751
rect -10710 -132795 -10702 -132751
rect -10610 -132795 -10602 -132751
rect -10510 -132795 -10502 -132751
rect -10410 -132795 -10402 -132751
rect -10310 -132795 -10302 -132751
rect -10210 -132795 -10202 -132751
rect -10110 -132795 -10102 -132751
rect -10010 -132795 -10002 -132751
rect -9910 -132795 -9902 -132751
rect -9810 -132795 -9802 -132751
rect -9310 -132795 -9302 -132751
rect -9210 -132795 -9202 -132751
rect -9110 -132795 -9102 -132751
rect -9010 -132795 -9002 -132751
rect -8910 -132795 -8902 -132751
rect -8810 -132795 -8802 -132751
rect -8710 -132795 -8702 -132751
rect -8610 -132795 -8602 -132751
rect -8510 -132795 -8502 -132751
rect -8410 -132795 -8402 -132751
rect -8310 -132795 -8302 -132751
rect -8210 -132795 -8202 -132751
rect -8110 -132795 -8102 -132751
rect -8010 -132795 -8002 -132751
rect -7910 -132795 -7902 -132751
rect -7810 -132795 -7802 -132751
rect -7310 -132795 -7302 -132751
rect -7210 -132795 -7202 -132751
rect -7110 -132795 -7102 -132751
rect -7010 -132795 -7002 -132751
rect -6910 -132795 -6902 -132751
rect -6810 -132795 -6802 -132751
rect -6710 -132795 -6702 -132751
rect -6610 -132795 -6602 -132751
rect -6510 -132795 -6502 -132751
rect -6410 -132795 -6402 -132751
rect -6310 -132795 -6302 -132751
rect -6210 -132795 -6202 -132751
rect -6110 -132795 -6102 -132751
rect -6010 -132795 -6002 -132751
rect -5910 -132795 -5902 -132751
rect -5810 -132795 -5802 -132751
rect 37387 -132785 37431 -132777
rect 37487 -132785 37531 -132777
rect 37587 -132785 37631 -132777
rect 37687 -132785 37731 -132777
rect 37787 -132785 37831 -132777
rect 37887 -132785 37931 -132777
rect 37987 -132785 38031 -132777
rect 38087 -132785 38131 -132777
rect 38187 -132785 38231 -132777
rect 38287 -132785 38331 -132777
rect 38387 -132785 38431 -132777
rect 38487 -132785 38531 -132777
rect 38587 -132785 38631 -132777
rect 38687 -132785 38731 -132777
rect 38787 -132785 38831 -132777
rect 38887 -132785 38931 -132777
rect 39387 -132785 39431 -132777
rect 39487 -132785 39531 -132777
rect 39587 -132785 39631 -132777
rect 39687 -132785 39731 -132777
rect 39787 -132785 39831 -132777
rect 39887 -132785 39931 -132777
rect 39987 -132785 40031 -132777
rect 40087 -132785 40131 -132777
rect 40187 -132785 40231 -132777
rect 40287 -132785 40331 -132777
rect 40387 -132785 40431 -132777
rect 40487 -132785 40531 -132777
rect 40587 -132785 40631 -132777
rect 40687 -132785 40731 -132777
rect 40787 -132785 40831 -132777
rect 40887 -132785 40931 -132777
rect 41387 -132785 41431 -132777
rect 41487 -132785 41531 -132777
rect 41587 -132785 41631 -132777
rect 41687 -132785 41731 -132777
rect 41787 -132785 41831 -132777
rect 41887 -132785 41931 -132777
rect 41987 -132785 42031 -132777
rect 42087 -132785 42131 -132777
rect 42187 -132785 42231 -132777
rect 42287 -132785 42331 -132777
rect 42387 -132785 42431 -132777
rect 42487 -132785 42531 -132777
rect 42587 -132785 42631 -132777
rect 42687 -132785 42731 -132777
rect 42787 -132785 42831 -132777
rect 42887 -132785 42931 -132777
rect 43387 -132785 43431 -132777
rect 43487 -132785 43531 -132777
rect 43587 -132785 43631 -132777
rect 43687 -132785 43731 -132777
rect 43787 -132785 43831 -132777
rect 43887 -132785 43931 -132777
rect 43987 -132785 44031 -132777
rect 44087 -132785 44131 -132777
rect 44187 -132785 44231 -132777
rect 44287 -132785 44331 -132777
rect 44387 -132785 44431 -132777
rect 44487 -132785 44531 -132777
rect 44587 -132785 44631 -132777
rect 44687 -132785 44731 -132777
rect 44787 -132785 44831 -132777
rect 44887 -132785 44931 -132777
rect 37431 -132829 37439 -132785
rect 37531 -132829 37539 -132785
rect 37631 -132829 37639 -132785
rect 37731 -132829 37739 -132785
rect 37831 -132829 37839 -132785
rect 37931 -132829 37939 -132785
rect 38031 -132829 38039 -132785
rect 38131 -132829 38139 -132785
rect 38231 -132829 38239 -132785
rect 38331 -132829 38339 -132785
rect 38431 -132829 38439 -132785
rect 38531 -132829 38539 -132785
rect 38631 -132829 38639 -132785
rect 38731 -132829 38739 -132785
rect 38831 -132829 38839 -132785
rect 38931 -132829 38939 -132785
rect 39431 -132829 39439 -132785
rect 39531 -132829 39539 -132785
rect 39631 -132829 39639 -132785
rect 39731 -132829 39739 -132785
rect 39831 -132829 39839 -132785
rect 39931 -132829 39939 -132785
rect 40031 -132829 40039 -132785
rect 40131 -132829 40139 -132785
rect 40231 -132829 40239 -132785
rect 40331 -132829 40339 -132785
rect 40431 -132829 40439 -132785
rect 40531 -132829 40539 -132785
rect 40631 -132829 40639 -132785
rect 40731 -132829 40739 -132785
rect 40831 -132829 40839 -132785
rect 40931 -132829 40939 -132785
rect 41431 -132829 41439 -132785
rect 41531 -132829 41539 -132785
rect 41631 -132829 41639 -132785
rect 41731 -132829 41739 -132785
rect 41831 -132829 41839 -132785
rect 41931 -132829 41939 -132785
rect 42031 -132829 42039 -132785
rect 42131 -132829 42139 -132785
rect 42231 -132829 42239 -132785
rect 42331 -132829 42339 -132785
rect 42431 -132829 42439 -132785
rect 42531 -132829 42539 -132785
rect 42631 -132829 42639 -132785
rect 42731 -132829 42739 -132785
rect 42831 -132829 42839 -132785
rect 42931 -132829 42939 -132785
rect 43431 -132829 43439 -132785
rect 43531 -132829 43539 -132785
rect 43631 -132829 43639 -132785
rect 43731 -132829 43739 -132785
rect 43831 -132829 43839 -132785
rect 43931 -132829 43939 -132785
rect 44031 -132829 44039 -132785
rect 44131 -132829 44139 -132785
rect 44231 -132829 44239 -132785
rect 44331 -132829 44339 -132785
rect 44431 -132829 44439 -132785
rect 44531 -132829 44539 -132785
rect 44631 -132829 44639 -132785
rect 44731 -132829 44739 -132785
rect 44831 -132829 44839 -132785
rect 44931 -132829 44939 -132785
rect 37387 -132885 37431 -132877
rect 37487 -132885 37531 -132877
rect 37587 -132885 37631 -132877
rect 37687 -132885 37731 -132877
rect 37787 -132885 37831 -132877
rect 37887 -132885 37931 -132877
rect 37987 -132885 38031 -132877
rect 38087 -132885 38131 -132877
rect 38187 -132885 38231 -132877
rect 38287 -132885 38331 -132877
rect 38387 -132885 38431 -132877
rect 38487 -132885 38531 -132877
rect 38587 -132885 38631 -132877
rect 38687 -132885 38731 -132877
rect 38787 -132885 38831 -132877
rect 38887 -132885 38931 -132877
rect 39387 -132885 39431 -132877
rect 39487 -132885 39531 -132877
rect 39587 -132885 39631 -132877
rect 39687 -132885 39731 -132877
rect 39787 -132885 39831 -132877
rect 39887 -132885 39931 -132877
rect 39987 -132885 40031 -132877
rect 40087 -132885 40131 -132877
rect 40187 -132885 40231 -132877
rect 40287 -132885 40331 -132877
rect 40387 -132885 40431 -132877
rect 40487 -132885 40531 -132877
rect 40587 -132885 40631 -132877
rect 40687 -132885 40731 -132877
rect 40787 -132885 40831 -132877
rect 40887 -132885 40931 -132877
rect 41387 -132885 41431 -132877
rect 41487 -132885 41531 -132877
rect 41587 -132885 41631 -132877
rect 41687 -132885 41731 -132877
rect 41787 -132885 41831 -132877
rect 41887 -132885 41931 -132877
rect 41987 -132885 42031 -132877
rect 42087 -132885 42131 -132877
rect 42187 -132885 42231 -132877
rect 42287 -132885 42331 -132877
rect 42387 -132885 42431 -132877
rect 42487 -132885 42531 -132877
rect 42587 -132885 42631 -132877
rect 42687 -132885 42731 -132877
rect 42787 -132885 42831 -132877
rect 42887 -132885 42931 -132877
rect 43387 -132885 43431 -132877
rect 43487 -132885 43531 -132877
rect 43587 -132885 43631 -132877
rect 43687 -132885 43731 -132877
rect 43787 -132885 43831 -132877
rect 43887 -132885 43931 -132877
rect 43987 -132885 44031 -132877
rect 44087 -132885 44131 -132877
rect 44187 -132885 44231 -132877
rect 44287 -132885 44331 -132877
rect 44387 -132885 44431 -132877
rect 44487 -132885 44531 -132877
rect 44587 -132885 44631 -132877
rect 44687 -132885 44731 -132877
rect 44787 -132885 44831 -132877
rect 44887 -132885 44931 -132877
rect 37431 -132929 37439 -132885
rect 37531 -132929 37539 -132885
rect 37631 -132929 37639 -132885
rect 37731 -132929 37739 -132885
rect 37831 -132929 37839 -132885
rect 37931 -132929 37939 -132885
rect 38031 -132929 38039 -132885
rect 38131 -132929 38139 -132885
rect 38231 -132929 38239 -132885
rect 38331 -132929 38339 -132885
rect 38431 -132929 38439 -132885
rect 38531 -132929 38539 -132885
rect 38631 -132929 38639 -132885
rect 38731 -132929 38739 -132885
rect 38831 -132929 38839 -132885
rect 38931 -132929 38939 -132885
rect 39431 -132929 39439 -132885
rect 39531 -132929 39539 -132885
rect 39631 -132929 39639 -132885
rect 39731 -132929 39739 -132885
rect 39831 -132929 39839 -132885
rect 39931 -132929 39939 -132885
rect 40031 -132929 40039 -132885
rect 40131 -132929 40139 -132885
rect 40231 -132929 40239 -132885
rect 40331 -132929 40339 -132885
rect 40431 -132929 40439 -132885
rect 40531 -132929 40539 -132885
rect 40631 -132929 40639 -132885
rect 40731 -132929 40739 -132885
rect 40831 -132929 40839 -132885
rect 40931 -132929 40939 -132885
rect 41431 -132929 41439 -132885
rect 41531 -132929 41539 -132885
rect 41631 -132929 41639 -132885
rect 41731 -132929 41739 -132885
rect 41831 -132929 41839 -132885
rect 41931 -132929 41939 -132885
rect 42031 -132929 42039 -132885
rect 42131 -132929 42139 -132885
rect 42231 -132929 42239 -132885
rect 42331 -132929 42339 -132885
rect 42431 -132929 42439 -132885
rect 42531 -132929 42539 -132885
rect 42631 -132929 42639 -132885
rect 42731 -132929 42739 -132885
rect 42831 -132929 42839 -132885
rect 42931 -132929 42939 -132885
rect 43431 -132929 43439 -132885
rect 43531 -132929 43539 -132885
rect 43631 -132929 43639 -132885
rect 43731 -132929 43739 -132885
rect 43831 -132929 43839 -132885
rect 43931 -132929 43939 -132885
rect 44031 -132929 44039 -132885
rect 44131 -132929 44139 -132885
rect 44231 -132929 44239 -132885
rect 44331 -132929 44339 -132885
rect 44431 -132929 44439 -132885
rect 44531 -132929 44539 -132885
rect 44631 -132929 44639 -132885
rect 44731 -132929 44739 -132885
rect 44831 -132929 44839 -132885
rect 44931 -132929 44939 -132885
rect -104783 -135314 -104739 -135306
rect -104683 -135314 -104639 -135306
rect -104583 -135314 -104539 -135306
rect -104483 -135314 -104439 -135306
rect -104383 -135314 -104339 -135306
rect -104283 -135314 -104239 -135306
rect -104183 -135314 -104139 -135306
rect -104083 -135314 -104039 -135306
rect -103983 -135314 -103939 -135306
rect -103883 -135314 -103839 -135306
rect -103783 -135314 -103739 -135306
rect -103683 -135314 -103639 -135306
rect -103583 -135314 -103539 -135306
rect -103483 -135314 -103439 -135306
rect -103383 -135314 -103339 -135306
rect -103283 -135314 -103239 -135306
rect -102783 -135314 -102739 -135306
rect -102683 -135314 -102639 -135306
rect -102583 -135314 -102539 -135306
rect -102483 -135314 -102439 -135306
rect -102383 -135314 -102339 -135306
rect -102283 -135314 -102239 -135306
rect -102183 -135314 -102139 -135306
rect -102083 -135314 -102039 -135306
rect -101983 -135314 -101939 -135306
rect -101883 -135314 -101839 -135306
rect -101783 -135314 -101739 -135306
rect -101683 -135314 -101639 -135306
rect -101583 -135314 -101539 -135306
rect -101483 -135314 -101439 -135306
rect -101383 -135314 -101339 -135306
rect -101283 -135314 -101239 -135306
rect -100783 -135314 -100739 -135306
rect -100683 -135314 -100639 -135306
rect -100583 -135314 -100539 -135306
rect -100483 -135314 -100439 -135306
rect -100383 -135314 -100339 -135306
rect -100283 -135314 -100239 -135306
rect -100183 -135314 -100139 -135306
rect -100083 -135314 -100039 -135306
rect -99983 -135314 -99939 -135306
rect -99883 -135314 -99839 -135306
rect -99783 -135314 -99739 -135306
rect -99683 -135314 -99639 -135306
rect -99583 -135314 -99539 -135306
rect -99483 -135314 -99439 -135306
rect -99383 -135314 -99339 -135306
rect -99283 -135314 -99239 -135306
rect -98783 -135314 -98739 -135306
rect -98683 -135314 -98639 -135306
rect -98583 -135314 -98539 -135306
rect -98483 -135314 -98439 -135306
rect -98383 -135314 -98339 -135306
rect -98283 -135314 -98239 -135306
rect -98183 -135314 -98139 -135306
rect -98083 -135314 -98039 -135306
rect -97983 -135314 -97939 -135306
rect -97883 -135314 -97839 -135306
rect -97783 -135314 -97739 -135306
rect -97683 -135314 -97639 -135306
rect -97583 -135314 -97539 -135306
rect -97483 -135314 -97439 -135306
rect -97383 -135314 -97339 -135306
rect -97283 -135314 -97239 -135306
rect -104739 -135358 -104731 -135314
rect -104639 -135358 -104631 -135314
rect -104539 -135358 -104531 -135314
rect -104439 -135358 -104431 -135314
rect -104339 -135358 -104331 -135314
rect -104239 -135358 -104231 -135314
rect -104139 -135358 -104131 -135314
rect -104039 -135358 -104031 -135314
rect -103939 -135358 -103931 -135314
rect -103839 -135358 -103831 -135314
rect -103739 -135358 -103731 -135314
rect -103639 -135358 -103631 -135314
rect -103539 -135358 -103531 -135314
rect -103439 -135358 -103431 -135314
rect -103339 -135358 -103331 -135314
rect -103239 -135358 -103231 -135314
rect -102739 -135358 -102731 -135314
rect -102639 -135358 -102631 -135314
rect -102539 -135358 -102531 -135314
rect -102439 -135358 -102431 -135314
rect -102339 -135358 -102331 -135314
rect -102239 -135358 -102231 -135314
rect -102139 -135358 -102131 -135314
rect -102039 -135358 -102031 -135314
rect -101939 -135358 -101931 -135314
rect -101839 -135358 -101831 -135314
rect -101739 -135358 -101731 -135314
rect -101639 -135358 -101631 -135314
rect -101539 -135358 -101531 -135314
rect -101439 -135358 -101431 -135314
rect -101339 -135358 -101331 -135314
rect -101239 -135358 -101231 -135314
rect -100739 -135358 -100731 -135314
rect -100639 -135358 -100631 -135314
rect -100539 -135358 -100531 -135314
rect -100439 -135358 -100431 -135314
rect -100339 -135358 -100331 -135314
rect -100239 -135358 -100231 -135314
rect -100139 -135358 -100131 -135314
rect -100039 -135358 -100031 -135314
rect -99939 -135358 -99931 -135314
rect -99839 -135358 -99831 -135314
rect -99739 -135358 -99731 -135314
rect -99639 -135358 -99631 -135314
rect -99539 -135358 -99531 -135314
rect -99439 -135358 -99431 -135314
rect -99339 -135358 -99331 -135314
rect -99239 -135358 -99231 -135314
rect -98739 -135358 -98731 -135314
rect -98639 -135358 -98631 -135314
rect -98539 -135358 -98531 -135314
rect -98439 -135358 -98431 -135314
rect -98339 -135358 -98331 -135314
rect -98239 -135358 -98231 -135314
rect -98139 -135358 -98131 -135314
rect -98039 -135358 -98031 -135314
rect -97939 -135358 -97931 -135314
rect -97839 -135358 -97831 -135314
rect -97739 -135358 -97731 -135314
rect -97639 -135358 -97631 -135314
rect -97539 -135358 -97531 -135314
rect -97439 -135358 -97431 -135314
rect -97339 -135358 -97331 -135314
rect -97239 -135358 -97231 -135314
rect -104783 -135414 -104739 -135406
rect -104683 -135414 -104639 -135406
rect -104583 -135414 -104539 -135406
rect -104483 -135414 -104439 -135406
rect -104383 -135414 -104339 -135406
rect -104283 -135414 -104239 -135406
rect -104183 -135414 -104139 -135406
rect -104083 -135414 -104039 -135406
rect -103983 -135414 -103939 -135406
rect -103883 -135414 -103839 -135406
rect -103783 -135414 -103739 -135406
rect -103683 -135414 -103639 -135406
rect -103583 -135414 -103539 -135406
rect -103483 -135414 -103439 -135406
rect -103383 -135414 -103339 -135406
rect -103283 -135414 -103239 -135406
rect -102783 -135414 -102739 -135406
rect -102683 -135414 -102639 -135406
rect -102583 -135414 -102539 -135406
rect -102483 -135414 -102439 -135406
rect -102383 -135414 -102339 -135406
rect -102283 -135414 -102239 -135406
rect -102183 -135414 -102139 -135406
rect -102083 -135414 -102039 -135406
rect -101983 -135414 -101939 -135406
rect -101883 -135414 -101839 -135406
rect -101783 -135414 -101739 -135406
rect -101683 -135414 -101639 -135406
rect -101583 -135414 -101539 -135406
rect -101483 -135414 -101439 -135406
rect -101383 -135414 -101339 -135406
rect -101283 -135414 -101239 -135406
rect -100783 -135414 -100739 -135406
rect -100683 -135414 -100639 -135406
rect -100583 -135414 -100539 -135406
rect -100483 -135414 -100439 -135406
rect -100383 -135414 -100339 -135406
rect -100283 -135414 -100239 -135406
rect -100183 -135414 -100139 -135406
rect -100083 -135414 -100039 -135406
rect -99983 -135414 -99939 -135406
rect -99883 -135414 -99839 -135406
rect -99783 -135414 -99739 -135406
rect -99683 -135414 -99639 -135406
rect -99583 -135414 -99539 -135406
rect -99483 -135414 -99439 -135406
rect -99383 -135414 -99339 -135406
rect -99283 -135414 -99239 -135406
rect -98783 -135414 -98739 -135406
rect -98683 -135414 -98639 -135406
rect -98583 -135414 -98539 -135406
rect -98483 -135414 -98439 -135406
rect -98383 -135414 -98339 -135406
rect -98283 -135414 -98239 -135406
rect -98183 -135414 -98139 -135406
rect -98083 -135414 -98039 -135406
rect -97983 -135414 -97939 -135406
rect -97883 -135414 -97839 -135406
rect -97783 -135414 -97739 -135406
rect -97683 -135414 -97639 -135406
rect -97583 -135414 -97539 -135406
rect -97483 -135414 -97439 -135406
rect -97383 -135414 -97339 -135406
rect -97283 -135414 -97239 -135406
rect -104739 -135458 -104731 -135414
rect -104639 -135458 -104631 -135414
rect -104539 -135458 -104531 -135414
rect -104439 -135458 -104431 -135414
rect -104339 -135458 -104331 -135414
rect -104239 -135458 -104231 -135414
rect -104139 -135458 -104131 -135414
rect -104039 -135458 -104031 -135414
rect -103939 -135458 -103931 -135414
rect -103839 -135458 -103831 -135414
rect -103739 -135458 -103731 -135414
rect -103639 -135458 -103631 -135414
rect -103539 -135458 -103531 -135414
rect -103439 -135458 -103431 -135414
rect -103339 -135458 -103331 -135414
rect -103239 -135458 -103231 -135414
rect -102739 -135458 -102731 -135414
rect -102639 -135458 -102631 -135414
rect -102539 -135458 -102531 -135414
rect -102439 -135458 -102431 -135414
rect -102339 -135458 -102331 -135414
rect -102239 -135458 -102231 -135414
rect -102139 -135458 -102131 -135414
rect -102039 -135458 -102031 -135414
rect -101939 -135458 -101931 -135414
rect -101839 -135458 -101831 -135414
rect -101739 -135458 -101731 -135414
rect -101639 -135458 -101631 -135414
rect -101539 -135458 -101531 -135414
rect -101439 -135458 -101431 -135414
rect -101339 -135458 -101331 -135414
rect -101239 -135458 -101231 -135414
rect -100739 -135458 -100731 -135414
rect -100639 -135458 -100631 -135414
rect -100539 -135458 -100531 -135414
rect -100439 -135458 -100431 -135414
rect -100339 -135458 -100331 -135414
rect -100239 -135458 -100231 -135414
rect -100139 -135458 -100131 -135414
rect -100039 -135458 -100031 -135414
rect -99939 -135458 -99931 -135414
rect -99839 -135458 -99831 -135414
rect -99739 -135458 -99731 -135414
rect -99639 -135458 -99631 -135414
rect -99539 -135458 -99531 -135414
rect -99439 -135458 -99431 -135414
rect -99339 -135458 -99331 -135414
rect -99239 -135458 -99231 -135414
rect -98739 -135458 -98731 -135414
rect -98639 -135458 -98631 -135414
rect -98539 -135458 -98531 -135414
rect -98439 -135458 -98431 -135414
rect -98339 -135458 -98331 -135414
rect -98239 -135458 -98231 -135414
rect -98139 -135458 -98131 -135414
rect -98039 -135458 -98031 -135414
rect -97939 -135458 -97931 -135414
rect -97839 -135458 -97831 -135414
rect -97739 -135458 -97731 -135414
rect -97639 -135458 -97631 -135414
rect -97539 -135458 -97531 -135414
rect -97439 -135458 -97431 -135414
rect -97339 -135458 -97331 -135414
rect -97239 -135458 -97231 -135414
rect -104783 -135514 -104739 -135506
rect -104683 -135514 -104639 -135506
rect -104583 -135514 -104539 -135506
rect -104483 -135514 -104439 -135506
rect -104383 -135514 -104339 -135506
rect -104283 -135514 -104239 -135506
rect -104183 -135514 -104139 -135506
rect -104083 -135514 -104039 -135506
rect -103983 -135514 -103939 -135506
rect -103883 -135514 -103839 -135506
rect -103783 -135514 -103739 -135506
rect -103683 -135514 -103639 -135506
rect -103583 -135514 -103539 -135506
rect -103483 -135514 -103439 -135506
rect -103383 -135514 -103339 -135506
rect -103283 -135514 -103239 -135506
rect -102783 -135514 -102739 -135506
rect -102683 -135514 -102639 -135506
rect -102583 -135514 -102539 -135506
rect -102483 -135514 -102439 -135506
rect -102383 -135514 -102339 -135506
rect -102283 -135514 -102239 -135506
rect -102183 -135514 -102139 -135506
rect -102083 -135514 -102039 -135506
rect -101983 -135514 -101939 -135506
rect -101883 -135514 -101839 -135506
rect -101783 -135514 -101739 -135506
rect -101683 -135514 -101639 -135506
rect -101583 -135514 -101539 -135506
rect -101483 -135514 -101439 -135506
rect -101383 -135514 -101339 -135506
rect -101283 -135514 -101239 -135506
rect -100783 -135514 -100739 -135506
rect -100683 -135514 -100639 -135506
rect -100583 -135514 -100539 -135506
rect -100483 -135514 -100439 -135506
rect -100383 -135514 -100339 -135506
rect -100283 -135514 -100239 -135506
rect -100183 -135514 -100139 -135506
rect -100083 -135514 -100039 -135506
rect -99983 -135514 -99939 -135506
rect -99883 -135514 -99839 -135506
rect -99783 -135514 -99739 -135506
rect -99683 -135514 -99639 -135506
rect -99583 -135514 -99539 -135506
rect -99483 -135514 -99439 -135506
rect -99383 -135514 -99339 -135506
rect -99283 -135514 -99239 -135506
rect -98783 -135514 -98739 -135506
rect -98683 -135514 -98639 -135506
rect -98583 -135514 -98539 -135506
rect -98483 -135514 -98439 -135506
rect -98383 -135514 -98339 -135506
rect -98283 -135514 -98239 -135506
rect -98183 -135514 -98139 -135506
rect -98083 -135514 -98039 -135506
rect -97983 -135514 -97939 -135506
rect -97883 -135514 -97839 -135506
rect -97783 -135514 -97739 -135506
rect -97683 -135514 -97639 -135506
rect -97583 -135514 -97539 -135506
rect -97483 -135514 -97439 -135506
rect -97383 -135514 -97339 -135506
rect -97283 -135514 -97239 -135506
rect -104739 -135558 -104731 -135514
rect -104639 -135558 -104631 -135514
rect -104539 -135558 -104531 -135514
rect -104439 -135558 -104431 -135514
rect -104339 -135558 -104331 -135514
rect -104239 -135558 -104231 -135514
rect -104139 -135558 -104131 -135514
rect -104039 -135558 -104031 -135514
rect -103939 -135558 -103931 -135514
rect -103839 -135558 -103831 -135514
rect -103739 -135558 -103731 -135514
rect -103639 -135558 -103631 -135514
rect -103539 -135558 -103531 -135514
rect -103439 -135558 -103431 -135514
rect -103339 -135558 -103331 -135514
rect -103239 -135558 -103231 -135514
rect -102739 -135558 -102731 -135514
rect -102639 -135558 -102631 -135514
rect -102539 -135558 -102531 -135514
rect -102439 -135558 -102431 -135514
rect -102339 -135558 -102331 -135514
rect -102239 -135558 -102231 -135514
rect -102139 -135558 -102131 -135514
rect -102039 -135558 -102031 -135514
rect -101939 -135558 -101931 -135514
rect -101839 -135558 -101831 -135514
rect -101739 -135558 -101731 -135514
rect -101639 -135558 -101631 -135514
rect -101539 -135558 -101531 -135514
rect -101439 -135558 -101431 -135514
rect -101339 -135558 -101331 -135514
rect -101239 -135558 -101231 -135514
rect -100739 -135558 -100731 -135514
rect -100639 -135558 -100631 -135514
rect -100539 -135558 -100531 -135514
rect -100439 -135558 -100431 -135514
rect -100339 -135558 -100331 -135514
rect -100239 -135558 -100231 -135514
rect -100139 -135558 -100131 -135514
rect -100039 -135558 -100031 -135514
rect -99939 -135558 -99931 -135514
rect -99839 -135558 -99831 -135514
rect -99739 -135558 -99731 -135514
rect -99639 -135558 -99631 -135514
rect -99539 -135558 -99531 -135514
rect -99439 -135558 -99431 -135514
rect -99339 -135558 -99331 -135514
rect -99239 -135558 -99231 -135514
rect -98739 -135558 -98731 -135514
rect -98639 -135558 -98631 -135514
rect -98539 -135558 -98531 -135514
rect -98439 -135558 -98431 -135514
rect -98339 -135558 -98331 -135514
rect -98239 -135558 -98231 -135514
rect -98139 -135558 -98131 -135514
rect -98039 -135558 -98031 -135514
rect -97939 -135558 -97931 -135514
rect -97839 -135558 -97831 -135514
rect -97739 -135558 -97731 -135514
rect -97639 -135558 -97631 -135514
rect -97539 -135558 -97531 -135514
rect -97439 -135558 -97431 -135514
rect -97339 -135558 -97331 -135514
rect -97239 -135558 -97231 -135514
rect -104783 -135614 -104739 -135606
rect -104683 -135614 -104639 -135606
rect -104583 -135614 -104539 -135606
rect -104483 -135614 -104439 -135606
rect -104383 -135614 -104339 -135606
rect -104283 -135614 -104239 -135606
rect -104183 -135614 -104139 -135606
rect -104083 -135614 -104039 -135606
rect -103983 -135614 -103939 -135606
rect -103883 -135614 -103839 -135606
rect -103783 -135614 -103739 -135606
rect -103683 -135614 -103639 -135606
rect -103583 -135614 -103539 -135606
rect -103483 -135614 -103439 -135606
rect -103383 -135614 -103339 -135606
rect -103283 -135614 -103239 -135606
rect -102783 -135614 -102739 -135606
rect -102683 -135614 -102639 -135606
rect -102583 -135614 -102539 -135606
rect -102483 -135614 -102439 -135606
rect -102383 -135614 -102339 -135606
rect -102283 -135614 -102239 -135606
rect -102183 -135614 -102139 -135606
rect -102083 -135614 -102039 -135606
rect -101983 -135614 -101939 -135606
rect -101883 -135614 -101839 -135606
rect -101783 -135614 -101739 -135606
rect -101683 -135614 -101639 -135606
rect -101583 -135614 -101539 -135606
rect -101483 -135614 -101439 -135606
rect -101383 -135614 -101339 -135606
rect -101283 -135614 -101239 -135606
rect -100783 -135614 -100739 -135606
rect -100683 -135614 -100639 -135606
rect -100583 -135614 -100539 -135606
rect -100483 -135614 -100439 -135606
rect -100383 -135614 -100339 -135606
rect -100283 -135614 -100239 -135606
rect -100183 -135614 -100139 -135606
rect -100083 -135614 -100039 -135606
rect -99983 -135614 -99939 -135606
rect -99883 -135614 -99839 -135606
rect -99783 -135614 -99739 -135606
rect -99683 -135614 -99639 -135606
rect -99583 -135614 -99539 -135606
rect -99483 -135614 -99439 -135606
rect -99383 -135614 -99339 -135606
rect -99283 -135614 -99239 -135606
rect -98783 -135614 -98739 -135606
rect -98683 -135614 -98639 -135606
rect -98583 -135614 -98539 -135606
rect -98483 -135614 -98439 -135606
rect -98383 -135614 -98339 -135606
rect -98283 -135614 -98239 -135606
rect -98183 -135614 -98139 -135606
rect -98083 -135614 -98039 -135606
rect -97983 -135614 -97939 -135606
rect -97883 -135614 -97839 -135606
rect -97783 -135614 -97739 -135606
rect -97683 -135614 -97639 -135606
rect -97583 -135614 -97539 -135606
rect -97483 -135614 -97439 -135606
rect -97383 -135614 -97339 -135606
rect -97283 -135614 -97239 -135606
rect -104739 -135658 -104731 -135614
rect -104639 -135658 -104631 -135614
rect -104539 -135658 -104531 -135614
rect -104439 -135658 -104431 -135614
rect -104339 -135658 -104331 -135614
rect -104239 -135658 -104231 -135614
rect -104139 -135658 -104131 -135614
rect -104039 -135658 -104031 -135614
rect -103939 -135658 -103931 -135614
rect -103839 -135658 -103831 -135614
rect -103739 -135658 -103731 -135614
rect -103639 -135658 -103631 -135614
rect -103539 -135658 -103531 -135614
rect -103439 -135658 -103431 -135614
rect -103339 -135658 -103331 -135614
rect -103239 -135658 -103231 -135614
rect -102739 -135658 -102731 -135614
rect -102639 -135658 -102631 -135614
rect -102539 -135658 -102531 -135614
rect -102439 -135658 -102431 -135614
rect -102339 -135658 -102331 -135614
rect -102239 -135658 -102231 -135614
rect -102139 -135658 -102131 -135614
rect -102039 -135658 -102031 -135614
rect -101939 -135658 -101931 -135614
rect -101839 -135658 -101831 -135614
rect -101739 -135658 -101731 -135614
rect -101639 -135658 -101631 -135614
rect -101539 -135658 -101531 -135614
rect -101439 -135658 -101431 -135614
rect -101339 -135658 -101331 -135614
rect -101239 -135658 -101231 -135614
rect -100739 -135658 -100731 -135614
rect -100639 -135658 -100631 -135614
rect -100539 -135658 -100531 -135614
rect -100439 -135658 -100431 -135614
rect -100339 -135658 -100331 -135614
rect -100239 -135658 -100231 -135614
rect -100139 -135658 -100131 -135614
rect -100039 -135658 -100031 -135614
rect -99939 -135658 -99931 -135614
rect -99839 -135658 -99831 -135614
rect -99739 -135658 -99731 -135614
rect -99639 -135658 -99631 -135614
rect -99539 -135658 -99531 -135614
rect -99439 -135658 -99431 -135614
rect -99339 -135658 -99331 -135614
rect -99239 -135658 -99231 -135614
rect -98739 -135658 -98731 -135614
rect -98639 -135658 -98631 -135614
rect -98539 -135658 -98531 -135614
rect -98439 -135658 -98431 -135614
rect -98339 -135658 -98331 -135614
rect -98239 -135658 -98231 -135614
rect -98139 -135658 -98131 -135614
rect -98039 -135658 -98031 -135614
rect -97939 -135658 -97931 -135614
rect -97839 -135658 -97831 -135614
rect -97739 -135658 -97731 -135614
rect -97639 -135658 -97631 -135614
rect -97539 -135658 -97531 -135614
rect -97439 -135658 -97431 -135614
rect -97339 -135658 -97331 -135614
rect -97239 -135658 -97231 -135614
rect -104783 -135714 -104739 -135706
rect -104683 -135714 -104639 -135706
rect -104583 -135714 -104539 -135706
rect -104483 -135714 -104439 -135706
rect -104383 -135714 -104339 -135706
rect -104283 -135714 -104239 -135706
rect -104183 -135714 -104139 -135706
rect -104083 -135714 -104039 -135706
rect -103983 -135714 -103939 -135706
rect -103883 -135714 -103839 -135706
rect -103783 -135714 -103739 -135706
rect -103683 -135714 -103639 -135706
rect -103583 -135714 -103539 -135706
rect -103483 -135714 -103439 -135706
rect -103383 -135714 -103339 -135706
rect -103283 -135714 -103239 -135706
rect -102783 -135714 -102739 -135706
rect -102683 -135714 -102639 -135706
rect -102583 -135714 -102539 -135706
rect -102483 -135714 -102439 -135706
rect -102383 -135714 -102339 -135706
rect -102283 -135714 -102239 -135706
rect -102183 -135714 -102139 -135706
rect -102083 -135714 -102039 -135706
rect -101983 -135714 -101939 -135706
rect -101883 -135714 -101839 -135706
rect -101783 -135714 -101739 -135706
rect -101683 -135714 -101639 -135706
rect -101583 -135714 -101539 -135706
rect -101483 -135714 -101439 -135706
rect -101383 -135714 -101339 -135706
rect -101283 -135714 -101239 -135706
rect -100783 -135714 -100739 -135706
rect -100683 -135714 -100639 -135706
rect -100583 -135714 -100539 -135706
rect -100483 -135714 -100439 -135706
rect -100383 -135714 -100339 -135706
rect -100283 -135714 -100239 -135706
rect -100183 -135714 -100139 -135706
rect -100083 -135714 -100039 -135706
rect -99983 -135714 -99939 -135706
rect -99883 -135714 -99839 -135706
rect -99783 -135714 -99739 -135706
rect -99683 -135714 -99639 -135706
rect -99583 -135714 -99539 -135706
rect -99483 -135714 -99439 -135706
rect -99383 -135714 -99339 -135706
rect -99283 -135714 -99239 -135706
rect -98783 -135714 -98739 -135706
rect -98683 -135714 -98639 -135706
rect -98583 -135714 -98539 -135706
rect -98483 -135714 -98439 -135706
rect -98383 -135714 -98339 -135706
rect -98283 -135714 -98239 -135706
rect -98183 -135714 -98139 -135706
rect -98083 -135714 -98039 -135706
rect -97983 -135714 -97939 -135706
rect -97883 -135714 -97839 -135706
rect -97783 -135714 -97739 -135706
rect -97683 -135714 -97639 -135706
rect -97583 -135714 -97539 -135706
rect -97483 -135714 -97439 -135706
rect -97383 -135714 -97339 -135706
rect -97283 -135714 -97239 -135706
rect -104739 -135758 -104731 -135714
rect -104639 -135758 -104631 -135714
rect -104539 -135758 -104531 -135714
rect -104439 -135758 -104431 -135714
rect -104339 -135758 -104331 -135714
rect -104239 -135758 -104231 -135714
rect -104139 -135758 -104131 -135714
rect -104039 -135758 -104031 -135714
rect -103939 -135758 -103931 -135714
rect -103839 -135758 -103831 -135714
rect -103739 -135758 -103731 -135714
rect -103639 -135758 -103631 -135714
rect -103539 -135758 -103531 -135714
rect -103439 -135758 -103431 -135714
rect -103339 -135758 -103331 -135714
rect -103239 -135758 -103231 -135714
rect -102739 -135758 -102731 -135714
rect -102639 -135758 -102631 -135714
rect -102539 -135758 -102531 -135714
rect -102439 -135758 -102431 -135714
rect -102339 -135758 -102331 -135714
rect -102239 -135758 -102231 -135714
rect -102139 -135758 -102131 -135714
rect -102039 -135758 -102031 -135714
rect -101939 -135758 -101931 -135714
rect -101839 -135758 -101831 -135714
rect -101739 -135758 -101731 -135714
rect -101639 -135758 -101631 -135714
rect -101539 -135758 -101531 -135714
rect -101439 -135758 -101431 -135714
rect -101339 -135758 -101331 -135714
rect -101239 -135758 -101231 -135714
rect -100739 -135758 -100731 -135714
rect -100639 -135758 -100631 -135714
rect -100539 -135758 -100531 -135714
rect -100439 -135758 -100431 -135714
rect -100339 -135758 -100331 -135714
rect -100239 -135758 -100231 -135714
rect -100139 -135758 -100131 -135714
rect -100039 -135758 -100031 -135714
rect -99939 -135758 -99931 -135714
rect -99839 -135758 -99831 -135714
rect -99739 -135758 -99731 -135714
rect -99639 -135758 -99631 -135714
rect -99539 -135758 -99531 -135714
rect -99439 -135758 -99431 -135714
rect -99339 -135758 -99331 -135714
rect -99239 -135758 -99231 -135714
rect -98739 -135758 -98731 -135714
rect -98639 -135758 -98631 -135714
rect -98539 -135758 -98531 -135714
rect -98439 -135758 -98431 -135714
rect -98339 -135758 -98331 -135714
rect -98239 -135758 -98231 -135714
rect -98139 -135758 -98131 -135714
rect -98039 -135758 -98031 -135714
rect -97939 -135758 -97931 -135714
rect -97839 -135758 -97831 -135714
rect -97739 -135758 -97731 -135714
rect -97639 -135758 -97631 -135714
rect -97539 -135758 -97531 -135714
rect -97439 -135758 -97431 -135714
rect -97339 -135758 -97331 -135714
rect -97239 -135758 -97231 -135714
rect -104783 -135814 -104739 -135806
rect -104683 -135814 -104639 -135806
rect -104583 -135814 -104539 -135806
rect -104483 -135814 -104439 -135806
rect -104383 -135814 -104339 -135806
rect -104283 -135814 -104239 -135806
rect -104183 -135814 -104139 -135806
rect -104083 -135814 -104039 -135806
rect -103983 -135814 -103939 -135806
rect -103883 -135814 -103839 -135806
rect -103783 -135814 -103739 -135806
rect -103683 -135814 -103639 -135806
rect -103583 -135814 -103539 -135806
rect -103483 -135814 -103439 -135806
rect -103383 -135814 -103339 -135806
rect -103283 -135814 -103239 -135806
rect -102783 -135814 -102739 -135806
rect -102683 -135814 -102639 -135806
rect -102583 -135814 -102539 -135806
rect -102483 -135814 -102439 -135806
rect -102383 -135814 -102339 -135806
rect -102283 -135814 -102239 -135806
rect -102183 -135814 -102139 -135806
rect -102083 -135814 -102039 -135806
rect -101983 -135814 -101939 -135806
rect -101883 -135814 -101839 -135806
rect -101783 -135814 -101739 -135806
rect -101683 -135814 -101639 -135806
rect -101583 -135814 -101539 -135806
rect -101483 -135814 -101439 -135806
rect -101383 -135814 -101339 -135806
rect -101283 -135814 -101239 -135806
rect -100783 -135814 -100739 -135806
rect -100683 -135814 -100639 -135806
rect -100583 -135814 -100539 -135806
rect -100483 -135814 -100439 -135806
rect -100383 -135814 -100339 -135806
rect -100283 -135814 -100239 -135806
rect -100183 -135814 -100139 -135806
rect -100083 -135814 -100039 -135806
rect -99983 -135814 -99939 -135806
rect -99883 -135814 -99839 -135806
rect -99783 -135814 -99739 -135806
rect -99683 -135814 -99639 -135806
rect -99583 -135814 -99539 -135806
rect -99483 -135814 -99439 -135806
rect -99383 -135814 -99339 -135806
rect -99283 -135814 -99239 -135806
rect -98783 -135814 -98739 -135806
rect -98683 -135814 -98639 -135806
rect -98583 -135814 -98539 -135806
rect -98483 -135814 -98439 -135806
rect -98383 -135814 -98339 -135806
rect -98283 -135814 -98239 -135806
rect -98183 -135814 -98139 -135806
rect -98083 -135814 -98039 -135806
rect -97983 -135814 -97939 -135806
rect -97883 -135814 -97839 -135806
rect -97783 -135814 -97739 -135806
rect -97683 -135814 -97639 -135806
rect -97583 -135814 -97539 -135806
rect -97483 -135814 -97439 -135806
rect -97383 -135814 -97339 -135806
rect -97283 -135814 -97239 -135806
rect -104739 -135858 -104731 -135814
rect -104639 -135858 -104631 -135814
rect -104539 -135858 -104531 -135814
rect -104439 -135858 -104431 -135814
rect -104339 -135858 -104331 -135814
rect -104239 -135858 -104231 -135814
rect -104139 -135858 -104131 -135814
rect -104039 -135858 -104031 -135814
rect -103939 -135858 -103931 -135814
rect -103839 -135858 -103831 -135814
rect -103739 -135858 -103731 -135814
rect -103639 -135858 -103631 -135814
rect -103539 -135858 -103531 -135814
rect -103439 -135858 -103431 -135814
rect -103339 -135858 -103331 -135814
rect -103239 -135858 -103231 -135814
rect -102739 -135858 -102731 -135814
rect -102639 -135858 -102631 -135814
rect -102539 -135858 -102531 -135814
rect -102439 -135858 -102431 -135814
rect -102339 -135858 -102331 -135814
rect -102239 -135858 -102231 -135814
rect -102139 -135858 -102131 -135814
rect -102039 -135858 -102031 -135814
rect -101939 -135858 -101931 -135814
rect -101839 -135858 -101831 -135814
rect -101739 -135858 -101731 -135814
rect -101639 -135858 -101631 -135814
rect -101539 -135858 -101531 -135814
rect -101439 -135858 -101431 -135814
rect -101339 -135858 -101331 -135814
rect -101239 -135858 -101231 -135814
rect -100739 -135858 -100731 -135814
rect -100639 -135858 -100631 -135814
rect -100539 -135858 -100531 -135814
rect -100439 -135858 -100431 -135814
rect -100339 -135858 -100331 -135814
rect -100239 -135858 -100231 -135814
rect -100139 -135858 -100131 -135814
rect -100039 -135858 -100031 -135814
rect -99939 -135858 -99931 -135814
rect -99839 -135858 -99831 -135814
rect -99739 -135858 -99731 -135814
rect -99639 -135858 -99631 -135814
rect -99539 -135858 -99531 -135814
rect -99439 -135858 -99431 -135814
rect -99339 -135858 -99331 -135814
rect -99239 -135858 -99231 -135814
rect -98739 -135858 -98731 -135814
rect -98639 -135858 -98631 -135814
rect -98539 -135858 -98531 -135814
rect -98439 -135858 -98431 -135814
rect -98339 -135858 -98331 -135814
rect -98239 -135858 -98231 -135814
rect -98139 -135858 -98131 -135814
rect -98039 -135858 -98031 -135814
rect -97939 -135858 -97931 -135814
rect -97839 -135858 -97831 -135814
rect -97739 -135858 -97731 -135814
rect -97639 -135858 -97631 -135814
rect -97539 -135858 -97531 -135814
rect -97439 -135858 -97431 -135814
rect -97339 -135858 -97331 -135814
rect -97239 -135858 -97231 -135814
rect -104783 -135914 -104739 -135906
rect -104683 -135914 -104639 -135906
rect -104583 -135914 -104539 -135906
rect -104483 -135914 -104439 -135906
rect -104383 -135914 -104339 -135906
rect -104283 -135914 -104239 -135906
rect -104183 -135914 -104139 -135906
rect -104083 -135914 -104039 -135906
rect -103983 -135914 -103939 -135906
rect -103883 -135914 -103839 -135906
rect -103783 -135914 -103739 -135906
rect -103683 -135914 -103639 -135906
rect -103583 -135914 -103539 -135906
rect -103483 -135914 -103439 -135906
rect -103383 -135914 -103339 -135906
rect -103283 -135914 -103239 -135906
rect -102783 -135914 -102739 -135906
rect -102683 -135914 -102639 -135906
rect -102583 -135914 -102539 -135906
rect -102483 -135914 -102439 -135906
rect -102383 -135914 -102339 -135906
rect -102283 -135914 -102239 -135906
rect -102183 -135914 -102139 -135906
rect -102083 -135914 -102039 -135906
rect -101983 -135914 -101939 -135906
rect -101883 -135914 -101839 -135906
rect -101783 -135914 -101739 -135906
rect -101683 -135914 -101639 -135906
rect -101583 -135914 -101539 -135906
rect -101483 -135914 -101439 -135906
rect -101383 -135914 -101339 -135906
rect -101283 -135914 -101239 -135906
rect -100783 -135914 -100739 -135906
rect -100683 -135914 -100639 -135906
rect -100583 -135914 -100539 -135906
rect -100483 -135914 -100439 -135906
rect -100383 -135914 -100339 -135906
rect -100283 -135914 -100239 -135906
rect -100183 -135914 -100139 -135906
rect -100083 -135914 -100039 -135906
rect -99983 -135914 -99939 -135906
rect -99883 -135914 -99839 -135906
rect -99783 -135914 -99739 -135906
rect -99683 -135914 -99639 -135906
rect -99583 -135914 -99539 -135906
rect -99483 -135914 -99439 -135906
rect -99383 -135914 -99339 -135906
rect -99283 -135914 -99239 -135906
rect -98783 -135914 -98739 -135906
rect -98683 -135914 -98639 -135906
rect -98583 -135914 -98539 -135906
rect -98483 -135914 -98439 -135906
rect -98383 -135914 -98339 -135906
rect -98283 -135914 -98239 -135906
rect -98183 -135914 -98139 -135906
rect -98083 -135914 -98039 -135906
rect -97983 -135914 -97939 -135906
rect -97883 -135914 -97839 -135906
rect -97783 -135914 -97739 -135906
rect -97683 -135914 -97639 -135906
rect -97583 -135914 -97539 -135906
rect -97483 -135914 -97439 -135906
rect -97383 -135914 -97339 -135906
rect -97283 -135914 -97239 -135906
rect -104739 -135958 -104731 -135914
rect -104639 -135958 -104631 -135914
rect -104539 -135958 -104531 -135914
rect -104439 -135958 -104431 -135914
rect -104339 -135958 -104331 -135914
rect -104239 -135958 -104231 -135914
rect -104139 -135958 -104131 -135914
rect -104039 -135958 -104031 -135914
rect -103939 -135958 -103931 -135914
rect -103839 -135958 -103831 -135914
rect -103739 -135958 -103731 -135914
rect -103639 -135958 -103631 -135914
rect -103539 -135958 -103531 -135914
rect -103439 -135958 -103431 -135914
rect -103339 -135958 -103331 -135914
rect -103239 -135958 -103231 -135914
rect -102739 -135958 -102731 -135914
rect -102639 -135958 -102631 -135914
rect -102539 -135958 -102531 -135914
rect -102439 -135958 -102431 -135914
rect -102339 -135958 -102331 -135914
rect -102239 -135958 -102231 -135914
rect -102139 -135958 -102131 -135914
rect -102039 -135958 -102031 -135914
rect -101939 -135958 -101931 -135914
rect -101839 -135958 -101831 -135914
rect -101739 -135958 -101731 -135914
rect -101639 -135958 -101631 -135914
rect -101539 -135958 -101531 -135914
rect -101439 -135958 -101431 -135914
rect -101339 -135958 -101331 -135914
rect -101239 -135958 -101231 -135914
rect -100739 -135958 -100731 -135914
rect -100639 -135958 -100631 -135914
rect -100539 -135958 -100531 -135914
rect -100439 -135958 -100431 -135914
rect -100339 -135958 -100331 -135914
rect -100239 -135958 -100231 -135914
rect -100139 -135958 -100131 -135914
rect -100039 -135958 -100031 -135914
rect -99939 -135958 -99931 -135914
rect -99839 -135958 -99831 -135914
rect -99739 -135958 -99731 -135914
rect -99639 -135958 -99631 -135914
rect -99539 -135958 -99531 -135914
rect -99439 -135958 -99431 -135914
rect -99339 -135958 -99331 -135914
rect -99239 -135958 -99231 -135914
rect -98739 -135958 -98731 -135914
rect -98639 -135958 -98631 -135914
rect -98539 -135958 -98531 -135914
rect -98439 -135958 -98431 -135914
rect -98339 -135958 -98331 -135914
rect -98239 -135958 -98231 -135914
rect -98139 -135958 -98131 -135914
rect -98039 -135958 -98031 -135914
rect -97939 -135958 -97931 -135914
rect -97839 -135958 -97831 -135914
rect -97739 -135958 -97731 -135914
rect -97639 -135958 -97631 -135914
rect -97539 -135958 -97531 -135914
rect -97439 -135958 -97431 -135914
rect -97339 -135958 -97331 -135914
rect -97239 -135958 -97231 -135914
rect -104783 -136014 -104739 -136006
rect -104683 -136014 -104639 -136006
rect -104583 -136014 -104539 -136006
rect -104483 -136014 -104439 -136006
rect -104383 -136014 -104339 -136006
rect -104283 -136014 -104239 -136006
rect -104183 -136014 -104139 -136006
rect -104083 -136014 -104039 -136006
rect -103983 -136014 -103939 -136006
rect -103883 -136014 -103839 -136006
rect -103783 -136014 -103739 -136006
rect -103683 -136014 -103639 -136006
rect -103583 -136014 -103539 -136006
rect -103483 -136014 -103439 -136006
rect -103383 -136014 -103339 -136006
rect -103283 -136014 -103239 -136006
rect -102783 -136014 -102739 -136006
rect -102683 -136014 -102639 -136006
rect -102583 -136014 -102539 -136006
rect -102483 -136014 -102439 -136006
rect -102383 -136014 -102339 -136006
rect -102283 -136014 -102239 -136006
rect -102183 -136014 -102139 -136006
rect -102083 -136014 -102039 -136006
rect -101983 -136014 -101939 -136006
rect -101883 -136014 -101839 -136006
rect -101783 -136014 -101739 -136006
rect -101683 -136014 -101639 -136006
rect -101583 -136014 -101539 -136006
rect -101483 -136014 -101439 -136006
rect -101383 -136014 -101339 -136006
rect -101283 -136014 -101239 -136006
rect -100783 -136014 -100739 -136006
rect -100683 -136014 -100639 -136006
rect -100583 -136014 -100539 -136006
rect -100483 -136014 -100439 -136006
rect -100383 -136014 -100339 -136006
rect -100283 -136014 -100239 -136006
rect -100183 -136014 -100139 -136006
rect -100083 -136014 -100039 -136006
rect -99983 -136014 -99939 -136006
rect -99883 -136014 -99839 -136006
rect -99783 -136014 -99739 -136006
rect -99683 -136014 -99639 -136006
rect -99583 -136014 -99539 -136006
rect -99483 -136014 -99439 -136006
rect -99383 -136014 -99339 -136006
rect -99283 -136014 -99239 -136006
rect -98783 -136014 -98739 -136006
rect -98683 -136014 -98639 -136006
rect -98583 -136014 -98539 -136006
rect -98483 -136014 -98439 -136006
rect -98383 -136014 -98339 -136006
rect -98283 -136014 -98239 -136006
rect -98183 -136014 -98139 -136006
rect -98083 -136014 -98039 -136006
rect -97983 -136014 -97939 -136006
rect -97883 -136014 -97839 -136006
rect -97783 -136014 -97739 -136006
rect -97683 -136014 -97639 -136006
rect -97583 -136014 -97539 -136006
rect -97483 -136014 -97439 -136006
rect -97383 -136014 -97339 -136006
rect -97283 -136014 -97239 -136006
rect -104739 -136058 -104731 -136014
rect -104639 -136058 -104631 -136014
rect -104539 -136058 -104531 -136014
rect -104439 -136058 -104431 -136014
rect -104339 -136058 -104331 -136014
rect -104239 -136058 -104231 -136014
rect -104139 -136058 -104131 -136014
rect -104039 -136058 -104031 -136014
rect -103939 -136058 -103931 -136014
rect -103839 -136058 -103831 -136014
rect -103739 -136058 -103731 -136014
rect -103639 -136058 -103631 -136014
rect -103539 -136058 -103531 -136014
rect -103439 -136058 -103431 -136014
rect -103339 -136058 -103331 -136014
rect -103239 -136058 -103231 -136014
rect -102739 -136058 -102731 -136014
rect -102639 -136058 -102631 -136014
rect -102539 -136058 -102531 -136014
rect -102439 -136058 -102431 -136014
rect -102339 -136058 -102331 -136014
rect -102239 -136058 -102231 -136014
rect -102139 -136058 -102131 -136014
rect -102039 -136058 -102031 -136014
rect -101939 -136058 -101931 -136014
rect -101839 -136058 -101831 -136014
rect -101739 -136058 -101731 -136014
rect -101639 -136058 -101631 -136014
rect -101539 -136058 -101531 -136014
rect -101439 -136058 -101431 -136014
rect -101339 -136058 -101331 -136014
rect -101239 -136058 -101231 -136014
rect -100739 -136058 -100731 -136014
rect -100639 -136058 -100631 -136014
rect -100539 -136058 -100531 -136014
rect -100439 -136058 -100431 -136014
rect -100339 -136058 -100331 -136014
rect -100239 -136058 -100231 -136014
rect -100139 -136058 -100131 -136014
rect -100039 -136058 -100031 -136014
rect -99939 -136058 -99931 -136014
rect -99839 -136058 -99831 -136014
rect -99739 -136058 -99731 -136014
rect -99639 -136058 -99631 -136014
rect -99539 -136058 -99531 -136014
rect -99439 -136058 -99431 -136014
rect -99339 -136058 -99331 -136014
rect -99239 -136058 -99231 -136014
rect -98739 -136058 -98731 -136014
rect -98639 -136058 -98631 -136014
rect -98539 -136058 -98531 -136014
rect -98439 -136058 -98431 -136014
rect -98339 -136058 -98331 -136014
rect -98239 -136058 -98231 -136014
rect -98139 -136058 -98131 -136014
rect -98039 -136058 -98031 -136014
rect -97939 -136058 -97931 -136014
rect -97839 -136058 -97831 -136014
rect -97739 -136058 -97731 -136014
rect -97639 -136058 -97631 -136014
rect -97539 -136058 -97531 -136014
rect -97439 -136058 -97431 -136014
rect -97339 -136058 -97331 -136014
rect -97239 -136058 -97231 -136014
rect -104783 -136114 -104739 -136106
rect -104683 -136114 -104639 -136106
rect -104583 -136114 -104539 -136106
rect -104483 -136114 -104439 -136106
rect -104383 -136114 -104339 -136106
rect -104283 -136114 -104239 -136106
rect -104183 -136114 -104139 -136106
rect -104083 -136114 -104039 -136106
rect -103983 -136114 -103939 -136106
rect -103883 -136114 -103839 -136106
rect -103783 -136114 -103739 -136106
rect -103683 -136114 -103639 -136106
rect -103583 -136114 -103539 -136106
rect -103483 -136114 -103439 -136106
rect -103383 -136114 -103339 -136106
rect -103283 -136114 -103239 -136106
rect -102783 -136114 -102739 -136106
rect -102683 -136114 -102639 -136106
rect -102583 -136114 -102539 -136106
rect -102483 -136114 -102439 -136106
rect -102383 -136114 -102339 -136106
rect -102283 -136114 -102239 -136106
rect -102183 -136114 -102139 -136106
rect -102083 -136114 -102039 -136106
rect -101983 -136114 -101939 -136106
rect -101883 -136114 -101839 -136106
rect -101783 -136114 -101739 -136106
rect -101683 -136114 -101639 -136106
rect -101583 -136114 -101539 -136106
rect -101483 -136114 -101439 -136106
rect -101383 -136114 -101339 -136106
rect -101283 -136114 -101239 -136106
rect -100783 -136114 -100739 -136106
rect -100683 -136114 -100639 -136106
rect -100583 -136114 -100539 -136106
rect -100483 -136114 -100439 -136106
rect -100383 -136114 -100339 -136106
rect -100283 -136114 -100239 -136106
rect -100183 -136114 -100139 -136106
rect -100083 -136114 -100039 -136106
rect -99983 -136114 -99939 -136106
rect -99883 -136114 -99839 -136106
rect -99783 -136114 -99739 -136106
rect -99683 -136114 -99639 -136106
rect -99583 -136114 -99539 -136106
rect -99483 -136114 -99439 -136106
rect -99383 -136114 -99339 -136106
rect -99283 -136114 -99239 -136106
rect -98783 -136114 -98739 -136106
rect -98683 -136114 -98639 -136106
rect -98583 -136114 -98539 -136106
rect -98483 -136114 -98439 -136106
rect -98383 -136114 -98339 -136106
rect -98283 -136114 -98239 -136106
rect -98183 -136114 -98139 -136106
rect -98083 -136114 -98039 -136106
rect -97983 -136114 -97939 -136106
rect -97883 -136114 -97839 -136106
rect -97783 -136114 -97739 -136106
rect -97683 -136114 -97639 -136106
rect -97583 -136114 -97539 -136106
rect -97483 -136114 -97439 -136106
rect -97383 -136114 -97339 -136106
rect -97283 -136114 -97239 -136106
rect -104739 -136158 -104731 -136114
rect -104639 -136158 -104631 -136114
rect -104539 -136158 -104531 -136114
rect -104439 -136158 -104431 -136114
rect -104339 -136158 -104331 -136114
rect -104239 -136158 -104231 -136114
rect -104139 -136158 -104131 -136114
rect -104039 -136158 -104031 -136114
rect -103939 -136158 -103931 -136114
rect -103839 -136158 -103831 -136114
rect -103739 -136158 -103731 -136114
rect -103639 -136158 -103631 -136114
rect -103539 -136158 -103531 -136114
rect -103439 -136158 -103431 -136114
rect -103339 -136158 -103331 -136114
rect -103239 -136158 -103231 -136114
rect -102739 -136158 -102731 -136114
rect -102639 -136158 -102631 -136114
rect -102539 -136158 -102531 -136114
rect -102439 -136158 -102431 -136114
rect -102339 -136158 -102331 -136114
rect -102239 -136158 -102231 -136114
rect -102139 -136158 -102131 -136114
rect -102039 -136158 -102031 -136114
rect -101939 -136158 -101931 -136114
rect -101839 -136158 -101831 -136114
rect -101739 -136158 -101731 -136114
rect -101639 -136158 -101631 -136114
rect -101539 -136158 -101531 -136114
rect -101439 -136158 -101431 -136114
rect -101339 -136158 -101331 -136114
rect -101239 -136158 -101231 -136114
rect -100739 -136158 -100731 -136114
rect -100639 -136158 -100631 -136114
rect -100539 -136158 -100531 -136114
rect -100439 -136158 -100431 -136114
rect -100339 -136158 -100331 -136114
rect -100239 -136158 -100231 -136114
rect -100139 -136158 -100131 -136114
rect -100039 -136158 -100031 -136114
rect -99939 -136158 -99931 -136114
rect -99839 -136158 -99831 -136114
rect -99739 -136158 -99731 -136114
rect -99639 -136158 -99631 -136114
rect -99539 -136158 -99531 -136114
rect -99439 -136158 -99431 -136114
rect -99339 -136158 -99331 -136114
rect -99239 -136158 -99231 -136114
rect -98739 -136158 -98731 -136114
rect -98639 -136158 -98631 -136114
rect -98539 -136158 -98531 -136114
rect -98439 -136158 -98431 -136114
rect -98339 -136158 -98331 -136114
rect -98239 -136158 -98231 -136114
rect -98139 -136158 -98131 -136114
rect -98039 -136158 -98031 -136114
rect -97939 -136158 -97931 -136114
rect -97839 -136158 -97831 -136114
rect -97739 -136158 -97731 -136114
rect -97639 -136158 -97631 -136114
rect -97539 -136158 -97531 -136114
rect -97439 -136158 -97431 -136114
rect -97339 -136158 -97331 -136114
rect -97239 -136158 -97231 -136114
rect -104783 -136214 -104739 -136206
rect -104683 -136214 -104639 -136206
rect -104583 -136214 -104539 -136206
rect -104483 -136214 -104439 -136206
rect -104383 -136214 -104339 -136206
rect -104283 -136214 -104239 -136206
rect -104183 -136214 -104139 -136206
rect -104083 -136214 -104039 -136206
rect -103983 -136214 -103939 -136206
rect -103883 -136214 -103839 -136206
rect -103783 -136214 -103739 -136206
rect -103683 -136214 -103639 -136206
rect -103583 -136214 -103539 -136206
rect -103483 -136214 -103439 -136206
rect -103383 -136214 -103339 -136206
rect -103283 -136214 -103239 -136206
rect -102783 -136214 -102739 -136206
rect -102683 -136214 -102639 -136206
rect -102583 -136214 -102539 -136206
rect -102483 -136214 -102439 -136206
rect -102383 -136214 -102339 -136206
rect -102283 -136214 -102239 -136206
rect -102183 -136214 -102139 -136206
rect -102083 -136214 -102039 -136206
rect -101983 -136214 -101939 -136206
rect -101883 -136214 -101839 -136206
rect -101783 -136214 -101739 -136206
rect -101683 -136214 -101639 -136206
rect -101583 -136214 -101539 -136206
rect -101483 -136214 -101439 -136206
rect -101383 -136214 -101339 -136206
rect -101283 -136214 -101239 -136206
rect -100783 -136214 -100739 -136206
rect -100683 -136214 -100639 -136206
rect -100583 -136214 -100539 -136206
rect -100483 -136214 -100439 -136206
rect -100383 -136214 -100339 -136206
rect -100283 -136214 -100239 -136206
rect -100183 -136214 -100139 -136206
rect -100083 -136214 -100039 -136206
rect -99983 -136214 -99939 -136206
rect -99883 -136214 -99839 -136206
rect -99783 -136214 -99739 -136206
rect -99683 -136214 -99639 -136206
rect -99583 -136214 -99539 -136206
rect -99483 -136214 -99439 -136206
rect -99383 -136214 -99339 -136206
rect -99283 -136214 -99239 -136206
rect -98783 -136214 -98739 -136206
rect -98683 -136214 -98639 -136206
rect -98583 -136214 -98539 -136206
rect -98483 -136214 -98439 -136206
rect -98383 -136214 -98339 -136206
rect -98283 -136214 -98239 -136206
rect -98183 -136214 -98139 -136206
rect -98083 -136214 -98039 -136206
rect -97983 -136214 -97939 -136206
rect -97883 -136214 -97839 -136206
rect -97783 -136214 -97739 -136206
rect -97683 -136214 -97639 -136206
rect -97583 -136214 -97539 -136206
rect -97483 -136214 -97439 -136206
rect -97383 -136214 -97339 -136206
rect -97283 -136214 -97239 -136206
rect -104739 -136258 -104731 -136214
rect -104639 -136258 -104631 -136214
rect -104539 -136258 -104531 -136214
rect -104439 -136258 -104431 -136214
rect -104339 -136258 -104331 -136214
rect -104239 -136258 -104231 -136214
rect -104139 -136258 -104131 -136214
rect -104039 -136258 -104031 -136214
rect -103939 -136258 -103931 -136214
rect -103839 -136258 -103831 -136214
rect -103739 -136258 -103731 -136214
rect -103639 -136258 -103631 -136214
rect -103539 -136258 -103531 -136214
rect -103439 -136258 -103431 -136214
rect -103339 -136258 -103331 -136214
rect -103239 -136258 -103231 -136214
rect -102739 -136258 -102731 -136214
rect -102639 -136258 -102631 -136214
rect -102539 -136258 -102531 -136214
rect -102439 -136258 -102431 -136214
rect -102339 -136258 -102331 -136214
rect -102239 -136258 -102231 -136214
rect -102139 -136258 -102131 -136214
rect -102039 -136258 -102031 -136214
rect -101939 -136258 -101931 -136214
rect -101839 -136258 -101831 -136214
rect -101739 -136258 -101731 -136214
rect -101639 -136258 -101631 -136214
rect -101539 -136258 -101531 -136214
rect -101439 -136258 -101431 -136214
rect -101339 -136258 -101331 -136214
rect -101239 -136258 -101231 -136214
rect -100739 -136258 -100731 -136214
rect -100639 -136258 -100631 -136214
rect -100539 -136258 -100531 -136214
rect -100439 -136258 -100431 -136214
rect -100339 -136258 -100331 -136214
rect -100239 -136258 -100231 -136214
rect -100139 -136258 -100131 -136214
rect -100039 -136258 -100031 -136214
rect -99939 -136258 -99931 -136214
rect -99839 -136258 -99831 -136214
rect -99739 -136258 -99731 -136214
rect -99639 -136258 -99631 -136214
rect -99539 -136258 -99531 -136214
rect -99439 -136258 -99431 -136214
rect -99339 -136258 -99331 -136214
rect -99239 -136258 -99231 -136214
rect -98739 -136258 -98731 -136214
rect -98639 -136258 -98631 -136214
rect -98539 -136258 -98531 -136214
rect -98439 -136258 -98431 -136214
rect -98339 -136258 -98331 -136214
rect -98239 -136258 -98231 -136214
rect -98139 -136258 -98131 -136214
rect -98039 -136258 -98031 -136214
rect -97939 -136258 -97931 -136214
rect -97839 -136258 -97831 -136214
rect -97739 -136258 -97731 -136214
rect -97639 -136258 -97631 -136214
rect -97539 -136258 -97531 -136214
rect -97439 -136258 -97431 -136214
rect -97339 -136258 -97331 -136214
rect -97239 -136258 -97231 -136214
rect -104783 -136314 -104739 -136306
rect -104683 -136314 -104639 -136306
rect -104583 -136314 -104539 -136306
rect -104483 -136314 -104439 -136306
rect -104383 -136314 -104339 -136306
rect -104283 -136314 -104239 -136306
rect -104183 -136314 -104139 -136306
rect -104083 -136314 -104039 -136306
rect -103983 -136314 -103939 -136306
rect -103883 -136314 -103839 -136306
rect -103783 -136314 -103739 -136306
rect -103683 -136314 -103639 -136306
rect -103583 -136314 -103539 -136306
rect -103483 -136314 -103439 -136306
rect -103383 -136314 -103339 -136306
rect -103283 -136314 -103239 -136306
rect -102783 -136314 -102739 -136306
rect -102683 -136314 -102639 -136306
rect -102583 -136314 -102539 -136306
rect -102483 -136314 -102439 -136306
rect -102383 -136314 -102339 -136306
rect -102283 -136314 -102239 -136306
rect -102183 -136314 -102139 -136306
rect -102083 -136314 -102039 -136306
rect -101983 -136314 -101939 -136306
rect -101883 -136314 -101839 -136306
rect -101783 -136314 -101739 -136306
rect -101683 -136314 -101639 -136306
rect -101583 -136314 -101539 -136306
rect -101483 -136314 -101439 -136306
rect -101383 -136314 -101339 -136306
rect -101283 -136314 -101239 -136306
rect -100783 -136314 -100739 -136306
rect -100683 -136314 -100639 -136306
rect -100583 -136314 -100539 -136306
rect -100483 -136314 -100439 -136306
rect -100383 -136314 -100339 -136306
rect -100283 -136314 -100239 -136306
rect -100183 -136314 -100139 -136306
rect -100083 -136314 -100039 -136306
rect -99983 -136314 -99939 -136306
rect -99883 -136314 -99839 -136306
rect -99783 -136314 -99739 -136306
rect -99683 -136314 -99639 -136306
rect -99583 -136314 -99539 -136306
rect -99483 -136314 -99439 -136306
rect -99383 -136314 -99339 -136306
rect -99283 -136314 -99239 -136306
rect -98783 -136314 -98739 -136306
rect -98683 -136314 -98639 -136306
rect -98583 -136314 -98539 -136306
rect -98483 -136314 -98439 -136306
rect -98383 -136314 -98339 -136306
rect -98283 -136314 -98239 -136306
rect -98183 -136314 -98139 -136306
rect -98083 -136314 -98039 -136306
rect -97983 -136314 -97939 -136306
rect -97883 -136314 -97839 -136306
rect -97783 -136314 -97739 -136306
rect -97683 -136314 -97639 -136306
rect -97583 -136314 -97539 -136306
rect -97483 -136314 -97439 -136306
rect -97383 -136314 -97339 -136306
rect -97283 -136314 -97239 -136306
rect -104739 -136358 -104731 -136314
rect -104639 -136358 -104631 -136314
rect -104539 -136358 -104531 -136314
rect -104439 -136358 -104431 -136314
rect -104339 -136358 -104331 -136314
rect -104239 -136358 -104231 -136314
rect -104139 -136358 -104131 -136314
rect -104039 -136358 -104031 -136314
rect -103939 -136358 -103931 -136314
rect -103839 -136358 -103831 -136314
rect -103739 -136358 -103731 -136314
rect -103639 -136358 -103631 -136314
rect -103539 -136358 -103531 -136314
rect -103439 -136358 -103431 -136314
rect -103339 -136358 -103331 -136314
rect -103239 -136358 -103231 -136314
rect -102739 -136358 -102731 -136314
rect -102639 -136358 -102631 -136314
rect -102539 -136358 -102531 -136314
rect -102439 -136358 -102431 -136314
rect -102339 -136358 -102331 -136314
rect -102239 -136358 -102231 -136314
rect -102139 -136358 -102131 -136314
rect -102039 -136358 -102031 -136314
rect -101939 -136358 -101931 -136314
rect -101839 -136358 -101831 -136314
rect -101739 -136358 -101731 -136314
rect -101639 -136358 -101631 -136314
rect -101539 -136358 -101531 -136314
rect -101439 -136358 -101431 -136314
rect -101339 -136358 -101331 -136314
rect -101239 -136358 -101231 -136314
rect -100739 -136358 -100731 -136314
rect -100639 -136358 -100631 -136314
rect -100539 -136358 -100531 -136314
rect -100439 -136358 -100431 -136314
rect -100339 -136358 -100331 -136314
rect -100239 -136358 -100231 -136314
rect -100139 -136358 -100131 -136314
rect -100039 -136358 -100031 -136314
rect -99939 -136358 -99931 -136314
rect -99839 -136358 -99831 -136314
rect -99739 -136358 -99731 -136314
rect -99639 -136358 -99631 -136314
rect -99539 -136358 -99531 -136314
rect -99439 -136358 -99431 -136314
rect -99339 -136358 -99331 -136314
rect -99239 -136358 -99231 -136314
rect -98739 -136358 -98731 -136314
rect -98639 -136358 -98631 -136314
rect -98539 -136358 -98531 -136314
rect -98439 -136358 -98431 -136314
rect -98339 -136358 -98331 -136314
rect -98239 -136358 -98231 -136314
rect -98139 -136358 -98131 -136314
rect -98039 -136358 -98031 -136314
rect -97939 -136358 -97931 -136314
rect -97839 -136358 -97831 -136314
rect -97739 -136358 -97731 -136314
rect -97639 -136358 -97631 -136314
rect -97539 -136358 -97531 -136314
rect -97439 -136358 -97431 -136314
rect -97339 -136358 -97331 -136314
rect -97239 -136358 -97231 -136314
rect -104783 -136414 -104739 -136406
rect -104683 -136414 -104639 -136406
rect -104583 -136414 -104539 -136406
rect -104483 -136414 -104439 -136406
rect -104383 -136414 -104339 -136406
rect -104283 -136414 -104239 -136406
rect -104183 -136414 -104139 -136406
rect -104083 -136414 -104039 -136406
rect -103983 -136414 -103939 -136406
rect -103883 -136414 -103839 -136406
rect -103783 -136414 -103739 -136406
rect -103683 -136414 -103639 -136406
rect -103583 -136414 -103539 -136406
rect -103483 -136414 -103439 -136406
rect -103383 -136414 -103339 -136406
rect -103283 -136414 -103239 -136406
rect -102783 -136414 -102739 -136406
rect -102683 -136414 -102639 -136406
rect -102583 -136414 -102539 -136406
rect -102483 -136414 -102439 -136406
rect -102383 -136414 -102339 -136406
rect -102283 -136414 -102239 -136406
rect -102183 -136414 -102139 -136406
rect -102083 -136414 -102039 -136406
rect -101983 -136414 -101939 -136406
rect -101883 -136414 -101839 -136406
rect -101783 -136414 -101739 -136406
rect -101683 -136414 -101639 -136406
rect -101583 -136414 -101539 -136406
rect -101483 -136414 -101439 -136406
rect -101383 -136414 -101339 -136406
rect -101283 -136414 -101239 -136406
rect -100783 -136414 -100739 -136406
rect -100683 -136414 -100639 -136406
rect -100583 -136414 -100539 -136406
rect -100483 -136414 -100439 -136406
rect -100383 -136414 -100339 -136406
rect -100283 -136414 -100239 -136406
rect -100183 -136414 -100139 -136406
rect -100083 -136414 -100039 -136406
rect -99983 -136414 -99939 -136406
rect -99883 -136414 -99839 -136406
rect -99783 -136414 -99739 -136406
rect -99683 -136414 -99639 -136406
rect -99583 -136414 -99539 -136406
rect -99483 -136414 -99439 -136406
rect -99383 -136414 -99339 -136406
rect -99283 -136414 -99239 -136406
rect -98783 -136414 -98739 -136406
rect -98683 -136414 -98639 -136406
rect -98583 -136414 -98539 -136406
rect -98483 -136414 -98439 -136406
rect -98383 -136414 -98339 -136406
rect -98283 -136414 -98239 -136406
rect -98183 -136414 -98139 -136406
rect -98083 -136414 -98039 -136406
rect -97983 -136414 -97939 -136406
rect -97883 -136414 -97839 -136406
rect -97783 -136414 -97739 -136406
rect -97683 -136414 -97639 -136406
rect -97583 -136414 -97539 -136406
rect -97483 -136414 -97439 -136406
rect -97383 -136414 -97339 -136406
rect -97283 -136414 -97239 -136406
rect -104739 -136458 -104731 -136414
rect -104639 -136458 -104631 -136414
rect -104539 -136458 -104531 -136414
rect -104439 -136458 -104431 -136414
rect -104339 -136458 -104331 -136414
rect -104239 -136458 -104231 -136414
rect -104139 -136458 -104131 -136414
rect -104039 -136458 -104031 -136414
rect -103939 -136458 -103931 -136414
rect -103839 -136458 -103831 -136414
rect -103739 -136458 -103731 -136414
rect -103639 -136458 -103631 -136414
rect -103539 -136458 -103531 -136414
rect -103439 -136458 -103431 -136414
rect -103339 -136458 -103331 -136414
rect -103239 -136458 -103231 -136414
rect -102739 -136458 -102731 -136414
rect -102639 -136458 -102631 -136414
rect -102539 -136458 -102531 -136414
rect -102439 -136458 -102431 -136414
rect -102339 -136458 -102331 -136414
rect -102239 -136458 -102231 -136414
rect -102139 -136458 -102131 -136414
rect -102039 -136458 -102031 -136414
rect -101939 -136458 -101931 -136414
rect -101839 -136458 -101831 -136414
rect -101739 -136458 -101731 -136414
rect -101639 -136458 -101631 -136414
rect -101539 -136458 -101531 -136414
rect -101439 -136458 -101431 -136414
rect -101339 -136458 -101331 -136414
rect -101239 -136458 -101231 -136414
rect -100739 -136458 -100731 -136414
rect -100639 -136458 -100631 -136414
rect -100539 -136458 -100531 -136414
rect -100439 -136458 -100431 -136414
rect -100339 -136458 -100331 -136414
rect -100239 -136458 -100231 -136414
rect -100139 -136458 -100131 -136414
rect -100039 -136458 -100031 -136414
rect -99939 -136458 -99931 -136414
rect -99839 -136458 -99831 -136414
rect -99739 -136458 -99731 -136414
rect -99639 -136458 -99631 -136414
rect -99539 -136458 -99531 -136414
rect -99439 -136458 -99431 -136414
rect -99339 -136458 -99331 -136414
rect -99239 -136458 -99231 -136414
rect -98739 -136458 -98731 -136414
rect -98639 -136458 -98631 -136414
rect -98539 -136458 -98531 -136414
rect -98439 -136458 -98431 -136414
rect -98339 -136458 -98331 -136414
rect -98239 -136458 -98231 -136414
rect -98139 -136458 -98131 -136414
rect -98039 -136458 -98031 -136414
rect -97939 -136458 -97931 -136414
rect -97839 -136458 -97831 -136414
rect -97739 -136458 -97731 -136414
rect -97639 -136458 -97631 -136414
rect -97539 -136458 -97531 -136414
rect -97439 -136458 -97431 -136414
rect -97339 -136458 -97331 -136414
rect -97239 -136458 -97231 -136414
rect -104783 -136514 -104739 -136506
rect -104683 -136514 -104639 -136506
rect -104583 -136514 -104539 -136506
rect -104483 -136514 -104439 -136506
rect -104383 -136514 -104339 -136506
rect -104283 -136514 -104239 -136506
rect -104183 -136514 -104139 -136506
rect -104083 -136514 -104039 -136506
rect -103983 -136514 -103939 -136506
rect -103883 -136514 -103839 -136506
rect -103783 -136514 -103739 -136506
rect -103683 -136514 -103639 -136506
rect -103583 -136514 -103539 -136506
rect -103483 -136514 -103439 -136506
rect -103383 -136514 -103339 -136506
rect -103283 -136514 -103239 -136506
rect -102783 -136514 -102739 -136506
rect -102683 -136514 -102639 -136506
rect -102583 -136514 -102539 -136506
rect -102483 -136514 -102439 -136506
rect -102383 -136514 -102339 -136506
rect -102283 -136514 -102239 -136506
rect -102183 -136514 -102139 -136506
rect -102083 -136514 -102039 -136506
rect -101983 -136514 -101939 -136506
rect -101883 -136514 -101839 -136506
rect -101783 -136514 -101739 -136506
rect -101683 -136514 -101639 -136506
rect -101583 -136514 -101539 -136506
rect -101483 -136514 -101439 -136506
rect -101383 -136514 -101339 -136506
rect -101283 -136514 -101239 -136506
rect -100783 -136514 -100739 -136506
rect -100683 -136514 -100639 -136506
rect -100583 -136514 -100539 -136506
rect -100483 -136514 -100439 -136506
rect -100383 -136514 -100339 -136506
rect -100283 -136514 -100239 -136506
rect -100183 -136514 -100139 -136506
rect -100083 -136514 -100039 -136506
rect -99983 -136514 -99939 -136506
rect -99883 -136514 -99839 -136506
rect -99783 -136514 -99739 -136506
rect -99683 -136514 -99639 -136506
rect -99583 -136514 -99539 -136506
rect -99483 -136514 -99439 -136506
rect -99383 -136514 -99339 -136506
rect -99283 -136514 -99239 -136506
rect -98783 -136514 -98739 -136506
rect -98683 -136514 -98639 -136506
rect -98583 -136514 -98539 -136506
rect -98483 -136514 -98439 -136506
rect -98383 -136514 -98339 -136506
rect -98283 -136514 -98239 -136506
rect -98183 -136514 -98139 -136506
rect -98083 -136514 -98039 -136506
rect -97983 -136514 -97939 -136506
rect -97883 -136514 -97839 -136506
rect -97783 -136514 -97739 -136506
rect -97683 -136514 -97639 -136506
rect -97583 -136514 -97539 -136506
rect -97483 -136514 -97439 -136506
rect -97383 -136514 -97339 -136506
rect -97283 -136514 -97239 -136506
rect -104739 -136558 -104731 -136514
rect -104639 -136558 -104631 -136514
rect -104539 -136558 -104531 -136514
rect -104439 -136558 -104431 -136514
rect -104339 -136558 -104331 -136514
rect -104239 -136558 -104231 -136514
rect -104139 -136558 -104131 -136514
rect -104039 -136558 -104031 -136514
rect -103939 -136558 -103931 -136514
rect -103839 -136558 -103831 -136514
rect -103739 -136558 -103731 -136514
rect -103639 -136558 -103631 -136514
rect -103539 -136558 -103531 -136514
rect -103439 -136558 -103431 -136514
rect -103339 -136558 -103331 -136514
rect -103239 -136558 -103231 -136514
rect -102739 -136558 -102731 -136514
rect -102639 -136558 -102631 -136514
rect -102539 -136558 -102531 -136514
rect -102439 -136558 -102431 -136514
rect -102339 -136558 -102331 -136514
rect -102239 -136558 -102231 -136514
rect -102139 -136558 -102131 -136514
rect -102039 -136558 -102031 -136514
rect -101939 -136558 -101931 -136514
rect -101839 -136558 -101831 -136514
rect -101739 -136558 -101731 -136514
rect -101639 -136558 -101631 -136514
rect -101539 -136558 -101531 -136514
rect -101439 -136558 -101431 -136514
rect -101339 -136558 -101331 -136514
rect -101239 -136558 -101231 -136514
rect -100739 -136558 -100731 -136514
rect -100639 -136558 -100631 -136514
rect -100539 -136558 -100531 -136514
rect -100439 -136558 -100431 -136514
rect -100339 -136558 -100331 -136514
rect -100239 -136558 -100231 -136514
rect -100139 -136558 -100131 -136514
rect -100039 -136558 -100031 -136514
rect -99939 -136558 -99931 -136514
rect -99839 -136558 -99831 -136514
rect -99739 -136558 -99731 -136514
rect -99639 -136558 -99631 -136514
rect -99539 -136558 -99531 -136514
rect -99439 -136558 -99431 -136514
rect -99339 -136558 -99331 -136514
rect -99239 -136558 -99231 -136514
rect -98739 -136558 -98731 -136514
rect -98639 -136558 -98631 -136514
rect -98539 -136558 -98531 -136514
rect -98439 -136558 -98431 -136514
rect -98339 -136558 -98331 -136514
rect -98239 -136558 -98231 -136514
rect -98139 -136558 -98131 -136514
rect -98039 -136558 -98031 -136514
rect -97939 -136558 -97931 -136514
rect -97839 -136558 -97831 -136514
rect -97739 -136558 -97731 -136514
rect -97639 -136558 -97631 -136514
rect -97539 -136558 -97531 -136514
rect -97439 -136558 -97431 -136514
rect -97339 -136558 -97331 -136514
rect -97239 -136558 -97231 -136514
rect -104783 -136614 -104739 -136606
rect -104683 -136614 -104639 -136606
rect -104583 -136614 -104539 -136606
rect -104483 -136614 -104439 -136606
rect -104383 -136614 -104339 -136606
rect -104283 -136614 -104239 -136606
rect -104183 -136614 -104139 -136606
rect -104083 -136614 -104039 -136606
rect -103983 -136614 -103939 -136606
rect -103883 -136614 -103839 -136606
rect -103783 -136614 -103739 -136606
rect -103683 -136614 -103639 -136606
rect -103583 -136614 -103539 -136606
rect -103483 -136614 -103439 -136606
rect -103383 -136614 -103339 -136606
rect -103283 -136614 -103239 -136606
rect -102783 -136614 -102739 -136606
rect -102683 -136614 -102639 -136606
rect -102583 -136614 -102539 -136606
rect -102483 -136614 -102439 -136606
rect -102383 -136614 -102339 -136606
rect -102283 -136614 -102239 -136606
rect -102183 -136614 -102139 -136606
rect -102083 -136614 -102039 -136606
rect -101983 -136614 -101939 -136606
rect -101883 -136614 -101839 -136606
rect -101783 -136614 -101739 -136606
rect -101683 -136614 -101639 -136606
rect -101583 -136614 -101539 -136606
rect -101483 -136614 -101439 -136606
rect -101383 -136614 -101339 -136606
rect -101283 -136614 -101239 -136606
rect -100783 -136614 -100739 -136606
rect -100683 -136614 -100639 -136606
rect -100583 -136614 -100539 -136606
rect -100483 -136614 -100439 -136606
rect -100383 -136614 -100339 -136606
rect -100283 -136614 -100239 -136606
rect -100183 -136614 -100139 -136606
rect -100083 -136614 -100039 -136606
rect -99983 -136614 -99939 -136606
rect -99883 -136614 -99839 -136606
rect -99783 -136614 -99739 -136606
rect -99683 -136614 -99639 -136606
rect -99583 -136614 -99539 -136606
rect -99483 -136614 -99439 -136606
rect -99383 -136614 -99339 -136606
rect -99283 -136614 -99239 -136606
rect -98783 -136614 -98739 -136606
rect -98683 -136614 -98639 -136606
rect -98583 -136614 -98539 -136606
rect -98483 -136614 -98439 -136606
rect -98383 -136614 -98339 -136606
rect -98283 -136614 -98239 -136606
rect -98183 -136614 -98139 -136606
rect -98083 -136614 -98039 -136606
rect -97983 -136614 -97939 -136606
rect -97883 -136614 -97839 -136606
rect -97783 -136614 -97739 -136606
rect -97683 -136614 -97639 -136606
rect -97583 -136614 -97539 -136606
rect -97483 -136614 -97439 -136606
rect -97383 -136614 -97339 -136606
rect -97283 -136614 -97239 -136606
rect -104739 -136658 -104731 -136614
rect -104639 -136658 -104631 -136614
rect -104539 -136658 -104531 -136614
rect -104439 -136658 -104431 -136614
rect -104339 -136658 -104331 -136614
rect -104239 -136658 -104231 -136614
rect -104139 -136658 -104131 -136614
rect -104039 -136658 -104031 -136614
rect -103939 -136658 -103931 -136614
rect -103839 -136658 -103831 -136614
rect -103739 -136658 -103731 -136614
rect -103639 -136658 -103631 -136614
rect -103539 -136658 -103531 -136614
rect -103439 -136658 -103431 -136614
rect -103339 -136658 -103331 -136614
rect -103239 -136658 -103231 -136614
rect -102739 -136658 -102731 -136614
rect -102639 -136658 -102631 -136614
rect -102539 -136658 -102531 -136614
rect -102439 -136658 -102431 -136614
rect -102339 -136658 -102331 -136614
rect -102239 -136658 -102231 -136614
rect -102139 -136658 -102131 -136614
rect -102039 -136658 -102031 -136614
rect -101939 -136658 -101931 -136614
rect -101839 -136658 -101831 -136614
rect -101739 -136658 -101731 -136614
rect -101639 -136658 -101631 -136614
rect -101539 -136658 -101531 -136614
rect -101439 -136658 -101431 -136614
rect -101339 -136658 -101331 -136614
rect -101239 -136658 -101231 -136614
rect -100739 -136658 -100731 -136614
rect -100639 -136658 -100631 -136614
rect -100539 -136658 -100531 -136614
rect -100439 -136658 -100431 -136614
rect -100339 -136658 -100331 -136614
rect -100239 -136658 -100231 -136614
rect -100139 -136658 -100131 -136614
rect -100039 -136658 -100031 -136614
rect -99939 -136658 -99931 -136614
rect -99839 -136658 -99831 -136614
rect -99739 -136658 -99731 -136614
rect -99639 -136658 -99631 -136614
rect -99539 -136658 -99531 -136614
rect -99439 -136658 -99431 -136614
rect -99339 -136658 -99331 -136614
rect -99239 -136658 -99231 -136614
rect -98739 -136658 -98731 -136614
rect -98639 -136658 -98631 -136614
rect -98539 -136658 -98531 -136614
rect -98439 -136658 -98431 -136614
rect -98339 -136658 -98331 -136614
rect -98239 -136658 -98231 -136614
rect -98139 -136658 -98131 -136614
rect -98039 -136658 -98031 -136614
rect -97939 -136658 -97931 -136614
rect -97839 -136658 -97831 -136614
rect -97739 -136658 -97731 -136614
rect -97639 -136658 -97631 -136614
rect -97539 -136658 -97531 -136614
rect -97439 -136658 -97431 -136614
rect -97339 -136658 -97331 -136614
rect -97239 -136658 -97231 -136614
rect -104783 -136714 -104739 -136706
rect -104683 -136714 -104639 -136706
rect -104583 -136714 -104539 -136706
rect -104483 -136714 -104439 -136706
rect -104383 -136714 -104339 -136706
rect -104283 -136714 -104239 -136706
rect -104183 -136714 -104139 -136706
rect -104083 -136714 -104039 -136706
rect -103983 -136714 -103939 -136706
rect -103883 -136714 -103839 -136706
rect -103783 -136714 -103739 -136706
rect -103683 -136714 -103639 -136706
rect -103583 -136714 -103539 -136706
rect -103483 -136714 -103439 -136706
rect -103383 -136714 -103339 -136706
rect -103283 -136714 -103239 -136706
rect -102783 -136714 -102739 -136706
rect -102683 -136714 -102639 -136706
rect -102583 -136714 -102539 -136706
rect -102483 -136714 -102439 -136706
rect -102383 -136714 -102339 -136706
rect -102283 -136714 -102239 -136706
rect -102183 -136714 -102139 -136706
rect -102083 -136714 -102039 -136706
rect -101983 -136714 -101939 -136706
rect -101883 -136714 -101839 -136706
rect -101783 -136714 -101739 -136706
rect -101683 -136714 -101639 -136706
rect -101583 -136714 -101539 -136706
rect -101483 -136714 -101439 -136706
rect -101383 -136714 -101339 -136706
rect -101283 -136714 -101239 -136706
rect -100783 -136714 -100739 -136706
rect -100683 -136714 -100639 -136706
rect -100583 -136714 -100539 -136706
rect -100483 -136714 -100439 -136706
rect -100383 -136714 -100339 -136706
rect -100283 -136714 -100239 -136706
rect -100183 -136714 -100139 -136706
rect -100083 -136714 -100039 -136706
rect -99983 -136714 -99939 -136706
rect -99883 -136714 -99839 -136706
rect -99783 -136714 -99739 -136706
rect -99683 -136714 -99639 -136706
rect -99583 -136714 -99539 -136706
rect -99483 -136714 -99439 -136706
rect -99383 -136714 -99339 -136706
rect -99283 -136714 -99239 -136706
rect -98783 -136714 -98739 -136706
rect -98683 -136714 -98639 -136706
rect -98583 -136714 -98539 -136706
rect -98483 -136714 -98439 -136706
rect -98383 -136714 -98339 -136706
rect -98283 -136714 -98239 -136706
rect -98183 -136714 -98139 -136706
rect -98083 -136714 -98039 -136706
rect -97983 -136714 -97939 -136706
rect -97883 -136714 -97839 -136706
rect -97783 -136714 -97739 -136706
rect -97683 -136714 -97639 -136706
rect -97583 -136714 -97539 -136706
rect -97483 -136714 -97439 -136706
rect -97383 -136714 -97339 -136706
rect -97283 -136714 -97239 -136706
rect -104739 -136758 -104731 -136714
rect -104639 -136758 -104631 -136714
rect -104539 -136758 -104531 -136714
rect -104439 -136758 -104431 -136714
rect -104339 -136758 -104331 -136714
rect -104239 -136758 -104231 -136714
rect -104139 -136758 -104131 -136714
rect -104039 -136758 -104031 -136714
rect -103939 -136758 -103931 -136714
rect -103839 -136758 -103831 -136714
rect -103739 -136758 -103731 -136714
rect -103639 -136758 -103631 -136714
rect -103539 -136758 -103531 -136714
rect -103439 -136758 -103431 -136714
rect -103339 -136758 -103331 -136714
rect -103239 -136758 -103231 -136714
rect -102739 -136758 -102731 -136714
rect -102639 -136758 -102631 -136714
rect -102539 -136758 -102531 -136714
rect -102439 -136758 -102431 -136714
rect -102339 -136758 -102331 -136714
rect -102239 -136758 -102231 -136714
rect -102139 -136758 -102131 -136714
rect -102039 -136758 -102031 -136714
rect -101939 -136758 -101931 -136714
rect -101839 -136758 -101831 -136714
rect -101739 -136758 -101731 -136714
rect -101639 -136758 -101631 -136714
rect -101539 -136758 -101531 -136714
rect -101439 -136758 -101431 -136714
rect -101339 -136758 -101331 -136714
rect -101239 -136758 -101231 -136714
rect -100739 -136758 -100731 -136714
rect -100639 -136758 -100631 -136714
rect -100539 -136758 -100531 -136714
rect -100439 -136758 -100431 -136714
rect -100339 -136758 -100331 -136714
rect -100239 -136758 -100231 -136714
rect -100139 -136758 -100131 -136714
rect -100039 -136758 -100031 -136714
rect -99939 -136758 -99931 -136714
rect -99839 -136758 -99831 -136714
rect -99739 -136758 -99731 -136714
rect -99639 -136758 -99631 -136714
rect -99539 -136758 -99531 -136714
rect -99439 -136758 -99431 -136714
rect -99339 -136758 -99331 -136714
rect -99239 -136758 -99231 -136714
rect -98739 -136758 -98731 -136714
rect -98639 -136758 -98631 -136714
rect -98539 -136758 -98531 -136714
rect -98439 -136758 -98431 -136714
rect -98339 -136758 -98331 -136714
rect -98239 -136758 -98231 -136714
rect -98139 -136758 -98131 -136714
rect -98039 -136758 -98031 -136714
rect -97939 -136758 -97931 -136714
rect -97839 -136758 -97831 -136714
rect -97739 -136758 -97731 -136714
rect -97639 -136758 -97631 -136714
rect -97539 -136758 -97531 -136714
rect -97439 -136758 -97431 -136714
rect -97339 -136758 -97331 -136714
rect -97239 -136758 -97231 -136714
rect -104783 -136814 -104739 -136806
rect -104683 -136814 -104639 -136806
rect -104583 -136814 -104539 -136806
rect -104483 -136814 -104439 -136806
rect -104383 -136814 -104339 -136806
rect -104283 -136814 -104239 -136806
rect -104183 -136814 -104139 -136806
rect -104083 -136814 -104039 -136806
rect -103983 -136814 -103939 -136806
rect -103883 -136814 -103839 -136806
rect -103783 -136814 -103739 -136806
rect -103683 -136814 -103639 -136806
rect -103583 -136814 -103539 -136806
rect -103483 -136814 -103439 -136806
rect -103383 -136814 -103339 -136806
rect -103283 -136814 -103239 -136806
rect -102783 -136814 -102739 -136806
rect -102683 -136814 -102639 -136806
rect -102583 -136814 -102539 -136806
rect -102483 -136814 -102439 -136806
rect -102383 -136814 -102339 -136806
rect -102283 -136814 -102239 -136806
rect -102183 -136814 -102139 -136806
rect -102083 -136814 -102039 -136806
rect -101983 -136814 -101939 -136806
rect -101883 -136814 -101839 -136806
rect -101783 -136814 -101739 -136806
rect -101683 -136814 -101639 -136806
rect -101583 -136814 -101539 -136806
rect -101483 -136814 -101439 -136806
rect -101383 -136814 -101339 -136806
rect -101283 -136814 -101239 -136806
rect -100783 -136814 -100739 -136806
rect -100683 -136814 -100639 -136806
rect -100583 -136814 -100539 -136806
rect -100483 -136814 -100439 -136806
rect -100383 -136814 -100339 -136806
rect -100283 -136814 -100239 -136806
rect -100183 -136814 -100139 -136806
rect -100083 -136814 -100039 -136806
rect -99983 -136814 -99939 -136806
rect -99883 -136814 -99839 -136806
rect -99783 -136814 -99739 -136806
rect -99683 -136814 -99639 -136806
rect -99583 -136814 -99539 -136806
rect -99483 -136814 -99439 -136806
rect -99383 -136814 -99339 -136806
rect -99283 -136814 -99239 -136806
rect -98783 -136814 -98739 -136806
rect -98683 -136814 -98639 -136806
rect -98583 -136814 -98539 -136806
rect -98483 -136814 -98439 -136806
rect -98383 -136814 -98339 -136806
rect -98283 -136814 -98239 -136806
rect -98183 -136814 -98139 -136806
rect -98083 -136814 -98039 -136806
rect -97983 -136814 -97939 -136806
rect -97883 -136814 -97839 -136806
rect -97783 -136814 -97739 -136806
rect -97683 -136814 -97639 -136806
rect -97583 -136814 -97539 -136806
rect -97483 -136814 -97439 -136806
rect -97383 -136814 -97339 -136806
rect -97283 -136814 -97239 -136806
rect -104739 -136858 -104731 -136814
rect -104639 -136858 -104631 -136814
rect -104539 -136858 -104531 -136814
rect -104439 -136858 -104431 -136814
rect -104339 -136858 -104331 -136814
rect -104239 -136858 -104231 -136814
rect -104139 -136858 -104131 -136814
rect -104039 -136858 -104031 -136814
rect -103939 -136858 -103931 -136814
rect -103839 -136858 -103831 -136814
rect -103739 -136858 -103731 -136814
rect -103639 -136858 -103631 -136814
rect -103539 -136858 -103531 -136814
rect -103439 -136858 -103431 -136814
rect -103339 -136858 -103331 -136814
rect -103239 -136858 -103231 -136814
rect -102739 -136858 -102731 -136814
rect -102639 -136858 -102631 -136814
rect -102539 -136858 -102531 -136814
rect -102439 -136858 -102431 -136814
rect -102339 -136858 -102331 -136814
rect -102239 -136858 -102231 -136814
rect -102139 -136858 -102131 -136814
rect -102039 -136858 -102031 -136814
rect -101939 -136858 -101931 -136814
rect -101839 -136858 -101831 -136814
rect -101739 -136858 -101731 -136814
rect -101639 -136858 -101631 -136814
rect -101539 -136858 -101531 -136814
rect -101439 -136858 -101431 -136814
rect -101339 -136858 -101331 -136814
rect -101239 -136858 -101231 -136814
rect -100739 -136858 -100731 -136814
rect -100639 -136858 -100631 -136814
rect -100539 -136858 -100531 -136814
rect -100439 -136858 -100431 -136814
rect -100339 -136858 -100331 -136814
rect -100239 -136858 -100231 -136814
rect -100139 -136858 -100131 -136814
rect -100039 -136858 -100031 -136814
rect -99939 -136858 -99931 -136814
rect -99839 -136858 -99831 -136814
rect -99739 -136858 -99731 -136814
rect -99639 -136858 -99631 -136814
rect -99539 -136858 -99531 -136814
rect -99439 -136858 -99431 -136814
rect -99339 -136858 -99331 -136814
rect -99239 -136858 -99231 -136814
rect -98739 -136858 -98731 -136814
rect -98639 -136858 -98631 -136814
rect -98539 -136858 -98531 -136814
rect -98439 -136858 -98431 -136814
rect -98339 -136858 -98331 -136814
rect -98239 -136858 -98231 -136814
rect -98139 -136858 -98131 -136814
rect -98039 -136858 -98031 -136814
rect -97939 -136858 -97931 -136814
rect -97839 -136858 -97831 -136814
rect -97739 -136858 -97731 -136814
rect -97639 -136858 -97631 -136814
rect -97539 -136858 -97531 -136814
rect -97439 -136858 -97431 -136814
rect -97339 -136858 -97331 -136814
rect -97239 -136858 -97231 -136814
rect 81632 -137966 81676 -137958
rect 81732 -137966 81776 -137958
rect 81832 -137966 81876 -137958
rect 81932 -137966 81976 -137958
rect 82032 -137966 82076 -137958
rect 82132 -137966 82176 -137958
rect 82232 -137966 82276 -137958
rect 82332 -137966 82376 -137958
rect 82432 -137966 82476 -137958
rect 82532 -137966 82576 -137958
rect 82632 -137966 82676 -137958
rect 82732 -137966 82776 -137958
rect 82832 -137966 82876 -137958
rect 82932 -137966 82976 -137958
rect 83032 -137966 83076 -137958
rect 83132 -137966 83176 -137958
rect 83632 -137966 83676 -137958
rect 83732 -137966 83776 -137958
rect 83832 -137966 83876 -137958
rect 83932 -137966 83976 -137958
rect 84032 -137966 84076 -137958
rect 84132 -137966 84176 -137958
rect 84232 -137966 84276 -137958
rect 84332 -137966 84376 -137958
rect 84432 -137966 84476 -137958
rect 84532 -137966 84576 -137958
rect 84632 -137966 84676 -137958
rect 84732 -137966 84776 -137958
rect 84832 -137966 84876 -137958
rect 84932 -137966 84976 -137958
rect 85032 -137966 85076 -137958
rect 85132 -137966 85176 -137958
rect 85632 -137966 85676 -137958
rect 85732 -137966 85776 -137958
rect 85832 -137966 85876 -137958
rect 85932 -137966 85976 -137958
rect 86032 -137966 86076 -137958
rect 86132 -137966 86176 -137958
rect 86232 -137966 86276 -137958
rect 86332 -137966 86376 -137958
rect 86432 -137966 86476 -137958
rect 86532 -137966 86576 -137958
rect 86632 -137966 86676 -137958
rect 86732 -137966 86776 -137958
rect 86832 -137966 86876 -137958
rect 86932 -137966 86976 -137958
rect 87032 -137966 87076 -137958
rect 87132 -137966 87176 -137958
rect 87632 -137966 87676 -137958
rect 87732 -137966 87776 -137958
rect 87832 -137966 87876 -137958
rect 87932 -137966 87976 -137958
rect 88032 -137966 88076 -137958
rect 88132 -137966 88176 -137958
rect 88232 -137966 88276 -137958
rect 88332 -137966 88376 -137958
rect 88432 -137966 88476 -137958
rect 88532 -137966 88576 -137958
rect 88632 -137966 88676 -137958
rect 88732 -137966 88776 -137958
rect 88832 -137966 88876 -137958
rect 88932 -137966 88976 -137958
rect 89032 -137966 89076 -137958
rect 89132 -137966 89176 -137958
rect 81676 -138010 81684 -137966
rect 81776 -138010 81784 -137966
rect 81876 -138010 81884 -137966
rect 81976 -138010 81984 -137966
rect 82076 -138010 82084 -137966
rect 82176 -138010 82184 -137966
rect 82276 -138010 82284 -137966
rect 82376 -138010 82384 -137966
rect 82476 -138010 82484 -137966
rect 82576 -138010 82584 -137966
rect 82676 -138010 82684 -137966
rect 82776 -138010 82784 -137966
rect 82876 -138010 82884 -137966
rect 82976 -138010 82984 -137966
rect 83076 -138010 83084 -137966
rect 83176 -138010 83184 -137966
rect 83676 -138010 83684 -137966
rect 83776 -138010 83784 -137966
rect 83876 -138010 83884 -137966
rect 83976 -138010 83984 -137966
rect 84076 -138010 84084 -137966
rect 84176 -138010 84184 -137966
rect 84276 -138010 84284 -137966
rect 84376 -138010 84384 -137966
rect 84476 -138010 84484 -137966
rect 84576 -138010 84584 -137966
rect 84676 -138010 84684 -137966
rect 84776 -138010 84784 -137966
rect 84876 -138010 84884 -137966
rect 84976 -138010 84984 -137966
rect 85076 -138010 85084 -137966
rect 85176 -138010 85184 -137966
rect 85676 -138010 85684 -137966
rect 85776 -138010 85784 -137966
rect 85876 -138010 85884 -137966
rect 85976 -138010 85984 -137966
rect 86076 -138010 86084 -137966
rect 86176 -138010 86184 -137966
rect 86276 -138010 86284 -137966
rect 86376 -138010 86384 -137966
rect 86476 -138010 86484 -137966
rect 86576 -138010 86584 -137966
rect 86676 -138010 86684 -137966
rect 86776 -138010 86784 -137966
rect 86876 -138010 86884 -137966
rect 86976 -138010 86984 -137966
rect 87076 -138010 87084 -137966
rect 87176 -138010 87184 -137966
rect 87676 -138010 87684 -137966
rect 87776 -138010 87784 -137966
rect 87876 -138010 87884 -137966
rect 87976 -138010 87984 -137966
rect 88076 -138010 88084 -137966
rect 88176 -138010 88184 -137966
rect 88276 -138010 88284 -137966
rect 88376 -138010 88384 -137966
rect 88476 -138010 88484 -137966
rect 88576 -138010 88584 -137966
rect 88676 -138010 88684 -137966
rect 88776 -138010 88784 -137966
rect 88876 -138010 88884 -137966
rect 88976 -138010 88984 -137966
rect 89076 -138010 89084 -137966
rect 89176 -138010 89184 -137966
rect 81632 -138066 81676 -138058
rect 81732 -138066 81776 -138058
rect 81832 -138066 81876 -138058
rect 81932 -138066 81976 -138058
rect 82032 -138066 82076 -138058
rect 82132 -138066 82176 -138058
rect 82232 -138066 82276 -138058
rect 82332 -138066 82376 -138058
rect 82432 -138066 82476 -138058
rect 82532 -138066 82576 -138058
rect 82632 -138066 82676 -138058
rect 82732 -138066 82776 -138058
rect 82832 -138066 82876 -138058
rect 82932 -138066 82976 -138058
rect 83032 -138066 83076 -138058
rect 83132 -138066 83176 -138058
rect 83632 -138066 83676 -138058
rect 83732 -138066 83776 -138058
rect 83832 -138066 83876 -138058
rect 83932 -138066 83976 -138058
rect 84032 -138066 84076 -138058
rect 84132 -138066 84176 -138058
rect 84232 -138066 84276 -138058
rect 84332 -138066 84376 -138058
rect 84432 -138066 84476 -138058
rect 84532 -138066 84576 -138058
rect 84632 -138066 84676 -138058
rect 84732 -138066 84776 -138058
rect 84832 -138066 84876 -138058
rect 84932 -138066 84976 -138058
rect 85032 -138066 85076 -138058
rect 85132 -138066 85176 -138058
rect 85632 -138066 85676 -138058
rect 85732 -138066 85776 -138058
rect 85832 -138066 85876 -138058
rect 85932 -138066 85976 -138058
rect 86032 -138066 86076 -138058
rect 86132 -138066 86176 -138058
rect 86232 -138066 86276 -138058
rect 86332 -138066 86376 -138058
rect 86432 -138066 86476 -138058
rect 86532 -138066 86576 -138058
rect 86632 -138066 86676 -138058
rect 86732 -138066 86776 -138058
rect 86832 -138066 86876 -138058
rect 86932 -138066 86976 -138058
rect 87032 -138066 87076 -138058
rect 87132 -138066 87176 -138058
rect 87632 -138066 87676 -138058
rect 87732 -138066 87776 -138058
rect 87832 -138066 87876 -138058
rect 87932 -138066 87976 -138058
rect 88032 -138066 88076 -138058
rect 88132 -138066 88176 -138058
rect 88232 -138066 88276 -138058
rect 88332 -138066 88376 -138058
rect 88432 -138066 88476 -138058
rect 88532 -138066 88576 -138058
rect 88632 -138066 88676 -138058
rect 88732 -138066 88776 -138058
rect 88832 -138066 88876 -138058
rect 88932 -138066 88976 -138058
rect 89032 -138066 89076 -138058
rect 89132 -138066 89176 -138058
rect 81676 -138110 81684 -138066
rect 81776 -138110 81784 -138066
rect 81876 -138110 81884 -138066
rect 81976 -138110 81984 -138066
rect 82076 -138110 82084 -138066
rect 82176 -138110 82184 -138066
rect 82276 -138110 82284 -138066
rect 82376 -138110 82384 -138066
rect 82476 -138110 82484 -138066
rect 82576 -138110 82584 -138066
rect 82676 -138110 82684 -138066
rect 82776 -138110 82784 -138066
rect 82876 -138110 82884 -138066
rect 82976 -138110 82984 -138066
rect 83076 -138110 83084 -138066
rect 83176 -138110 83184 -138066
rect 83676 -138110 83684 -138066
rect 83776 -138110 83784 -138066
rect 83876 -138110 83884 -138066
rect 83976 -138110 83984 -138066
rect 84076 -138110 84084 -138066
rect 84176 -138110 84184 -138066
rect 84276 -138110 84284 -138066
rect 84376 -138110 84384 -138066
rect 84476 -138110 84484 -138066
rect 84576 -138110 84584 -138066
rect 84676 -138110 84684 -138066
rect 84776 -138110 84784 -138066
rect 84876 -138110 84884 -138066
rect 84976 -138110 84984 -138066
rect 85076 -138110 85084 -138066
rect 85176 -138110 85184 -138066
rect 85676 -138110 85684 -138066
rect 85776 -138110 85784 -138066
rect 85876 -138110 85884 -138066
rect 85976 -138110 85984 -138066
rect 86076 -138110 86084 -138066
rect 86176 -138110 86184 -138066
rect 86276 -138110 86284 -138066
rect 86376 -138110 86384 -138066
rect 86476 -138110 86484 -138066
rect 86576 -138110 86584 -138066
rect 86676 -138110 86684 -138066
rect 86776 -138110 86784 -138066
rect 86876 -138110 86884 -138066
rect 86976 -138110 86984 -138066
rect 87076 -138110 87084 -138066
rect 87176 -138110 87184 -138066
rect 87676 -138110 87684 -138066
rect 87776 -138110 87784 -138066
rect 87876 -138110 87884 -138066
rect 87976 -138110 87984 -138066
rect 88076 -138110 88084 -138066
rect 88176 -138110 88184 -138066
rect 88276 -138110 88284 -138066
rect 88376 -138110 88384 -138066
rect 88476 -138110 88484 -138066
rect 88576 -138110 88584 -138066
rect 88676 -138110 88684 -138066
rect 88776 -138110 88784 -138066
rect 88876 -138110 88884 -138066
rect 88976 -138110 88984 -138066
rect 89076 -138110 89084 -138066
rect 89176 -138110 89184 -138066
rect 81632 -138166 81676 -138158
rect 81732 -138166 81776 -138158
rect 81832 -138166 81876 -138158
rect 81932 -138166 81976 -138158
rect 82032 -138166 82076 -138158
rect 82132 -138166 82176 -138158
rect 82232 -138166 82276 -138158
rect 82332 -138166 82376 -138158
rect 82432 -138166 82476 -138158
rect 82532 -138166 82576 -138158
rect 82632 -138166 82676 -138158
rect 82732 -138166 82776 -138158
rect 82832 -138166 82876 -138158
rect 82932 -138166 82976 -138158
rect 83032 -138166 83076 -138158
rect 83132 -138166 83176 -138158
rect 83632 -138166 83676 -138158
rect 83732 -138166 83776 -138158
rect 83832 -138166 83876 -138158
rect 83932 -138166 83976 -138158
rect 84032 -138166 84076 -138158
rect 84132 -138166 84176 -138158
rect 84232 -138166 84276 -138158
rect 84332 -138166 84376 -138158
rect 84432 -138166 84476 -138158
rect 84532 -138166 84576 -138158
rect 84632 -138166 84676 -138158
rect 84732 -138166 84776 -138158
rect 84832 -138166 84876 -138158
rect 84932 -138166 84976 -138158
rect 85032 -138166 85076 -138158
rect 85132 -138166 85176 -138158
rect 85632 -138166 85676 -138158
rect 85732 -138166 85776 -138158
rect 85832 -138166 85876 -138158
rect 85932 -138166 85976 -138158
rect 86032 -138166 86076 -138158
rect 86132 -138166 86176 -138158
rect 86232 -138166 86276 -138158
rect 86332 -138166 86376 -138158
rect 86432 -138166 86476 -138158
rect 86532 -138166 86576 -138158
rect 86632 -138166 86676 -138158
rect 86732 -138166 86776 -138158
rect 86832 -138166 86876 -138158
rect 86932 -138166 86976 -138158
rect 87032 -138166 87076 -138158
rect 87132 -138166 87176 -138158
rect 87632 -138166 87676 -138158
rect 87732 -138166 87776 -138158
rect 87832 -138166 87876 -138158
rect 87932 -138166 87976 -138158
rect 88032 -138166 88076 -138158
rect 88132 -138166 88176 -138158
rect 88232 -138166 88276 -138158
rect 88332 -138166 88376 -138158
rect 88432 -138166 88476 -138158
rect 88532 -138166 88576 -138158
rect 88632 -138166 88676 -138158
rect 88732 -138166 88776 -138158
rect 88832 -138166 88876 -138158
rect 88932 -138166 88976 -138158
rect 89032 -138166 89076 -138158
rect 89132 -138166 89176 -138158
rect 81676 -138210 81684 -138166
rect 81776 -138210 81784 -138166
rect 81876 -138210 81884 -138166
rect 81976 -138210 81984 -138166
rect 82076 -138210 82084 -138166
rect 82176 -138210 82184 -138166
rect 82276 -138210 82284 -138166
rect 82376 -138210 82384 -138166
rect 82476 -138210 82484 -138166
rect 82576 -138210 82584 -138166
rect 82676 -138210 82684 -138166
rect 82776 -138210 82784 -138166
rect 82876 -138210 82884 -138166
rect 82976 -138210 82984 -138166
rect 83076 -138210 83084 -138166
rect 83176 -138210 83184 -138166
rect 83676 -138210 83684 -138166
rect 83776 -138210 83784 -138166
rect 83876 -138210 83884 -138166
rect 83976 -138210 83984 -138166
rect 84076 -138210 84084 -138166
rect 84176 -138210 84184 -138166
rect 84276 -138210 84284 -138166
rect 84376 -138210 84384 -138166
rect 84476 -138210 84484 -138166
rect 84576 -138210 84584 -138166
rect 84676 -138210 84684 -138166
rect 84776 -138210 84784 -138166
rect 84876 -138210 84884 -138166
rect 84976 -138210 84984 -138166
rect 85076 -138210 85084 -138166
rect 85176 -138210 85184 -138166
rect 85676 -138210 85684 -138166
rect 85776 -138210 85784 -138166
rect 85876 -138210 85884 -138166
rect 85976 -138210 85984 -138166
rect 86076 -138210 86084 -138166
rect 86176 -138210 86184 -138166
rect 86276 -138210 86284 -138166
rect 86376 -138210 86384 -138166
rect 86476 -138210 86484 -138166
rect 86576 -138210 86584 -138166
rect 86676 -138210 86684 -138166
rect 86776 -138210 86784 -138166
rect 86876 -138210 86884 -138166
rect 86976 -138210 86984 -138166
rect 87076 -138210 87084 -138166
rect 87176 -138210 87184 -138166
rect 87676 -138210 87684 -138166
rect 87776 -138210 87784 -138166
rect 87876 -138210 87884 -138166
rect 87976 -138210 87984 -138166
rect 88076 -138210 88084 -138166
rect 88176 -138210 88184 -138166
rect 88276 -138210 88284 -138166
rect 88376 -138210 88384 -138166
rect 88476 -138210 88484 -138166
rect 88576 -138210 88584 -138166
rect 88676 -138210 88684 -138166
rect 88776 -138210 88784 -138166
rect 88876 -138210 88884 -138166
rect 88976 -138210 88984 -138166
rect 89076 -138210 89084 -138166
rect 89176 -138210 89184 -138166
rect 81632 -138266 81676 -138258
rect 81732 -138266 81776 -138258
rect 81832 -138266 81876 -138258
rect 81932 -138266 81976 -138258
rect 82032 -138266 82076 -138258
rect 82132 -138266 82176 -138258
rect 82232 -138266 82276 -138258
rect 82332 -138266 82376 -138258
rect 82432 -138266 82476 -138258
rect 82532 -138266 82576 -138258
rect 82632 -138266 82676 -138258
rect 82732 -138266 82776 -138258
rect 82832 -138266 82876 -138258
rect 82932 -138266 82976 -138258
rect 83032 -138266 83076 -138258
rect 83132 -138266 83176 -138258
rect 83632 -138266 83676 -138258
rect 83732 -138266 83776 -138258
rect 83832 -138266 83876 -138258
rect 83932 -138266 83976 -138258
rect 84032 -138266 84076 -138258
rect 84132 -138266 84176 -138258
rect 84232 -138266 84276 -138258
rect 84332 -138266 84376 -138258
rect 84432 -138266 84476 -138258
rect 84532 -138266 84576 -138258
rect 84632 -138266 84676 -138258
rect 84732 -138266 84776 -138258
rect 84832 -138266 84876 -138258
rect 84932 -138266 84976 -138258
rect 85032 -138266 85076 -138258
rect 85132 -138266 85176 -138258
rect 85632 -138266 85676 -138258
rect 85732 -138266 85776 -138258
rect 85832 -138266 85876 -138258
rect 85932 -138266 85976 -138258
rect 86032 -138266 86076 -138258
rect 86132 -138266 86176 -138258
rect 86232 -138266 86276 -138258
rect 86332 -138266 86376 -138258
rect 86432 -138266 86476 -138258
rect 86532 -138266 86576 -138258
rect 86632 -138266 86676 -138258
rect 86732 -138266 86776 -138258
rect 86832 -138266 86876 -138258
rect 86932 -138266 86976 -138258
rect 87032 -138266 87076 -138258
rect 87132 -138266 87176 -138258
rect 87632 -138266 87676 -138258
rect 87732 -138266 87776 -138258
rect 87832 -138266 87876 -138258
rect 87932 -138266 87976 -138258
rect 88032 -138266 88076 -138258
rect 88132 -138266 88176 -138258
rect 88232 -138266 88276 -138258
rect 88332 -138266 88376 -138258
rect 88432 -138266 88476 -138258
rect 88532 -138266 88576 -138258
rect 88632 -138266 88676 -138258
rect 88732 -138266 88776 -138258
rect 88832 -138266 88876 -138258
rect 88932 -138266 88976 -138258
rect 89032 -138266 89076 -138258
rect 89132 -138266 89176 -138258
rect 81676 -138310 81684 -138266
rect 81776 -138310 81784 -138266
rect 81876 -138310 81884 -138266
rect 81976 -138310 81984 -138266
rect 82076 -138310 82084 -138266
rect 82176 -138310 82184 -138266
rect 82276 -138310 82284 -138266
rect 82376 -138310 82384 -138266
rect 82476 -138310 82484 -138266
rect 82576 -138310 82584 -138266
rect 82676 -138310 82684 -138266
rect 82776 -138310 82784 -138266
rect 82876 -138310 82884 -138266
rect 82976 -138310 82984 -138266
rect 83076 -138310 83084 -138266
rect 83176 -138310 83184 -138266
rect 83676 -138310 83684 -138266
rect 83776 -138310 83784 -138266
rect 83876 -138310 83884 -138266
rect 83976 -138310 83984 -138266
rect 84076 -138310 84084 -138266
rect 84176 -138310 84184 -138266
rect 84276 -138310 84284 -138266
rect 84376 -138310 84384 -138266
rect 84476 -138310 84484 -138266
rect 84576 -138310 84584 -138266
rect 84676 -138310 84684 -138266
rect 84776 -138310 84784 -138266
rect 84876 -138310 84884 -138266
rect 84976 -138310 84984 -138266
rect 85076 -138310 85084 -138266
rect 85176 -138310 85184 -138266
rect 85676 -138310 85684 -138266
rect 85776 -138310 85784 -138266
rect 85876 -138310 85884 -138266
rect 85976 -138310 85984 -138266
rect 86076 -138310 86084 -138266
rect 86176 -138310 86184 -138266
rect 86276 -138310 86284 -138266
rect 86376 -138310 86384 -138266
rect 86476 -138310 86484 -138266
rect 86576 -138310 86584 -138266
rect 86676 -138310 86684 -138266
rect 86776 -138310 86784 -138266
rect 86876 -138310 86884 -138266
rect 86976 -138310 86984 -138266
rect 87076 -138310 87084 -138266
rect 87176 -138310 87184 -138266
rect 87676 -138310 87684 -138266
rect 87776 -138310 87784 -138266
rect 87876 -138310 87884 -138266
rect 87976 -138310 87984 -138266
rect 88076 -138310 88084 -138266
rect 88176 -138310 88184 -138266
rect 88276 -138310 88284 -138266
rect 88376 -138310 88384 -138266
rect 88476 -138310 88484 -138266
rect 88576 -138310 88584 -138266
rect 88676 -138310 88684 -138266
rect 88776 -138310 88784 -138266
rect 88876 -138310 88884 -138266
rect 88976 -138310 88984 -138266
rect 89076 -138310 89084 -138266
rect 89176 -138310 89184 -138266
rect 81632 -138366 81676 -138358
rect 81732 -138366 81776 -138358
rect 81832 -138366 81876 -138358
rect 81932 -138366 81976 -138358
rect 82032 -138366 82076 -138358
rect 82132 -138366 82176 -138358
rect 82232 -138366 82276 -138358
rect 82332 -138366 82376 -138358
rect 82432 -138366 82476 -138358
rect 82532 -138366 82576 -138358
rect 82632 -138366 82676 -138358
rect 82732 -138366 82776 -138358
rect 82832 -138366 82876 -138358
rect 82932 -138366 82976 -138358
rect 83032 -138366 83076 -138358
rect 83132 -138366 83176 -138358
rect 83632 -138366 83676 -138358
rect 83732 -138366 83776 -138358
rect 83832 -138366 83876 -138358
rect 83932 -138366 83976 -138358
rect 84032 -138366 84076 -138358
rect 84132 -138366 84176 -138358
rect 84232 -138366 84276 -138358
rect 84332 -138366 84376 -138358
rect 84432 -138366 84476 -138358
rect 84532 -138366 84576 -138358
rect 84632 -138366 84676 -138358
rect 84732 -138366 84776 -138358
rect 84832 -138366 84876 -138358
rect 84932 -138366 84976 -138358
rect 85032 -138366 85076 -138358
rect 85132 -138366 85176 -138358
rect 85632 -138366 85676 -138358
rect 85732 -138366 85776 -138358
rect 85832 -138366 85876 -138358
rect 85932 -138366 85976 -138358
rect 86032 -138366 86076 -138358
rect 86132 -138366 86176 -138358
rect 86232 -138366 86276 -138358
rect 86332 -138366 86376 -138358
rect 86432 -138366 86476 -138358
rect 86532 -138366 86576 -138358
rect 86632 -138366 86676 -138358
rect 86732 -138366 86776 -138358
rect 86832 -138366 86876 -138358
rect 86932 -138366 86976 -138358
rect 87032 -138366 87076 -138358
rect 87132 -138366 87176 -138358
rect 87632 -138366 87676 -138358
rect 87732 -138366 87776 -138358
rect 87832 -138366 87876 -138358
rect 87932 -138366 87976 -138358
rect 88032 -138366 88076 -138358
rect 88132 -138366 88176 -138358
rect 88232 -138366 88276 -138358
rect 88332 -138366 88376 -138358
rect 88432 -138366 88476 -138358
rect 88532 -138366 88576 -138358
rect 88632 -138366 88676 -138358
rect 88732 -138366 88776 -138358
rect 88832 -138366 88876 -138358
rect 88932 -138366 88976 -138358
rect 89032 -138366 89076 -138358
rect 89132 -138366 89176 -138358
rect 81676 -138410 81684 -138366
rect 81776 -138410 81784 -138366
rect 81876 -138410 81884 -138366
rect 81976 -138410 81984 -138366
rect 82076 -138410 82084 -138366
rect 82176 -138410 82184 -138366
rect 82276 -138410 82284 -138366
rect 82376 -138410 82384 -138366
rect 82476 -138410 82484 -138366
rect 82576 -138410 82584 -138366
rect 82676 -138410 82684 -138366
rect 82776 -138410 82784 -138366
rect 82876 -138410 82884 -138366
rect 82976 -138410 82984 -138366
rect 83076 -138410 83084 -138366
rect 83176 -138410 83184 -138366
rect 83676 -138410 83684 -138366
rect 83776 -138410 83784 -138366
rect 83876 -138410 83884 -138366
rect 83976 -138410 83984 -138366
rect 84076 -138410 84084 -138366
rect 84176 -138410 84184 -138366
rect 84276 -138410 84284 -138366
rect 84376 -138410 84384 -138366
rect 84476 -138410 84484 -138366
rect 84576 -138410 84584 -138366
rect 84676 -138410 84684 -138366
rect 84776 -138410 84784 -138366
rect 84876 -138410 84884 -138366
rect 84976 -138410 84984 -138366
rect 85076 -138410 85084 -138366
rect 85176 -138410 85184 -138366
rect 85676 -138410 85684 -138366
rect 85776 -138410 85784 -138366
rect 85876 -138410 85884 -138366
rect 85976 -138410 85984 -138366
rect 86076 -138410 86084 -138366
rect 86176 -138410 86184 -138366
rect 86276 -138410 86284 -138366
rect 86376 -138410 86384 -138366
rect 86476 -138410 86484 -138366
rect 86576 -138410 86584 -138366
rect 86676 -138410 86684 -138366
rect 86776 -138410 86784 -138366
rect 86876 -138410 86884 -138366
rect 86976 -138410 86984 -138366
rect 87076 -138410 87084 -138366
rect 87176 -138410 87184 -138366
rect 87676 -138410 87684 -138366
rect 87776 -138410 87784 -138366
rect 87876 -138410 87884 -138366
rect 87976 -138410 87984 -138366
rect 88076 -138410 88084 -138366
rect 88176 -138410 88184 -138366
rect 88276 -138410 88284 -138366
rect 88376 -138410 88384 -138366
rect 88476 -138410 88484 -138366
rect 88576 -138410 88584 -138366
rect 88676 -138410 88684 -138366
rect 88776 -138410 88784 -138366
rect 88876 -138410 88884 -138366
rect 88976 -138410 88984 -138366
rect 89076 -138410 89084 -138366
rect 89176 -138410 89184 -138366
rect 81632 -138466 81676 -138458
rect 81732 -138466 81776 -138458
rect 81832 -138466 81876 -138458
rect 81932 -138466 81976 -138458
rect 82032 -138466 82076 -138458
rect 82132 -138466 82176 -138458
rect 82232 -138466 82276 -138458
rect 82332 -138466 82376 -138458
rect 82432 -138466 82476 -138458
rect 82532 -138466 82576 -138458
rect 82632 -138466 82676 -138458
rect 82732 -138466 82776 -138458
rect 82832 -138466 82876 -138458
rect 82932 -138466 82976 -138458
rect 83032 -138466 83076 -138458
rect 83132 -138466 83176 -138458
rect 83632 -138466 83676 -138458
rect 83732 -138466 83776 -138458
rect 83832 -138466 83876 -138458
rect 83932 -138466 83976 -138458
rect 84032 -138466 84076 -138458
rect 84132 -138466 84176 -138458
rect 84232 -138466 84276 -138458
rect 84332 -138466 84376 -138458
rect 84432 -138466 84476 -138458
rect 84532 -138466 84576 -138458
rect 84632 -138466 84676 -138458
rect 84732 -138466 84776 -138458
rect 84832 -138466 84876 -138458
rect 84932 -138466 84976 -138458
rect 85032 -138466 85076 -138458
rect 85132 -138466 85176 -138458
rect 85632 -138466 85676 -138458
rect 85732 -138466 85776 -138458
rect 85832 -138466 85876 -138458
rect 85932 -138466 85976 -138458
rect 86032 -138466 86076 -138458
rect 86132 -138466 86176 -138458
rect 86232 -138466 86276 -138458
rect 86332 -138466 86376 -138458
rect 86432 -138466 86476 -138458
rect 86532 -138466 86576 -138458
rect 86632 -138466 86676 -138458
rect 86732 -138466 86776 -138458
rect 86832 -138466 86876 -138458
rect 86932 -138466 86976 -138458
rect 87032 -138466 87076 -138458
rect 87132 -138466 87176 -138458
rect 87632 -138466 87676 -138458
rect 87732 -138466 87776 -138458
rect 87832 -138466 87876 -138458
rect 87932 -138466 87976 -138458
rect 88032 -138466 88076 -138458
rect 88132 -138466 88176 -138458
rect 88232 -138466 88276 -138458
rect 88332 -138466 88376 -138458
rect 88432 -138466 88476 -138458
rect 88532 -138466 88576 -138458
rect 88632 -138466 88676 -138458
rect 88732 -138466 88776 -138458
rect 88832 -138466 88876 -138458
rect 88932 -138466 88976 -138458
rect 89032 -138466 89076 -138458
rect 89132 -138466 89176 -138458
rect 81676 -138510 81684 -138466
rect 81776 -138510 81784 -138466
rect 81876 -138510 81884 -138466
rect 81976 -138510 81984 -138466
rect 82076 -138510 82084 -138466
rect 82176 -138510 82184 -138466
rect 82276 -138510 82284 -138466
rect 82376 -138510 82384 -138466
rect 82476 -138510 82484 -138466
rect 82576 -138510 82584 -138466
rect 82676 -138510 82684 -138466
rect 82776 -138510 82784 -138466
rect 82876 -138510 82884 -138466
rect 82976 -138510 82984 -138466
rect 83076 -138510 83084 -138466
rect 83176 -138510 83184 -138466
rect 83676 -138510 83684 -138466
rect 83776 -138510 83784 -138466
rect 83876 -138510 83884 -138466
rect 83976 -138510 83984 -138466
rect 84076 -138510 84084 -138466
rect 84176 -138510 84184 -138466
rect 84276 -138510 84284 -138466
rect 84376 -138510 84384 -138466
rect 84476 -138510 84484 -138466
rect 84576 -138510 84584 -138466
rect 84676 -138510 84684 -138466
rect 84776 -138510 84784 -138466
rect 84876 -138510 84884 -138466
rect 84976 -138510 84984 -138466
rect 85076 -138510 85084 -138466
rect 85176 -138510 85184 -138466
rect 85676 -138510 85684 -138466
rect 85776 -138510 85784 -138466
rect 85876 -138510 85884 -138466
rect 85976 -138510 85984 -138466
rect 86076 -138510 86084 -138466
rect 86176 -138510 86184 -138466
rect 86276 -138510 86284 -138466
rect 86376 -138510 86384 -138466
rect 86476 -138510 86484 -138466
rect 86576 -138510 86584 -138466
rect 86676 -138510 86684 -138466
rect 86776 -138510 86784 -138466
rect 86876 -138510 86884 -138466
rect 86976 -138510 86984 -138466
rect 87076 -138510 87084 -138466
rect 87176 -138510 87184 -138466
rect 87676 -138510 87684 -138466
rect 87776 -138510 87784 -138466
rect 87876 -138510 87884 -138466
rect 87976 -138510 87984 -138466
rect 88076 -138510 88084 -138466
rect 88176 -138510 88184 -138466
rect 88276 -138510 88284 -138466
rect 88376 -138510 88384 -138466
rect 88476 -138510 88484 -138466
rect 88576 -138510 88584 -138466
rect 88676 -138510 88684 -138466
rect 88776 -138510 88784 -138466
rect 88876 -138510 88884 -138466
rect 88976 -138510 88984 -138466
rect 89076 -138510 89084 -138466
rect 89176 -138510 89184 -138466
rect 81632 -138566 81676 -138558
rect 81732 -138566 81776 -138558
rect 81832 -138566 81876 -138558
rect 81932 -138566 81976 -138558
rect 82032 -138566 82076 -138558
rect 82132 -138566 82176 -138558
rect 82232 -138566 82276 -138558
rect 82332 -138566 82376 -138558
rect 82432 -138566 82476 -138558
rect 82532 -138566 82576 -138558
rect 82632 -138566 82676 -138558
rect 82732 -138566 82776 -138558
rect 82832 -138566 82876 -138558
rect 82932 -138566 82976 -138558
rect 83032 -138566 83076 -138558
rect 83132 -138566 83176 -138558
rect 83632 -138566 83676 -138558
rect 83732 -138566 83776 -138558
rect 83832 -138566 83876 -138558
rect 83932 -138566 83976 -138558
rect 84032 -138566 84076 -138558
rect 84132 -138566 84176 -138558
rect 84232 -138566 84276 -138558
rect 84332 -138566 84376 -138558
rect 84432 -138566 84476 -138558
rect 84532 -138566 84576 -138558
rect 84632 -138566 84676 -138558
rect 84732 -138566 84776 -138558
rect 84832 -138566 84876 -138558
rect 84932 -138566 84976 -138558
rect 85032 -138566 85076 -138558
rect 85132 -138566 85176 -138558
rect 85632 -138566 85676 -138558
rect 85732 -138566 85776 -138558
rect 85832 -138566 85876 -138558
rect 85932 -138566 85976 -138558
rect 86032 -138566 86076 -138558
rect 86132 -138566 86176 -138558
rect 86232 -138566 86276 -138558
rect 86332 -138566 86376 -138558
rect 86432 -138566 86476 -138558
rect 86532 -138566 86576 -138558
rect 86632 -138566 86676 -138558
rect 86732 -138566 86776 -138558
rect 86832 -138566 86876 -138558
rect 86932 -138566 86976 -138558
rect 87032 -138566 87076 -138558
rect 87132 -138566 87176 -138558
rect 87632 -138566 87676 -138558
rect 87732 -138566 87776 -138558
rect 87832 -138566 87876 -138558
rect 87932 -138566 87976 -138558
rect 88032 -138566 88076 -138558
rect 88132 -138566 88176 -138558
rect 88232 -138566 88276 -138558
rect 88332 -138566 88376 -138558
rect 88432 -138566 88476 -138558
rect 88532 -138566 88576 -138558
rect 88632 -138566 88676 -138558
rect 88732 -138566 88776 -138558
rect 88832 -138566 88876 -138558
rect 88932 -138566 88976 -138558
rect 89032 -138566 89076 -138558
rect 89132 -138566 89176 -138558
rect 81676 -138610 81684 -138566
rect 81776 -138610 81784 -138566
rect 81876 -138610 81884 -138566
rect 81976 -138610 81984 -138566
rect 82076 -138610 82084 -138566
rect 82176 -138610 82184 -138566
rect 82276 -138610 82284 -138566
rect 82376 -138610 82384 -138566
rect 82476 -138610 82484 -138566
rect 82576 -138610 82584 -138566
rect 82676 -138610 82684 -138566
rect 82776 -138610 82784 -138566
rect 82876 -138610 82884 -138566
rect 82976 -138610 82984 -138566
rect 83076 -138610 83084 -138566
rect 83176 -138610 83184 -138566
rect 83676 -138610 83684 -138566
rect 83776 -138610 83784 -138566
rect 83876 -138610 83884 -138566
rect 83976 -138610 83984 -138566
rect 84076 -138610 84084 -138566
rect 84176 -138610 84184 -138566
rect 84276 -138610 84284 -138566
rect 84376 -138610 84384 -138566
rect 84476 -138610 84484 -138566
rect 84576 -138610 84584 -138566
rect 84676 -138610 84684 -138566
rect 84776 -138610 84784 -138566
rect 84876 -138610 84884 -138566
rect 84976 -138610 84984 -138566
rect 85076 -138610 85084 -138566
rect 85176 -138610 85184 -138566
rect 85676 -138610 85684 -138566
rect 85776 -138610 85784 -138566
rect 85876 -138610 85884 -138566
rect 85976 -138610 85984 -138566
rect 86076 -138610 86084 -138566
rect 86176 -138610 86184 -138566
rect 86276 -138610 86284 -138566
rect 86376 -138610 86384 -138566
rect 86476 -138610 86484 -138566
rect 86576 -138610 86584 -138566
rect 86676 -138610 86684 -138566
rect 86776 -138610 86784 -138566
rect 86876 -138610 86884 -138566
rect 86976 -138610 86984 -138566
rect 87076 -138610 87084 -138566
rect 87176 -138610 87184 -138566
rect 87676 -138610 87684 -138566
rect 87776 -138610 87784 -138566
rect 87876 -138610 87884 -138566
rect 87976 -138610 87984 -138566
rect 88076 -138610 88084 -138566
rect 88176 -138610 88184 -138566
rect 88276 -138610 88284 -138566
rect 88376 -138610 88384 -138566
rect 88476 -138610 88484 -138566
rect 88576 -138610 88584 -138566
rect 88676 -138610 88684 -138566
rect 88776 -138610 88784 -138566
rect 88876 -138610 88884 -138566
rect 88976 -138610 88984 -138566
rect 89076 -138610 89084 -138566
rect 89176 -138610 89184 -138566
rect 81632 -138666 81676 -138658
rect 81732 -138666 81776 -138658
rect 81832 -138666 81876 -138658
rect 81932 -138666 81976 -138658
rect 82032 -138666 82076 -138658
rect 82132 -138666 82176 -138658
rect 82232 -138666 82276 -138658
rect 82332 -138666 82376 -138658
rect 82432 -138666 82476 -138658
rect 82532 -138666 82576 -138658
rect 82632 -138666 82676 -138658
rect 82732 -138666 82776 -138658
rect 82832 -138666 82876 -138658
rect 82932 -138666 82976 -138658
rect 83032 -138666 83076 -138658
rect 83132 -138666 83176 -138658
rect 83632 -138666 83676 -138658
rect 83732 -138666 83776 -138658
rect 83832 -138666 83876 -138658
rect 83932 -138666 83976 -138658
rect 84032 -138666 84076 -138658
rect 84132 -138666 84176 -138658
rect 84232 -138666 84276 -138658
rect 84332 -138666 84376 -138658
rect 84432 -138666 84476 -138658
rect 84532 -138666 84576 -138658
rect 84632 -138666 84676 -138658
rect 84732 -138666 84776 -138658
rect 84832 -138666 84876 -138658
rect 84932 -138666 84976 -138658
rect 85032 -138666 85076 -138658
rect 85132 -138666 85176 -138658
rect 85632 -138666 85676 -138658
rect 85732 -138666 85776 -138658
rect 85832 -138666 85876 -138658
rect 85932 -138666 85976 -138658
rect 86032 -138666 86076 -138658
rect 86132 -138666 86176 -138658
rect 86232 -138666 86276 -138658
rect 86332 -138666 86376 -138658
rect 86432 -138666 86476 -138658
rect 86532 -138666 86576 -138658
rect 86632 -138666 86676 -138658
rect 86732 -138666 86776 -138658
rect 86832 -138666 86876 -138658
rect 86932 -138666 86976 -138658
rect 87032 -138666 87076 -138658
rect 87132 -138666 87176 -138658
rect 87632 -138666 87676 -138658
rect 87732 -138666 87776 -138658
rect 87832 -138666 87876 -138658
rect 87932 -138666 87976 -138658
rect 88032 -138666 88076 -138658
rect 88132 -138666 88176 -138658
rect 88232 -138666 88276 -138658
rect 88332 -138666 88376 -138658
rect 88432 -138666 88476 -138658
rect 88532 -138666 88576 -138658
rect 88632 -138666 88676 -138658
rect 88732 -138666 88776 -138658
rect 88832 -138666 88876 -138658
rect 88932 -138666 88976 -138658
rect 89032 -138666 89076 -138658
rect 89132 -138666 89176 -138658
rect 81676 -138710 81684 -138666
rect 81776 -138710 81784 -138666
rect 81876 -138710 81884 -138666
rect 81976 -138710 81984 -138666
rect 82076 -138710 82084 -138666
rect 82176 -138710 82184 -138666
rect 82276 -138710 82284 -138666
rect 82376 -138710 82384 -138666
rect 82476 -138710 82484 -138666
rect 82576 -138710 82584 -138666
rect 82676 -138710 82684 -138666
rect 82776 -138710 82784 -138666
rect 82876 -138710 82884 -138666
rect 82976 -138710 82984 -138666
rect 83076 -138710 83084 -138666
rect 83176 -138710 83184 -138666
rect 83676 -138710 83684 -138666
rect 83776 -138710 83784 -138666
rect 83876 -138710 83884 -138666
rect 83976 -138710 83984 -138666
rect 84076 -138710 84084 -138666
rect 84176 -138710 84184 -138666
rect 84276 -138710 84284 -138666
rect 84376 -138710 84384 -138666
rect 84476 -138710 84484 -138666
rect 84576 -138710 84584 -138666
rect 84676 -138710 84684 -138666
rect 84776 -138710 84784 -138666
rect 84876 -138710 84884 -138666
rect 84976 -138710 84984 -138666
rect 85076 -138710 85084 -138666
rect 85176 -138710 85184 -138666
rect 85676 -138710 85684 -138666
rect 85776 -138710 85784 -138666
rect 85876 -138710 85884 -138666
rect 85976 -138710 85984 -138666
rect 86076 -138710 86084 -138666
rect 86176 -138710 86184 -138666
rect 86276 -138710 86284 -138666
rect 86376 -138710 86384 -138666
rect 86476 -138710 86484 -138666
rect 86576 -138710 86584 -138666
rect 86676 -138710 86684 -138666
rect 86776 -138710 86784 -138666
rect 86876 -138710 86884 -138666
rect 86976 -138710 86984 -138666
rect 87076 -138710 87084 -138666
rect 87176 -138710 87184 -138666
rect 87676 -138710 87684 -138666
rect 87776 -138710 87784 -138666
rect 87876 -138710 87884 -138666
rect 87976 -138710 87984 -138666
rect 88076 -138710 88084 -138666
rect 88176 -138710 88184 -138666
rect 88276 -138710 88284 -138666
rect 88376 -138710 88384 -138666
rect 88476 -138710 88484 -138666
rect 88576 -138710 88584 -138666
rect 88676 -138710 88684 -138666
rect 88776 -138710 88784 -138666
rect 88876 -138710 88884 -138666
rect 88976 -138710 88984 -138666
rect 89076 -138710 89084 -138666
rect 89176 -138710 89184 -138666
rect 81632 -138766 81676 -138758
rect 81732 -138766 81776 -138758
rect 81832 -138766 81876 -138758
rect 81932 -138766 81976 -138758
rect 82032 -138766 82076 -138758
rect 82132 -138766 82176 -138758
rect 82232 -138766 82276 -138758
rect 82332 -138766 82376 -138758
rect 82432 -138766 82476 -138758
rect 82532 -138766 82576 -138758
rect 82632 -138766 82676 -138758
rect 82732 -138766 82776 -138758
rect 82832 -138766 82876 -138758
rect 82932 -138766 82976 -138758
rect 83032 -138766 83076 -138758
rect 83132 -138766 83176 -138758
rect 83632 -138766 83676 -138758
rect 83732 -138766 83776 -138758
rect 83832 -138766 83876 -138758
rect 83932 -138766 83976 -138758
rect 84032 -138766 84076 -138758
rect 84132 -138766 84176 -138758
rect 84232 -138766 84276 -138758
rect 84332 -138766 84376 -138758
rect 84432 -138766 84476 -138758
rect 84532 -138766 84576 -138758
rect 84632 -138766 84676 -138758
rect 84732 -138766 84776 -138758
rect 84832 -138766 84876 -138758
rect 84932 -138766 84976 -138758
rect 85032 -138766 85076 -138758
rect 85132 -138766 85176 -138758
rect 85632 -138766 85676 -138758
rect 85732 -138766 85776 -138758
rect 85832 -138766 85876 -138758
rect 85932 -138766 85976 -138758
rect 86032 -138766 86076 -138758
rect 86132 -138766 86176 -138758
rect 86232 -138766 86276 -138758
rect 86332 -138766 86376 -138758
rect 86432 -138766 86476 -138758
rect 86532 -138766 86576 -138758
rect 86632 -138766 86676 -138758
rect 86732 -138766 86776 -138758
rect 86832 -138766 86876 -138758
rect 86932 -138766 86976 -138758
rect 87032 -138766 87076 -138758
rect 87132 -138766 87176 -138758
rect 87632 -138766 87676 -138758
rect 87732 -138766 87776 -138758
rect 87832 -138766 87876 -138758
rect 87932 -138766 87976 -138758
rect 88032 -138766 88076 -138758
rect 88132 -138766 88176 -138758
rect 88232 -138766 88276 -138758
rect 88332 -138766 88376 -138758
rect 88432 -138766 88476 -138758
rect 88532 -138766 88576 -138758
rect 88632 -138766 88676 -138758
rect 88732 -138766 88776 -138758
rect 88832 -138766 88876 -138758
rect 88932 -138766 88976 -138758
rect 89032 -138766 89076 -138758
rect 89132 -138766 89176 -138758
rect -105728 -142783 -105726 -138783
rect -105662 -142783 -105660 -138783
rect 81676 -138810 81684 -138766
rect 81776 -138810 81784 -138766
rect 81876 -138810 81884 -138766
rect 81976 -138810 81984 -138766
rect 82076 -138810 82084 -138766
rect 82176 -138810 82184 -138766
rect 82276 -138810 82284 -138766
rect 82376 -138810 82384 -138766
rect 82476 -138810 82484 -138766
rect 82576 -138810 82584 -138766
rect 82676 -138810 82684 -138766
rect 82776 -138810 82784 -138766
rect 82876 -138810 82884 -138766
rect 82976 -138810 82984 -138766
rect 83076 -138810 83084 -138766
rect 83176 -138810 83184 -138766
rect 83676 -138810 83684 -138766
rect 83776 -138810 83784 -138766
rect 83876 -138810 83884 -138766
rect 83976 -138810 83984 -138766
rect 84076 -138810 84084 -138766
rect 84176 -138810 84184 -138766
rect 84276 -138810 84284 -138766
rect 84376 -138810 84384 -138766
rect 84476 -138810 84484 -138766
rect 84576 -138810 84584 -138766
rect 84676 -138810 84684 -138766
rect 84776 -138810 84784 -138766
rect 84876 -138810 84884 -138766
rect 84976 -138810 84984 -138766
rect 85076 -138810 85084 -138766
rect 85176 -138810 85184 -138766
rect 85676 -138810 85684 -138766
rect 85776 -138810 85784 -138766
rect 85876 -138810 85884 -138766
rect 85976 -138810 85984 -138766
rect 86076 -138810 86084 -138766
rect 86176 -138810 86184 -138766
rect 86276 -138810 86284 -138766
rect 86376 -138810 86384 -138766
rect 86476 -138810 86484 -138766
rect 86576 -138810 86584 -138766
rect 86676 -138810 86684 -138766
rect 86776 -138810 86784 -138766
rect 86876 -138810 86884 -138766
rect 86976 -138810 86984 -138766
rect 87076 -138810 87084 -138766
rect 87176 -138810 87184 -138766
rect 87676 -138810 87684 -138766
rect 87776 -138810 87784 -138766
rect 87876 -138810 87884 -138766
rect 87976 -138810 87984 -138766
rect 88076 -138810 88084 -138766
rect 88176 -138810 88184 -138766
rect 88276 -138810 88284 -138766
rect 88376 -138810 88384 -138766
rect 88476 -138810 88484 -138766
rect 88576 -138810 88584 -138766
rect 88676 -138810 88684 -138766
rect 88776 -138810 88784 -138766
rect 88876 -138810 88884 -138766
rect 88976 -138810 88984 -138766
rect 89076 -138810 89084 -138766
rect 89176 -138810 89184 -138766
rect 81632 -138866 81676 -138858
rect 81732 -138866 81776 -138858
rect 81832 -138866 81876 -138858
rect 81932 -138866 81976 -138858
rect 82032 -138866 82076 -138858
rect 82132 -138866 82176 -138858
rect 82232 -138866 82276 -138858
rect 82332 -138866 82376 -138858
rect 82432 -138866 82476 -138858
rect 82532 -138866 82576 -138858
rect 82632 -138866 82676 -138858
rect 82732 -138866 82776 -138858
rect 82832 -138866 82876 -138858
rect 82932 -138866 82976 -138858
rect 83032 -138866 83076 -138858
rect 83132 -138866 83176 -138858
rect 83632 -138866 83676 -138858
rect 83732 -138866 83776 -138858
rect 83832 -138866 83876 -138858
rect 83932 -138866 83976 -138858
rect 84032 -138866 84076 -138858
rect 84132 -138866 84176 -138858
rect 84232 -138866 84276 -138858
rect 84332 -138866 84376 -138858
rect 84432 -138866 84476 -138858
rect 84532 -138866 84576 -138858
rect 84632 -138866 84676 -138858
rect 84732 -138866 84776 -138858
rect 84832 -138866 84876 -138858
rect 84932 -138866 84976 -138858
rect 85032 -138866 85076 -138858
rect 85132 -138866 85176 -138858
rect 85632 -138866 85676 -138858
rect 85732 -138866 85776 -138858
rect 85832 -138866 85876 -138858
rect 85932 -138866 85976 -138858
rect 86032 -138866 86076 -138858
rect 86132 -138866 86176 -138858
rect 86232 -138866 86276 -138858
rect 86332 -138866 86376 -138858
rect 86432 -138866 86476 -138858
rect 86532 -138866 86576 -138858
rect 86632 -138866 86676 -138858
rect 86732 -138866 86776 -138858
rect 86832 -138866 86876 -138858
rect 86932 -138866 86976 -138858
rect 87032 -138866 87076 -138858
rect 87132 -138866 87176 -138858
rect 87632 -138866 87676 -138858
rect 87732 -138866 87776 -138858
rect 87832 -138866 87876 -138858
rect 87932 -138866 87976 -138858
rect 88032 -138866 88076 -138858
rect 88132 -138866 88176 -138858
rect 88232 -138866 88276 -138858
rect 88332 -138866 88376 -138858
rect 88432 -138866 88476 -138858
rect 88532 -138866 88576 -138858
rect 88632 -138866 88676 -138858
rect 88732 -138866 88776 -138858
rect 88832 -138866 88876 -138858
rect 88932 -138866 88976 -138858
rect 89032 -138866 89076 -138858
rect 89132 -138866 89176 -138858
rect 81676 -138910 81684 -138866
rect 81776 -138910 81784 -138866
rect 81876 -138910 81884 -138866
rect 81976 -138910 81984 -138866
rect 82076 -138910 82084 -138866
rect 82176 -138910 82184 -138866
rect 82276 -138910 82284 -138866
rect 82376 -138910 82384 -138866
rect 82476 -138910 82484 -138866
rect 82576 -138910 82584 -138866
rect 82676 -138910 82684 -138866
rect 82776 -138910 82784 -138866
rect 82876 -138910 82884 -138866
rect 82976 -138910 82984 -138866
rect 83076 -138910 83084 -138866
rect 83176 -138910 83184 -138866
rect 83676 -138910 83684 -138866
rect 83776 -138910 83784 -138866
rect 83876 -138910 83884 -138866
rect 83976 -138910 83984 -138866
rect 84076 -138910 84084 -138866
rect 84176 -138910 84184 -138866
rect 84276 -138910 84284 -138866
rect 84376 -138910 84384 -138866
rect 84476 -138910 84484 -138866
rect 84576 -138910 84584 -138866
rect 84676 -138910 84684 -138866
rect 84776 -138910 84784 -138866
rect 84876 -138910 84884 -138866
rect 84976 -138910 84984 -138866
rect 85076 -138910 85084 -138866
rect 85176 -138910 85184 -138866
rect 85676 -138910 85684 -138866
rect 85776 -138910 85784 -138866
rect 85876 -138910 85884 -138866
rect 85976 -138910 85984 -138866
rect 86076 -138910 86084 -138866
rect 86176 -138910 86184 -138866
rect 86276 -138910 86284 -138866
rect 86376 -138910 86384 -138866
rect 86476 -138910 86484 -138866
rect 86576 -138910 86584 -138866
rect 86676 -138910 86684 -138866
rect 86776 -138910 86784 -138866
rect 86876 -138910 86884 -138866
rect 86976 -138910 86984 -138866
rect 87076 -138910 87084 -138866
rect 87176 -138910 87184 -138866
rect 87676 -138910 87684 -138866
rect 87776 -138910 87784 -138866
rect 87876 -138910 87884 -138866
rect 87976 -138910 87984 -138866
rect 88076 -138910 88084 -138866
rect 88176 -138910 88184 -138866
rect 88276 -138910 88284 -138866
rect 88376 -138910 88384 -138866
rect 88476 -138910 88484 -138866
rect 88576 -138910 88584 -138866
rect 88676 -138910 88684 -138866
rect 88776 -138910 88784 -138866
rect 88876 -138910 88884 -138866
rect 88976 -138910 88984 -138866
rect 89076 -138910 89084 -138866
rect 89176 -138910 89184 -138866
rect 81632 -138966 81676 -138958
rect 81732 -138966 81776 -138958
rect 81832 -138966 81876 -138958
rect 81932 -138966 81976 -138958
rect 82032 -138966 82076 -138958
rect 82132 -138966 82176 -138958
rect 82232 -138966 82276 -138958
rect 82332 -138966 82376 -138958
rect 82432 -138966 82476 -138958
rect 82532 -138966 82576 -138958
rect 82632 -138966 82676 -138958
rect 82732 -138966 82776 -138958
rect 82832 -138966 82876 -138958
rect 82932 -138966 82976 -138958
rect 83032 -138966 83076 -138958
rect 83132 -138966 83176 -138958
rect 83632 -138966 83676 -138958
rect 83732 -138966 83776 -138958
rect 83832 -138966 83876 -138958
rect 83932 -138966 83976 -138958
rect 84032 -138966 84076 -138958
rect 84132 -138966 84176 -138958
rect 84232 -138966 84276 -138958
rect 84332 -138966 84376 -138958
rect 84432 -138966 84476 -138958
rect 84532 -138966 84576 -138958
rect 84632 -138966 84676 -138958
rect 84732 -138966 84776 -138958
rect 84832 -138966 84876 -138958
rect 84932 -138966 84976 -138958
rect 85032 -138966 85076 -138958
rect 85132 -138966 85176 -138958
rect 85632 -138966 85676 -138958
rect 85732 -138966 85776 -138958
rect 85832 -138966 85876 -138958
rect 85932 -138966 85976 -138958
rect 86032 -138966 86076 -138958
rect 86132 -138966 86176 -138958
rect 86232 -138966 86276 -138958
rect 86332 -138966 86376 -138958
rect 86432 -138966 86476 -138958
rect 86532 -138966 86576 -138958
rect 86632 -138966 86676 -138958
rect 86732 -138966 86776 -138958
rect 86832 -138966 86876 -138958
rect 86932 -138966 86976 -138958
rect 87032 -138966 87076 -138958
rect 87132 -138966 87176 -138958
rect 87632 -138966 87676 -138958
rect 87732 -138966 87776 -138958
rect 87832 -138966 87876 -138958
rect 87932 -138966 87976 -138958
rect 88032 -138966 88076 -138958
rect 88132 -138966 88176 -138958
rect 88232 -138966 88276 -138958
rect 88332 -138966 88376 -138958
rect 88432 -138966 88476 -138958
rect 88532 -138966 88576 -138958
rect 88632 -138966 88676 -138958
rect 88732 -138966 88776 -138958
rect 88832 -138966 88876 -138958
rect 88932 -138966 88976 -138958
rect 89032 -138966 89076 -138958
rect 89132 -138966 89176 -138958
rect 81676 -139010 81684 -138966
rect 81776 -139010 81784 -138966
rect 81876 -139010 81884 -138966
rect 81976 -139010 81984 -138966
rect 82076 -139010 82084 -138966
rect 82176 -139010 82184 -138966
rect 82276 -139010 82284 -138966
rect 82376 -139010 82384 -138966
rect 82476 -139010 82484 -138966
rect 82576 -139010 82584 -138966
rect 82676 -139010 82684 -138966
rect 82776 -139010 82784 -138966
rect 82876 -139010 82884 -138966
rect 82976 -139010 82984 -138966
rect 83076 -139010 83084 -138966
rect 83176 -139010 83184 -138966
rect 83676 -139010 83684 -138966
rect 83776 -139010 83784 -138966
rect 83876 -139010 83884 -138966
rect 83976 -139010 83984 -138966
rect 84076 -139010 84084 -138966
rect 84176 -139010 84184 -138966
rect 84276 -139010 84284 -138966
rect 84376 -139010 84384 -138966
rect 84476 -139010 84484 -138966
rect 84576 -139010 84584 -138966
rect 84676 -139010 84684 -138966
rect 84776 -139010 84784 -138966
rect 84876 -139010 84884 -138966
rect 84976 -139010 84984 -138966
rect 85076 -139010 85084 -138966
rect 85176 -139010 85184 -138966
rect 85676 -139010 85684 -138966
rect 85776 -139010 85784 -138966
rect 85876 -139010 85884 -138966
rect 85976 -139010 85984 -138966
rect 86076 -139010 86084 -138966
rect 86176 -139010 86184 -138966
rect 86276 -139010 86284 -138966
rect 86376 -139010 86384 -138966
rect 86476 -139010 86484 -138966
rect 86576 -139010 86584 -138966
rect 86676 -139010 86684 -138966
rect 86776 -139010 86784 -138966
rect 86876 -139010 86884 -138966
rect 86976 -139010 86984 -138966
rect 87076 -139010 87084 -138966
rect 87176 -139010 87184 -138966
rect 87676 -139010 87684 -138966
rect 87776 -139010 87784 -138966
rect 87876 -139010 87884 -138966
rect 87976 -139010 87984 -138966
rect 88076 -139010 88084 -138966
rect 88176 -139010 88184 -138966
rect 88276 -139010 88284 -138966
rect 88376 -139010 88384 -138966
rect 88476 -139010 88484 -138966
rect 88576 -139010 88584 -138966
rect 88676 -139010 88684 -138966
rect 88776 -139010 88784 -138966
rect 88876 -139010 88884 -138966
rect 88976 -139010 88984 -138966
rect 89076 -139010 89084 -138966
rect 89176 -139010 89184 -138966
rect 81632 -139066 81676 -139058
rect 81732 -139066 81776 -139058
rect 81832 -139066 81876 -139058
rect 81932 -139066 81976 -139058
rect 82032 -139066 82076 -139058
rect 82132 -139066 82176 -139058
rect 82232 -139066 82276 -139058
rect 82332 -139066 82376 -139058
rect 82432 -139066 82476 -139058
rect 82532 -139066 82576 -139058
rect 82632 -139066 82676 -139058
rect 82732 -139066 82776 -139058
rect 82832 -139066 82876 -139058
rect 82932 -139066 82976 -139058
rect 83032 -139066 83076 -139058
rect 83132 -139066 83176 -139058
rect 83632 -139066 83676 -139058
rect 83732 -139066 83776 -139058
rect 83832 -139066 83876 -139058
rect 83932 -139066 83976 -139058
rect 84032 -139066 84076 -139058
rect 84132 -139066 84176 -139058
rect 84232 -139066 84276 -139058
rect 84332 -139066 84376 -139058
rect 84432 -139066 84476 -139058
rect 84532 -139066 84576 -139058
rect 84632 -139066 84676 -139058
rect 84732 -139066 84776 -139058
rect 84832 -139066 84876 -139058
rect 84932 -139066 84976 -139058
rect 85032 -139066 85076 -139058
rect 85132 -139066 85176 -139058
rect 85632 -139066 85676 -139058
rect 85732 -139066 85776 -139058
rect 85832 -139066 85876 -139058
rect 85932 -139066 85976 -139058
rect 86032 -139066 86076 -139058
rect 86132 -139066 86176 -139058
rect 86232 -139066 86276 -139058
rect 86332 -139066 86376 -139058
rect 86432 -139066 86476 -139058
rect 86532 -139066 86576 -139058
rect 86632 -139066 86676 -139058
rect 86732 -139066 86776 -139058
rect 86832 -139066 86876 -139058
rect 86932 -139066 86976 -139058
rect 87032 -139066 87076 -139058
rect 87132 -139066 87176 -139058
rect 87632 -139066 87676 -139058
rect 87732 -139066 87776 -139058
rect 87832 -139066 87876 -139058
rect 87932 -139066 87976 -139058
rect 88032 -139066 88076 -139058
rect 88132 -139066 88176 -139058
rect 88232 -139066 88276 -139058
rect 88332 -139066 88376 -139058
rect 88432 -139066 88476 -139058
rect 88532 -139066 88576 -139058
rect 88632 -139066 88676 -139058
rect 88732 -139066 88776 -139058
rect 88832 -139066 88876 -139058
rect 88932 -139066 88976 -139058
rect 89032 -139066 89076 -139058
rect 89132 -139066 89176 -139058
rect 81676 -139110 81684 -139066
rect 81776 -139110 81784 -139066
rect 81876 -139110 81884 -139066
rect 81976 -139110 81984 -139066
rect 82076 -139110 82084 -139066
rect 82176 -139110 82184 -139066
rect 82276 -139110 82284 -139066
rect 82376 -139110 82384 -139066
rect 82476 -139110 82484 -139066
rect 82576 -139110 82584 -139066
rect 82676 -139110 82684 -139066
rect 82776 -139110 82784 -139066
rect 82876 -139110 82884 -139066
rect 82976 -139110 82984 -139066
rect 83076 -139110 83084 -139066
rect 83176 -139110 83184 -139066
rect 83676 -139110 83684 -139066
rect 83776 -139110 83784 -139066
rect 83876 -139110 83884 -139066
rect 83976 -139110 83984 -139066
rect 84076 -139110 84084 -139066
rect 84176 -139110 84184 -139066
rect 84276 -139110 84284 -139066
rect 84376 -139110 84384 -139066
rect 84476 -139110 84484 -139066
rect 84576 -139110 84584 -139066
rect 84676 -139110 84684 -139066
rect 84776 -139110 84784 -139066
rect 84876 -139110 84884 -139066
rect 84976 -139110 84984 -139066
rect 85076 -139110 85084 -139066
rect 85176 -139110 85184 -139066
rect 85676 -139110 85684 -139066
rect 85776 -139110 85784 -139066
rect 85876 -139110 85884 -139066
rect 85976 -139110 85984 -139066
rect 86076 -139110 86084 -139066
rect 86176 -139110 86184 -139066
rect 86276 -139110 86284 -139066
rect 86376 -139110 86384 -139066
rect 86476 -139110 86484 -139066
rect 86576 -139110 86584 -139066
rect 86676 -139110 86684 -139066
rect 86776 -139110 86784 -139066
rect 86876 -139110 86884 -139066
rect 86976 -139110 86984 -139066
rect 87076 -139110 87084 -139066
rect 87176 -139110 87184 -139066
rect 87676 -139110 87684 -139066
rect 87776 -139110 87784 -139066
rect 87876 -139110 87884 -139066
rect 87976 -139110 87984 -139066
rect 88076 -139110 88084 -139066
rect 88176 -139110 88184 -139066
rect 88276 -139110 88284 -139066
rect 88376 -139110 88384 -139066
rect 88476 -139110 88484 -139066
rect 88576 -139110 88584 -139066
rect 88676 -139110 88684 -139066
rect 88776 -139110 88784 -139066
rect 88876 -139110 88884 -139066
rect 88976 -139110 88984 -139066
rect 89076 -139110 89084 -139066
rect 89176 -139110 89184 -139066
rect 81632 -139166 81676 -139158
rect 81732 -139166 81776 -139158
rect 81832 -139166 81876 -139158
rect 81932 -139166 81976 -139158
rect 82032 -139166 82076 -139158
rect 82132 -139166 82176 -139158
rect 82232 -139166 82276 -139158
rect 82332 -139166 82376 -139158
rect 82432 -139166 82476 -139158
rect 82532 -139166 82576 -139158
rect 82632 -139166 82676 -139158
rect 82732 -139166 82776 -139158
rect 82832 -139166 82876 -139158
rect 82932 -139166 82976 -139158
rect 83032 -139166 83076 -139158
rect 83132 -139166 83176 -139158
rect 83632 -139166 83676 -139158
rect 83732 -139166 83776 -139158
rect 83832 -139166 83876 -139158
rect 83932 -139166 83976 -139158
rect 84032 -139166 84076 -139158
rect 84132 -139166 84176 -139158
rect 84232 -139166 84276 -139158
rect 84332 -139166 84376 -139158
rect 84432 -139166 84476 -139158
rect 84532 -139166 84576 -139158
rect 84632 -139166 84676 -139158
rect 84732 -139166 84776 -139158
rect 84832 -139166 84876 -139158
rect 84932 -139166 84976 -139158
rect 85032 -139166 85076 -139158
rect 85132 -139166 85176 -139158
rect 85632 -139166 85676 -139158
rect 85732 -139166 85776 -139158
rect 85832 -139166 85876 -139158
rect 85932 -139166 85976 -139158
rect 86032 -139166 86076 -139158
rect 86132 -139166 86176 -139158
rect 86232 -139166 86276 -139158
rect 86332 -139166 86376 -139158
rect 86432 -139166 86476 -139158
rect 86532 -139166 86576 -139158
rect 86632 -139166 86676 -139158
rect 86732 -139166 86776 -139158
rect 86832 -139166 86876 -139158
rect 86932 -139166 86976 -139158
rect 87032 -139166 87076 -139158
rect 87132 -139166 87176 -139158
rect 87632 -139166 87676 -139158
rect 87732 -139166 87776 -139158
rect 87832 -139166 87876 -139158
rect 87932 -139166 87976 -139158
rect 88032 -139166 88076 -139158
rect 88132 -139166 88176 -139158
rect 88232 -139166 88276 -139158
rect 88332 -139166 88376 -139158
rect 88432 -139166 88476 -139158
rect 88532 -139166 88576 -139158
rect 88632 -139166 88676 -139158
rect 88732 -139166 88776 -139158
rect 88832 -139166 88876 -139158
rect 88932 -139166 88976 -139158
rect 89032 -139166 89076 -139158
rect 89132 -139166 89176 -139158
rect 81676 -139210 81684 -139166
rect 81776 -139210 81784 -139166
rect 81876 -139210 81884 -139166
rect 81976 -139210 81984 -139166
rect 82076 -139210 82084 -139166
rect 82176 -139210 82184 -139166
rect 82276 -139210 82284 -139166
rect 82376 -139210 82384 -139166
rect 82476 -139210 82484 -139166
rect 82576 -139210 82584 -139166
rect 82676 -139210 82684 -139166
rect 82776 -139210 82784 -139166
rect 82876 -139210 82884 -139166
rect 82976 -139210 82984 -139166
rect 83076 -139210 83084 -139166
rect 83176 -139210 83184 -139166
rect 83676 -139210 83684 -139166
rect 83776 -139210 83784 -139166
rect 83876 -139210 83884 -139166
rect 83976 -139210 83984 -139166
rect 84076 -139210 84084 -139166
rect 84176 -139210 84184 -139166
rect 84276 -139210 84284 -139166
rect 84376 -139210 84384 -139166
rect 84476 -139210 84484 -139166
rect 84576 -139210 84584 -139166
rect 84676 -139210 84684 -139166
rect 84776 -139210 84784 -139166
rect 84876 -139210 84884 -139166
rect 84976 -139210 84984 -139166
rect 85076 -139210 85084 -139166
rect 85176 -139210 85184 -139166
rect 85676 -139210 85684 -139166
rect 85776 -139210 85784 -139166
rect 85876 -139210 85884 -139166
rect 85976 -139210 85984 -139166
rect 86076 -139210 86084 -139166
rect 86176 -139210 86184 -139166
rect 86276 -139210 86284 -139166
rect 86376 -139210 86384 -139166
rect 86476 -139210 86484 -139166
rect 86576 -139210 86584 -139166
rect 86676 -139210 86684 -139166
rect 86776 -139210 86784 -139166
rect 86876 -139210 86884 -139166
rect 86976 -139210 86984 -139166
rect 87076 -139210 87084 -139166
rect 87176 -139210 87184 -139166
rect 87676 -139210 87684 -139166
rect 87776 -139210 87784 -139166
rect 87876 -139210 87884 -139166
rect 87976 -139210 87984 -139166
rect 88076 -139210 88084 -139166
rect 88176 -139210 88184 -139166
rect 88276 -139210 88284 -139166
rect 88376 -139210 88384 -139166
rect 88476 -139210 88484 -139166
rect 88576 -139210 88584 -139166
rect 88676 -139210 88684 -139166
rect 88776 -139210 88784 -139166
rect 88876 -139210 88884 -139166
rect 88976 -139210 88984 -139166
rect 89076 -139210 89084 -139166
rect 89176 -139210 89184 -139166
rect 81632 -139266 81676 -139258
rect 81732 -139266 81776 -139258
rect 81832 -139266 81876 -139258
rect 81932 -139266 81976 -139258
rect 82032 -139266 82076 -139258
rect 82132 -139266 82176 -139258
rect 82232 -139266 82276 -139258
rect 82332 -139266 82376 -139258
rect 82432 -139266 82476 -139258
rect 82532 -139266 82576 -139258
rect 82632 -139266 82676 -139258
rect 82732 -139266 82776 -139258
rect 82832 -139266 82876 -139258
rect 82932 -139266 82976 -139258
rect 83032 -139266 83076 -139258
rect 83132 -139266 83176 -139258
rect 83632 -139266 83676 -139258
rect 83732 -139266 83776 -139258
rect 83832 -139266 83876 -139258
rect 83932 -139266 83976 -139258
rect 84032 -139266 84076 -139258
rect 84132 -139266 84176 -139258
rect 84232 -139266 84276 -139258
rect 84332 -139266 84376 -139258
rect 84432 -139266 84476 -139258
rect 84532 -139266 84576 -139258
rect 84632 -139266 84676 -139258
rect 84732 -139266 84776 -139258
rect 84832 -139266 84876 -139258
rect 84932 -139266 84976 -139258
rect 85032 -139266 85076 -139258
rect 85132 -139266 85176 -139258
rect 85632 -139266 85676 -139258
rect 85732 -139266 85776 -139258
rect 85832 -139266 85876 -139258
rect 85932 -139266 85976 -139258
rect 86032 -139266 86076 -139258
rect 86132 -139266 86176 -139258
rect 86232 -139266 86276 -139258
rect 86332 -139266 86376 -139258
rect 86432 -139266 86476 -139258
rect 86532 -139266 86576 -139258
rect 86632 -139266 86676 -139258
rect 86732 -139266 86776 -139258
rect 86832 -139266 86876 -139258
rect 86932 -139266 86976 -139258
rect 87032 -139266 87076 -139258
rect 87132 -139266 87176 -139258
rect 87632 -139266 87676 -139258
rect 87732 -139266 87776 -139258
rect 87832 -139266 87876 -139258
rect 87932 -139266 87976 -139258
rect 88032 -139266 88076 -139258
rect 88132 -139266 88176 -139258
rect 88232 -139266 88276 -139258
rect 88332 -139266 88376 -139258
rect 88432 -139266 88476 -139258
rect 88532 -139266 88576 -139258
rect 88632 -139266 88676 -139258
rect 88732 -139266 88776 -139258
rect 88832 -139266 88876 -139258
rect 88932 -139266 88976 -139258
rect 89032 -139266 89076 -139258
rect 89132 -139266 89176 -139258
rect 81676 -139310 81684 -139266
rect 81776 -139310 81784 -139266
rect 81876 -139310 81884 -139266
rect 81976 -139310 81984 -139266
rect 82076 -139310 82084 -139266
rect 82176 -139310 82184 -139266
rect 82276 -139310 82284 -139266
rect 82376 -139310 82384 -139266
rect 82476 -139310 82484 -139266
rect 82576 -139310 82584 -139266
rect 82676 -139310 82684 -139266
rect 82776 -139310 82784 -139266
rect 82876 -139310 82884 -139266
rect 82976 -139310 82984 -139266
rect 83076 -139310 83084 -139266
rect 83176 -139310 83184 -139266
rect 83676 -139310 83684 -139266
rect 83776 -139310 83784 -139266
rect 83876 -139310 83884 -139266
rect 83976 -139310 83984 -139266
rect 84076 -139310 84084 -139266
rect 84176 -139310 84184 -139266
rect 84276 -139310 84284 -139266
rect 84376 -139310 84384 -139266
rect 84476 -139310 84484 -139266
rect 84576 -139310 84584 -139266
rect 84676 -139310 84684 -139266
rect 84776 -139310 84784 -139266
rect 84876 -139310 84884 -139266
rect 84976 -139310 84984 -139266
rect 85076 -139310 85084 -139266
rect 85176 -139310 85184 -139266
rect 85676 -139310 85684 -139266
rect 85776 -139310 85784 -139266
rect 85876 -139310 85884 -139266
rect 85976 -139310 85984 -139266
rect 86076 -139310 86084 -139266
rect 86176 -139310 86184 -139266
rect 86276 -139310 86284 -139266
rect 86376 -139310 86384 -139266
rect 86476 -139310 86484 -139266
rect 86576 -139310 86584 -139266
rect 86676 -139310 86684 -139266
rect 86776 -139310 86784 -139266
rect 86876 -139310 86884 -139266
rect 86976 -139310 86984 -139266
rect 87076 -139310 87084 -139266
rect 87176 -139310 87184 -139266
rect 87676 -139310 87684 -139266
rect 87776 -139310 87784 -139266
rect 87876 -139310 87884 -139266
rect 87976 -139310 87984 -139266
rect 88076 -139310 88084 -139266
rect 88176 -139310 88184 -139266
rect 88276 -139310 88284 -139266
rect 88376 -139310 88384 -139266
rect 88476 -139310 88484 -139266
rect 88576 -139310 88584 -139266
rect 88676 -139310 88684 -139266
rect 88776 -139310 88784 -139266
rect 88876 -139310 88884 -139266
rect 88976 -139310 88984 -139266
rect 89076 -139310 89084 -139266
rect 89176 -139310 89184 -139266
rect 81632 -139366 81676 -139358
rect 81732 -139366 81776 -139358
rect 81832 -139366 81876 -139358
rect 81932 -139366 81976 -139358
rect 82032 -139366 82076 -139358
rect 82132 -139366 82176 -139358
rect 82232 -139366 82276 -139358
rect 82332 -139366 82376 -139358
rect 82432 -139366 82476 -139358
rect 82532 -139366 82576 -139358
rect 82632 -139366 82676 -139358
rect 82732 -139366 82776 -139358
rect 82832 -139366 82876 -139358
rect 82932 -139366 82976 -139358
rect 83032 -139366 83076 -139358
rect 83132 -139366 83176 -139358
rect 83632 -139366 83676 -139358
rect 83732 -139366 83776 -139358
rect 83832 -139366 83876 -139358
rect 83932 -139366 83976 -139358
rect 84032 -139366 84076 -139358
rect 84132 -139366 84176 -139358
rect 84232 -139366 84276 -139358
rect 84332 -139366 84376 -139358
rect 84432 -139366 84476 -139358
rect 84532 -139366 84576 -139358
rect 84632 -139366 84676 -139358
rect 84732 -139366 84776 -139358
rect 84832 -139366 84876 -139358
rect 84932 -139366 84976 -139358
rect 85032 -139366 85076 -139358
rect 85132 -139366 85176 -139358
rect 85632 -139366 85676 -139358
rect 85732 -139366 85776 -139358
rect 85832 -139366 85876 -139358
rect 85932 -139366 85976 -139358
rect 86032 -139366 86076 -139358
rect 86132 -139366 86176 -139358
rect 86232 -139366 86276 -139358
rect 86332 -139366 86376 -139358
rect 86432 -139366 86476 -139358
rect 86532 -139366 86576 -139358
rect 86632 -139366 86676 -139358
rect 86732 -139366 86776 -139358
rect 86832 -139366 86876 -139358
rect 86932 -139366 86976 -139358
rect 87032 -139366 87076 -139358
rect 87132 -139366 87176 -139358
rect 87632 -139366 87676 -139358
rect 87732 -139366 87776 -139358
rect 87832 -139366 87876 -139358
rect 87932 -139366 87976 -139358
rect 88032 -139366 88076 -139358
rect 88132 -139366 88176 -139358
rect 88232 -139366 88276 -139358
rect 88332 -139366 88376 -139358
rect 88432 -139366 88476 -139358
rect 88532 -139366 88576 -139358
rect 88632 -139366 88676 -139358
rect 88732 -139366 88776 -139358
rect 88832 -139366 88876 -139358
rect 88932 -139366 88976 -139358
rect 89032 -139366 89076 -139358
rect 89132 -139366 89176 -139358
rect 81676 -139410 81684 -139366
rect 81776 -139410 81784 -139366
rect 81876 -139410 81884 -139366
rect 81976 -139410 81984 -139366
rect 82076 -139410 82084 -139366
rect 82176 -139410 82184 -139366
rect 82276 -139410 82284 -139366
rect 82376 -139410 82384 -139366
rect 82476 -139410 82484 -139366
rect 82576 -139410 82584 -139366
rect 82676 -139410 82684 -139366
rect 82776 -139410 82784 -139366
rect 82876 -139410 82884 -139366
rect 82976 -139410 82984 -139366
rect 83076 -139410 83084 -139366
rect 83176 -139410 83184 -139366
rect 83676 -139410 83684 -139366
rect 83776 -139410 83784 -139366
rect 83876 -139410 83884 -139366
rect 83976 -139410 83984 -139366
rect 84076 -139410 84084 -139366
rect 84176 -139410 84184 -139366
rect 84276 -139410 84284 -139366
rect 84376 -139410 84384 -139366
rect 84476 -139410 84484 -139366
rect 84576 -139410 84584 -139366
rect 84676 -139410 84684 -139366
rect 84776 -139410 84784 -139366
rect 84876 -139410 84884 -139366
rect 84976 -139410 84984 -139366
rect 85076 -139410 85084 -139366
rect 85176 -139410 85184 -139366
rect 85676 -139410 85684 -139366
rect 85776 -139410 85784 -139366
rect 85876 -139410 85884 -139366
rect 85976 -139410 85984 -139366
rect 86076 -139410 86084 -139366
rect 86176 -139410 86184 -139366
rect 86276 -139410 86284 -139366
rect 86376 -139410 86384 -139366
rect 86476 -139410 86484 -139366
rect 86576 -139410 86584 -139366
rect 86676 -139410 86684 -139366
rect 86776 -139410 86784 -139366
rect 86876 -139410 86884 -139366
rect 86976 -139410 86984 -139366
rect 87076 -139410 87084 -139366
rect 87176 -139410 87184 -139366
rect 87676 -139410 87684 -139366
rect 87776 -139410 87784 -139366
rect 87876 -139410 87884 -139366
rect 87976 -139410 87984 -139366
rect 88076 -139410 88084 -139366
rect 88176 -139410 88184 -139366
rect 88276 -139410 88284 -139366
rect 88376 -139410 88384 -139366
rect 88476 -139410 88484 -139366
rect 88576 -139410 88584 -139366
rect 88676 -139410 88684 -139366
rect 88776 -139410 88784 -139366
rect 88876 -139410 88884 -139366
rect 88976 -139410 88984 -139366
rect 89076 -139410 89084 -139366
rect 89176 -139410 89184 -139366
rect 81632 -139466 81676 -139458
rect 81732 -139466 81776 -139458
rect 81832 -139466 81876 -139458
rect 81932 -139466 81976 -139458
rect 82032 -139466 82076 -139458
rect 82132 -139466 82176 -139458
rect 82232 -139466 82276 -139458
rect 82332 -139466 82376 -139458
rect 82432 -139466 82476 -139458
rect 82532 -139466 82576 -139458
rect 82632 -139466 82676 -139458
rect 82732 -139466 82776 -139458
rect 82832 -139466 82876 -139458
rect 82932 -139466 82976 -139458
rect 83032 -139466 83076 -139458
rect 83132 -139466 83176 -139458
rect 83632 -139466 83676 -139458
rect 83732 -139466 83776 -139458
rect 83832 -139466 83876 -139458
rect 83932 -139466 83976 -139458
rect 84032 -139466 84076 -139458
rect 84132 -139466 84176 -139458
rect 84232 -139466 84276 -139458
rect 84332 -139466 84376 -139458
rect 84432 -139466 84476 -139458
rect 84532 -139466 84576 -139458
rect 84632 -139466 84676 -139458
rect 84732 -139466 84776 -139458
rect 84832 -139466 84876 -139458
rect 84932 -139466 84976 -139458
rect 85032 -139466 85076 -139458
rect 85132 -139466 85176 -139458
rect 85632 -139466 85676 -139458
rect 85732 -139466 85776 -139458
rect 85832 -139466 85876 -139458
rect 85932 -139466 85976 -139458
rect 86032 -139466 86076 -139458
rect 86132 -139466 86176 -139458
rect 86232 -139466 86276 -139458
rect 86332 -139466 86376 -139458
rect 86432 -139466 86476 -139458
rect 86532 -139466 86576 -139458
rect 86632 -139466 86676 -139458
rect 86732 -139466 86776 -139458
rect 86832 -139466 86876 -139458
rect 86932 -139466 86976 -139458
rect 87032 -139466 87076 -139458
rect 87132 -139466 87176 -139458
rect 87632 -139466 87676 -139458
rect 87732 -139466 87776 -139458
rect 87832 -139466 87876 -139458
rect 87932 -139466 87976 -139458
rect 88032 -139466 88076 -139458
rect 88132 -139466 88176 -139458
rect 88232 -139466 88276 -139458
rect 88332 -139466 88376 -139458
rect 88432 -139466 88476 -139458
rect 88532 -139466 88576 -139458
rect 88632 -139466 88676 -139458
rect 88732 -139466 88776 -139458
rect 88832 -139466 88876 -139458
rect 88932 -139466 88976 -139458
rect 89032 -139466 89076 -139458
rect 89132 -139466 89176 -139458
rect 81676 -139510 81684 -139466
rect 81776 -139510 81784 -139466
rect 81876 -139510 81884 -139466
rect 81976 -139510 81984 -139466
rect 82076 -139510 82084 -139466
rect 82176 -139510 82184 -139466
rect 82276 -139510 82284 -139466
rect 82376 -139510 82384 -139466
rect 82476 -139510 82484 -139466
rect 82576 -139510 82584 -139466
rect 82676 -139510 82684 -139466
rect 82776 -139510 82784 -139466
rect 82876 -139510 82884 -139466
rect 82976 -139510 82984 -139466
rect 83076 -139510 83084 -139466
rect 83176 -139510 83184 -139466
rect 83676 -139510 83684 -139466
rect 83776 -139510 83784 -139466
rect 83876 -139510 83884 -139466
rect 83976 -139510 83984 -139466
rect 84076 -139510 84084 -139466
rect 84176 -139510 84184 -139466
rect 84276 -139510 84284 -139466
rect 84376 -139510 84384 -139466
rect 84476 -139510 84484 -139466
rect 84576 -139510 84584 -139466
rect 84676 -139510 84684 -139466
rect 84776 -139510 84784 -139466
rect 84876 -139510 84884 -139466
rect 84976 -139510 84984 -139466
rect 85076 -139510 85084 -139466
rect 85176 -139510 85184 -139466
rect 85676 -139510 85684 -139466
rect 85776 -139510 85784 -139466
rect 85876 -139510 85884 -139466
rect 85976 -139510 85984 -139466
rect 86076 -139510 86084 -139466
rect 86176 -139510 86184 -139466
rect 86276 -139510 86284 -139466
rect 86376 -139510 86384 -139466
rect 86476 -139510 86484 -139466
rect 86576 -139510 86584 -139466
rect 86676 -139510 86684 -139466
rect 86776 -139510 86784 -139466
rect 86876 -139510 86884 -139466
rect 86976 -139510 86984 -139466
rect 87076 -139510 87084 -139466
rect 87176 -139510 87184 -139466
rect 87676 -139510 87684 -139466
rect 87776 -139510 87784 -139466
rect 87876 -139510 87884 -139466
rect 87976 -139510 87984 -139466
rect 88076 -139510 88084 -139466
rect 88176 -139510 88184 -139466
rect 88276 -139510 88284 -139466
rect 88376 -139510 88384 -139466
rect 88476 -139510 88484 -139466
rect 88576 -139510 88584 -139466
rect 88676 -139510 88684 -139466
rect 88776 -139510 88784 -139466
rect 88876 -139510 88884 -139466
rect 88976 -139510 88984 -139466
rect 89076 -139510 89084 -139466
rect 89176 -139510 89184 -139466
rect -83265 -140231 -83221 -140223
rect -83165 -140231 -83121 -140223
rect -83065 -140231 -83021 -140223
rect -82965 -140231 -82921 -140223
rect -82865 -140231 -82821 -140223
rect -82765 -140231 -82721 -140223
rect -82665 -140231 -82621 -140223
rect -82565 -140231 -82521 -140223
rect -82465 -140231 -82421 -140223
rect -82365 -140231 -82321 -140223
rect -82265 -140231 -82221 -140223
rect -82165 -140231 -82121 -140223
rect -82065 -140231 -82021 -140223
rect -81965 -140231 -81921 -140223
rect -81865 -140231 -81821 -140223
rect -81765 -140231 -81721 -140223
rect -81265 -140231 -81221 -140223
rect -81165 -140231 -81121 -140223
rect -81065 -140231 -81021 -140223
rect -80965 -140231 -80921 -140223
rect -80865 -140231 -80821 -140223
rect -80765 -140231 -80721 -140223
rect -80665 -140231 -80621 -140223
rect -80565 -140231 -80521 -140223
rect -80465 -140231 -80421 -140223
rect -80365 -140231 -80321 -140223
rect -80265 -140231 -80221 -140223
rect -80165 -140231 -80121 -140223
rect -80065 -140231 -80021 -140223
rect -79965 -140231 -79921 -140223
rect -79865 -140231 -79821 -140223
rect -79765 -140231 -79721 -140223
rect -79265 -140231 -79221 -140223
rect -79165 -140231 -79121 -140223
rect -79065 -140231 -79021 -140223
rect -78965 -140231 -78921 -140223
rect -78865 -140231 -78821 -140223
rect -78765 -140231 -78721 -140223
rect -78665 -140231 -78621 -140223
rect -78565 -140231 -78521 -140223
rect -78465 -140231 -78421 -140223
rect -78365 -140231 -78321 -140223
rect -78265 -140231 -78221 -140223
rect -78165 -140231 -78121 -140223
rect -78065 -140231 -78021 -140223
rect -77965 -140231 -77921 -140223
rect -77865 -140231 -77821 -140223
rect -77765 -140231 -77721 -140223
rect -77265 -140231 -77221 -140223
rect -77165 -140231 -77121 -140223
rect -77065 -140231 -77021 -140223
rect -76965 -140231 -76921 -140223
rect -76865 -140231 -76821 -140223
rect -76765 -140231 -76721 -140223
rect -76665 -140231 -76621 -140223
rect -76565 -140231 -76521 -140223
rect -76465 -140231 -76421 -140223
rect -76365 -140231 -76321 -140223
rect -76265 -140231 -76221 -140223
rect -76165 -140231 -76121 -140223
rect -76065 -140231 -76021 -140223
rect -75965 -140231 -75921 -140223
rect -75865 -140231 -75821 -140223
rect -75765 -140231 -75721 -140223
rect -83221 -140275 -83213 -140231
rect -83121 -140275 -83113 -140231
rect -83021 -140275 -83013 -140231
rect -82921 -140275 -82913 -140231
rect -82821 -140275 -82813 -140231
rect -82721 -140275 -82713 -140231
rect -82621 -140275 -82613 -140231
rect -82521 -140275 -82513 -140231
rect -82421 -140275 -82413 -140231
rect -82321 -140275 -82313 -140231
rect -82221 -140275 -82213 -140231
rect -82121 -140275 -82113 -140231
rect -82021 -140275 -82013 -140231
rect -81921 -140275 -81913 -140231
rect -81821 -140275 -81813 -140231
rect -81721 -140275 -81713 -140231
rect -81221 -140275 -81213 -140231
rect -81121 -140275 -81113 -140231
rect -81021 -140275 -81013 -140231
rect -80921 -140275 -80913 -140231
rect -80821 -140275 -80813 -140231
rect -80721 -140275 -80713 -140231
rect -80621 -140275 -80613 -140231
rect -80521 -140275 -80513 -140231
rect -80421 -140275 -80413 -140231
rect -80321 -140275 -80313 -140231
rect -80221 -140275 -80213 -140231
rect -80121 -140275 -80113 -140231
rect -80021 -140275 -80013 -140231
rect -79921 -140275 -79913 -140231
rect -79821 -140275 -79813 -140231
rect -79721 -140275 -79713 -140231
rect -79221 -140275 -79213 -140231
rect -79121 -140275 -79113 -140231
rect -79021 -140275 -79013 -140231
rect -78921 -140275 -78913 -140231
rect -78821 -140275 -78813 -140231
rect -78721 -140275 -78713 -140231
rect -78621 -140275 -78613 -140231
rect -78521 -140275 -78513 -140231
rect -78421 -140275 -78413 -140231
rect -78321 -140275 -78313 -140231
rect -78221 -140275 -78213 -140231
rect -78121 -140275 -78113 -140231
rect -78021 -140275 -78013 -140231
rect -77921 -140275 -77913 -140231
rect -77821 -140275 -77813 -140231
rect -77721 -140275 -77713 -140231
rect -77221 -140275 -77213 -140231
rect -77121 -140275 -77113 -140231
rect -77021 -140275 -77013 -140231
rect -76921 -140275 -76913 -140231
rect -76821 -140275 -76813 -140231
rect -76721 -140275 -76713 -140231
rect -76621 -140275 -76613 -140231
rect -76521 -140275 -76513 -140231
rect -76421 -140275 -76413 -140231
rect -76321 -140275 -76313 -140231
rect -76221 -140275 -76213 -140231
rect -76121 -140275 -76113 -140231
rect -76021 -140275 -76013 -140231
rect -75921 -140275 -75913 -140231
rect -75821 -140275 -75813 -140231
rect -75721 -140275 -75713 -140231
rect -83265 -140331 -83221 -140323
rect -83165 -140331 -83121 -140323
rect -83065 -140331 -83021 -140323
rect -82965 -140331 -82921 -140323
rect -82865 -140331 -82821 -140323
rect -82765 -140331 -82721 -140323
rect -82665 -140331 -82621 -140323
rect -82565 -140331 -82521 -140323
rect -82465 -140331 -82421 -140323
rect -82365 -140331 -82321 -140323
rect -82265 -140331 -82221 -140323
rect -82165 -140331 -82121 -140323
rect -82065 -140331 -82021 -140323
rect -81965 -140331 -81921 -140323
rect -81865 -140331 -81821 -140323
rect -81765 -140331 -81721 -140323
rect -81265 -140331 -81221 -140323
rect -81165 -140331 -81121 -140323
rect -81065 -140331 -81021 -140323
rect -80965 -140331 -80921 -140323
rect -80865 -140331 -80821 -140323
rect -80765 -140331 -80721 -140323
rect -80665 -140331 -80621 -140323
rect -80565 -140331 -80521 -140323
rect -80465 -140331 -80421 -140323
rect -80365 -140331 -80321 -140323
rect -80265 -140331 -80221 -140323
rect -80165 -140331 -80121 -140323
rect -80065 -140331 -80021 -140323
rect -79965 -140331 -79921 -140323
rect -79865 -140331 -79821 -140323
rect -79765 -140331 -79721 -140323
rect -79265 -140331 -79221 -140323
rect -79165 -140331 -79121 -140323
rect -79065 -140331 -79021 -140323
rect -78965 -140331 -78921 -140323
rect -78865 -140331 -78821 -140323
rect -78765 -140331 -78721 -140323
rect -78665 -140331 -78621 -140323
rect -78565 -140331 -78521 -140323
rect -78465 -140331 -78421 -140323
rect -78365 -140331 -78321 -140323
rect -78265 -140331 -78221 -140323
rect -78165 -140331 -78121 -140323
rect -78065 -140331 -78021 -140323
rect -77965 -140331 -77921 -140323
rect -77865 -140331 -77821 -140323
rect -77765 -140331 -77721 -140323
rect -77265 -140331 -77221 -140323
rect -77165 -140331 -77121 -140323
rect -77065 -140331 -77021 -140323
rect -76965 -140331 -76921 -140323
rect -76865 -140331 -76821 -140323
rect -76765 -140331 -76721 -140323
rect -76665 -140331 -76621 -140323
rect -76565 -140331 -76521 -140323
rect -76465 -140331 -76421 -140323
rect -76365 -140331 -76321 -140323
rect -76265 -140331 -76221 -140323
rect -76165 -140331 -76121 -140323
rect -76065 -140331 -76021 -140323
rect -75965 -140331 -75921 -140323
rect -75865 -140331 -75821 -140323
rect -75765 -140331 -75721 -140323
rect -83221 -140375 -83213 -140331
rect -83121 -140375 -83113 -140331
rect -83021 -140375 -83013 -140331
rect -82921 -140375 -82913 -140331
rect -82821 -140375 -82813 -140331
rect -82721 -140375 -82713 -140331
rect -82621 -140375 -82613 -140331
rect -82521 -140375 -82513 -140331
rect -82421 -140375 -82413 -140331
rect -82321 -140375 -82313 -140331
rect -82221 -140375 -82213 -140331
rect -82121 -140375 -82113 -140331
rect -82021 -140375 -82013 -140331
rect -81921 -140375 -81913 -140331
rect -81821 -140375 -81813 -140331
rect -81721 -140375 -81713 -140331
rect -81221 -140375 -81213 -140331
rect -81121 -140375 -81113 -140331
rect -81021 -140375 -81013 -140331
rect -80921 -140375 -80913 -140331
rect -80821 -140375 -80813 -140331
rect -80721 -140375 -80713 -140331
rect -80621 -140375 -80613 -140331
rect -80521 -140375 -80513 -140331
rect -80421 -140375 -80413 -140331
rect -80321 -140375 -80313 -140331
rect -80221 -140375 -80213 -140331
rect -80121 -140375 -80113 -140331
rect -80021 -140375 -80013 -140331
rect -79921 -140375 -79913 -140331
rect -79821 -140375 -79813 -140331
rect -79721 -140375 -79713 -140331
rect -79221 -140375 -79213 -140331
rect -79121 -140375 -79113 -140331
rect -79021 -140375 -79013 -140331
rect -78921 -140375 -78913 -140331
rect -78821 -140375 -78813 -140331
rect -78721 -140375 -78713 -140331
rect -78621 -140375 -78613 -140331
rect -78521 -140375 -78513 -140331
rect -78421 -140375 -78413 -140331
rect -78321 -140375 -78313 -140331
rect -78221 -140375 -78213 -140331
rect -78121 -140375 -78113 -140331
rect -78021 -140375 -78013 -140331
rect -77921 -140375 -77913 -140331
rect -77821 -140375 -77813 -140331
rect -77721 -140375 -77713 -140331
rect -77221 -140375 -77213 -140331
rect -77121 -140375 -77113 -140331
rect -77021 -140375 -77013 -140331
rect -76921 -140375 -76913 -140331
rect -76821 -140375 -76813 -140331
rect -76721 -140375 -76713 -140331
rect -76621 -140375 -76613 -140331
rect -76521 -140375 -76513 -140331
rect -76421 -140375 -76413 -140331
rect -76321 -140375 -76313 -140331
rect -76221 -140375 -76213 -140331
rect -76121 -140375 -76113 -140331
rect -76021 -140375 -76013 -140331
rect -75921 -140375 -75913 -140331
rect -75821 -140375 -75813 -140331
rect -75721 -140375 -75713 -140331
rect -83265 -140431 -83221 -140423
rect -83165 -140431 -83121 -140423
rect -83065 -140431 -83021 -140423
rect -82965 -140431 -82921 -140423
rect -82865 -140431 -82821 -140423
rect -82765 -140431 -82721 -140423
rect -82665 -140431 -82621 -140423
rect -82565 -140431 -82521 -140423
rect -82465 -140431 -82421 -140423
rect -82365 -140431 -82321 -140423
rect -82265 -140431 -82221 -140423
rect -82165 -140431 -82121 -140423
rect -82065 -140431 -82021 -140423
rect -81965 -140431 -81921 -140423
rect -81865 -140431 -81821 -140423
rect -81765 -140431 -81721 -140423
rect -81265 -140431 -81221 -140423
rect -81165 -140431 -81121 -140423
rect -81065 -140431 -81021 -140423
rect -80965 -140431 -80921 -140423
rect -80865 -140431 -80821 -140423
rect -80765 -140431 -80721 -140423
rect -80665 -140431 -80621 -140423
rect -80565 -140431 -80521 -140423
rect -80465 -140431 -80421 -140423
rect -80365 -140431 -80321 -140423
rect -80265 -140431 -80221 -140423
rect -80165 -140431 -80121 -140423
rect -80065 -140431 -80021 -140423
rect -79965 -140431 -79921 -140423
rect -79865 -140431 -79821 -140423
rect -79765 -140431 -79721 -140423
rect -79265 -140431 -79221 -140423
rect -79165 -140431 -79121 -140423
rect -79065 -140431 -79021 -140423
rect -78965 -140431 -78921 -140423
rect -78865 -140431 -78821 -140423
rect -78765 -140431 -78721 -140423
rect -78665 -140431 -78621 -140423
rect -78565 -140431 -78521 -140423
rect -78465 -140431 -78421 -140423
rect -78365 -140431 -78321 -140423
rect -78265 -140431 -78221 -140423
rect -78165 -140431 -78121 -140423
rect -78065 -140431 -78021 -140423
rect -77965 -140431 -77921 -140423
rect -77865 -140431 -77821 -140423
rect -77765 -140431 -77721 -140423
rect -77265 -140431 -77221 -140423
rect -77165 -140431 -77121 -140423
rect -77065 -140431 -77021 -140423
rect -76965 -140431 -76921 -140423
rect -76865 -140431 -76821 -140423
rect -76765 -140431 -76721 -140423
rect -76665 -140431 -76621 -140423
rect -76565 -140431 -76521 -140423
rect -76465 -140431 -76421 -140423
rect -76365 -140431 -76321 -140423
rect -76265 -140431 -76221 -140423
rect -76165 -140431 -76121 -140423
rect -76065 -140431 -76021 -140423
rect -75965 -140431 -75921 -140423
rect -75865 -140431 -75821 -140423
rect -75765 -140431 -75721 -140423
rect -83221 -140475 -83213 -140431
rect -83121 -140475 -83113 -140431
rect -83021 -140475 -83013 -140431
rect -82921 -140475 -82913 -140431
rect -82821 -140475 -82813 -140431
rect -82721 -140475 -82713 -140431
rect -82621 -140475 -82613 -140431
rect -82521 -140475 -82513 -140431
rect -82421 -140475 -82413 -140431
rect -82321 -140475 -82313 -140431
rect -82221 -140475 -82213 -140431
rect -82121 -140475 -82113 -140431
rect -82021 -140475 -82013 -140431
rect -81921 -140475 -81913 -140431
rect -81821 -140475 -81813 -140431
rect -81721 -140475 -81713 -140431
rect -81221 -140475 -81213 -140431
rect -81121 -140475 -81113 -140431
rect -81021 -140475 -81013 -140431
rect -80921 -140475 -80913 -140431
rect -80821 -140475 -80813 -140431
rect -80721 -140475 -80713 -140431
rect -80621 -140475 -80613 -140431
rect -80521 -140475 -80513 -140431
rect -80421 -140475 -80413 -140431
rect -80321 -140475 -80313 -140431
rect -80221 -140475 -80213 -140431
rect -80121 -140475 -80113 -140431
rect -80021 -140475 -80013 -140431
rect -79921 -140475 -79913 -140431
rect -79821 -140475 -79813 -140431
rect -79721 -140475 -79713 -140431
rect -79221 -140475 -79213 -140431
rect -79121 -140475 -79113 -140431
rect -79021 -140475 -79013 -140431
rect -78921 -140475 -78913 -140431
rect -78821 -140475 -78813 -140431
rect -78721 -140475 -78713 -140431
rect -78621 -140475 -78613 -140431
rect -78521 -140475 -78513 -140431
rect -78421 -140475 -78413 -140431
rect -78321 -140475 -78313 -140431
rect -78221 -140475 -78213 -140431
rect -78121 -140475 -78113 -140431
rect -78021 -140475 -78013 -140431
rect -77921 -140475 -77913 -140431
rect -77821 -140475 -77813 -140431
rect -77721 -140475 -77713 -140431
rect -77221 -140475 -77213 -140431
rect -77121 -140475 -77113 -140431
rect -77021 -140475 -77013 -140431
rect -76921 -140475 -76913 -140431
rect -76821 -140475 -76813 -140431
rect -76721 -140475 -76713 -140431
rect -76621 -140475 -76613 -140431
rect -76521 -140475 -76513 -140431
rect -76421 -140475 -76413 -140431
rect -76321 -140475 -76313 -140431
rect -76221 -140475 -76213 -140431
rect -76121 -140475 -76113 -140431
rect -76021 -140475 -76013 -140431
rect -75921 -140475 -75913 -140431
rect -75821 -140475 -75813 -140431
rect -75721 -140475 -75713 -140431
rect -83265 -140531 -83221 -140523
rect -83165 -140531 -83121 -140523
rect -83065 -140531 -83021 -140523
rect -82965 -140531 -82921 -140523
rect -82865 -140531 -82821 -140523
rect -82765 -140531 -82721 -140523
rect -82665 -140531 -82621 -140523
rect -82565 -140531 -82521 -140523
rect -82465 -140531 -82421 -140523
rect -82365 -140531 -82321 -140523
rect -82265 -140531 -82221 -140523
rect -82165 -140531 -82121 -140523
rect -82065 -140531 -82021 -140523
rect -81965 -140531 -81921 -140523
rect -81865 -140531 -81821 -140523
rect -81765 -140531 -81721 -140523
rect -81265 -140531 -81221 -140523
rect -81165 -140531 -81121 -140523
rect -81065 -140531 -81021 -140523
rect -80965 -140531 -80921 -140523
rect -80865 -140531 -80821 -140523
rect -80765 -140531 -80721 -140523
rect -80665 -140531 -80621 -140523
rect -80565 -140531 -80521 -140523
rect -80465 -140531 -80421 -140523
rect -80365 -140531 -80321 -140523
rect -80265 -140531 -80221 -140523
rect -80165 -140531 -80121 -140523
rect -80065 -140531 -80021 -140523
rect -79965 -140531 -79921 -140523
rect -79865 -140531 -79821 -140523
rect -79765 -140531 -79721 -140523
rect -79265 -140531 -79221 -140523
rect -79165 -140531 -79121 -140523
rect -79065 -140531 -79021 -140523
rect -78965 -140531 -78921 -140523
rect -78865 -140531 -78821 -140523
rect -78765 -140531 -78721 -140523
rect -78665 -140531 -78621 -140523
rect -78565 -140531 -78521 -140523
rect -78465 -140531 -78421 -140523
rect -78365 -140531 -78321 -140523
rect -78265 -140531 -78221 -140523
rect -78165 -140531 -78121 -140523
rect -78065 -140531 -78021 -140523
rect -77965 -140531 -77921 -140523
rect -77865 -140531 -77821 -140523
rect -77765 -140531 -77721 -140523
rect -77265 -140531 -77221 -140523
rect -77165 -140531 -77121 -140523
rect -77065 -140531 -77021 -140523
rect -76965 -140531 -76921 -140523
rect -76865 -140531 -76821 -140523
rect -76765 -140531 -76721 -140523
rect -76665 -140531 -76621 -140523
rect -76565 -140531 -76521 -140523
rect -76465 -140531 -76421 -140523
rect -76365 -140531 -76321 -140523
rect -76265 -140531 -76221 -140523
rect -76165 -140531 -76121 -140523
rect -76065 -140531 -76021 -140523
rect -75965 -140531 -75921 -140523
rect -75865 -140531 -75821 -140523
rect -75765 -140531 -75721 -140523
rect -83221 -140575 -83213 -140531
rect -83121 -140575 -83113 -140531
rect -83021 -140575 -83013 -140531
rect -82921 -140575 -82913 -140531
rect -82821 -140575 -82813 -140531
rect -82721 -140575 -82713 -140531
rect -82621 -140575 -82613 -140531
rect -82521 -140575 -82513 -140531
rect -82421 -140575 -82413 -140531
rect -82321 -140575 -82313 -140531
rect -82221 -140575 -82213 -140531
rect -82121 -140575 -82113 -140531
rect -82021 -140575 -82013 -140531
rect -81921 -140575 -81913 -140531
rect -81821 -140575 -81813 -140531
rect -81721 -140575 -81713 -140531
rect -81221 -140575 -81213 -140531
rect -81121 -140575 -81113 -140531
rect -81021 -140575 -81013 -140531
rect -80921 -140575 -80913 -140531
rect -80821 -140575 -80813 -140531
rect -80721 -140575 -80713 -140531
rect -80621 -140575 -80613 -140531
rect -80521 -140575 -80513 -140531
rect -80421 -140575 -80413 -140531
rect -80321 -140575 -80313 -140531
rect -80221 -140575 -80213 -140531
rect -80121 -140575 -80113 -140531
rect -80021 -140575 -80013 -140531
rect -79921 -140575 -79913 -140531
rect -79821 -140575 -79813 -140531
rect -79721 -140575 -79713 -140531
rect -79221 -140575 -79213 -140531
rect -79121 -140575 -79113 -140531
rect -79021 -140575 -79013 -140531
rect -78921 -140575 -78913 -140531
rect -78821 -140575 -78813 -140531
rect -78721 -140575 -78713 -140531
rect -78621 -140575 -78613 -140531
rect -78521 -140575 -78513 -140531
rect -78421 -140575 -78413 -140531
rect -78321 -140575 -78313 -140531
rect -78221 -140575 -78213 -140531
rect -78121 -140575 -78113 -140531
rect -78021 -140575 -78013 -140531
rect -77921 -140575 -77913 -140531
rect -77821 -140575 -77813 -140531
rect -77721 -140575 -77713 -140531
rect -77221 -140575 -77213 -140531
rect -77121 -140575 -77113 -140531
rect -77021 -140575 -77013 -140531
rect -76921 -140575 -76913 -140531
rect -76821 -140575 -76813 -140531
rect -76721 -140575 -76713 -140531
rect -76621 -140575 -76613 -140531
rect -76521 -140575 -76513 -140531
rect -76421 -140575 -76413 -140531
rect -76321 -140575 -76313 -140531
rect -76221 -140575 -76213 -140531
rect -76121 -140575 -76113 -140531
rect -76021 -140575 -76013 -140531
rect -75921 -140575 -75913 -140531
rect -75821 -140575 -75813 -140531
rect -75721 -140575 -75713 -140531
rect -83265 -140631 -83221 -140623
rect -83165 -140631 -83121 -140623
rect -83065 -140631 -83021 -140623
rect -82965 -140631 -82921 -140623
rect -82865 -140631 -82821 -140623
rect -82765 -140631 -82721 -140623
rect -82665 -140631 -82621 -140623
rect -82565 -140631 -82521 -140623
rect -82465 -140631 -82421 -140623
rect -82365 -140631 -82321 -140623
rect -82265 -140631 -82221 -140623
rect -82165 -140631 -82121 -140623
rect -82065 -140631 -82021 -140623
rect -81965 -140631 -81921 -140623
rect -81865 -140631 -81821 -140623
rect -81765 -140631 -81721 -140623
rect -81265 -140631 -81221 -140623
rect -81165 -140631 -81121 -140623
rect -81065 -140631 -81021 -140623
rect -80965 -140631 -80921 -140623
rect -80865 -140631 -80821 -140623
rect -80765 -140631 -80721 -140623
rect -80665 -140631 -80621 -140623
rect -80565 -140631 -80521 -140623
rect -80465 -140631 -80421 -140623
rect -80365 -140631 -80321 -140623
rect -80265 -140631 -80221 -140623
rect -80165 -140631 -80121 -140623
rect -80065 -140631 -80021 -140623
rect -79965 -140631 -79921 -140623
rect -79865 -140631 -79821 -140623
rect -79765 -140631 -79721 -140623
rect -79265 -140631 -79221 -140623
rect -79165 -140631 -79121 -140623
rect -79065 -140631 -79021 -140623
rect -78965 -140631 -78921 -140623
rect -78865 -140631 -78821 -140623
rect -78765 -140631 -78721 -140623
rect -78665 -140631 -78621 -140623
rect -78565 -140631 -78521 -140623
rect -78465 -140631 -78421 -140623
rect -78365 -140631 -78321 -140623
rect -78265 -140631 -78221 -140623
rect -78165 -140631 -78121 -140623
rect -78065 -140631 -78021 -140623
rect -77965 -140631 -77921 -140623
rect -77865 -140631 -77821 -140623
rect -77765 -140631 -77721 -140623
rect -77265 -140631 -77221 -140623
rect -77165 -140631 -77121 -140623
rect -77065 -140631 -77021 -140623
rect -76965 -140631 -76921 -140623
rect -76865 -140631 -76821 -140623
rect -76765 -140631 -76721 -140623
rect -76665 -140631 -76621 -140623
rect -76565 -140631 -76521 -140623
rect -76465 -140631 -76421 -140623
rect -76365 -140631 -76321 -140623
rect -76265 -140631 -76221 -140623
rect -76165 -140631 -76121 -140623
rect -76065 -140631 -76021 -140623
rect -75965 -140631 -75921 -140623
rect -75865 -140631 -75821 -140623
rect -75765 -140631 -75721 -140623
rect -83221 -140675 -83213 -140631
rect -83121 -140675 -83113 -140631
rect -83021 -140675 -83013 -140631
rect -82921 -140675 -82913 -140631
rect -82821 -140675 -82813 -140631
rect -82721 -140675 -82713 -140631
rect -82621 -140675 -82613 -140631
rect -82521 -140675 -82513 -140631
rect -82421 -140675 -82413 -140631
rect -82321 -140675 -82313 -140631
rect -82221 -140675 -82213 -140631
rect -82121 -140675 -82113 -140631
rect -82021 -140675 -82013 -140631
rect -81921 -140675 -81913 -140631
rect -81821 -140675 -81813 -140631
rect -81721 -140675 -81713 -140631
rect -81221 -140675 -81213 -140631
rect -81121 -140675 -81113 -140631
rect -81021 -140675 -81013 -140631
rect -80921 -140675 -80913 -140631
rect -80821 -140675 -80813 -140631
rect -80721 -140675 -80713 -140631
rect -80621 -140675 -80613 -140631
rect -80521 -140675 -80513 -140631
rect -80421 -140675 -80413 -140631
rect -80321 -140675 -80313 -140631
rect -80221 -140675 -80213 -140631
rect -80121 -140675 -80113 -140631
rect -80021 -140675 -80013 -140631
rect -79921 -140675 -79913 -140631
rect -79821 -140675 -79813 -140631
rect -79721 -140675 -79713 -140631
rect -79221 -140675 -79213 -140631
rect -79121 -140675 -79113 -140631
rect -79021 -140675 -79013 -140631
rect -78921 -140675 -78913 -140631
rect -78821 -140675 -78813 -140631
rect -78721 -140675 -78713 -140631
rect -78621 -140675 -78613 -140631
rect -78521 -140675 -78513 -140631
rect -78421 -140675 -78413 -140631
rect -78321 -140675 -78313 -140631
rect -78221 -140675 -78213 -140631
rect -78121 -140675 -78113 -140631
rect -78021 -140675 -78013 -140631
rect -77921 -140675 -77913 -140631
rect -77821 -140675 -77813 -140631
rect -77721 -140675 -77713 -140631
rect -77221 -140675 -77213 -140631
rect -77121 -140675 -77113 -140631
rect -77021 -140675 -77013 -140631
rect -76921 -140675 -76913 -140631
rect -76821 -140675 -76813 -140631
rect -76721 -140675 -76713 -140631
rect -76621 -140675 -76613 -140631
rect -76521 -140675 -76513 -140631
rect -76421 -140675 -76413 -140631
rect -76321 -140675 -76313 -140631
rect -76221 -140675 -76213 -140631
rect -76121 -140675 -76113 -140631
rect -76021 -140675 -76013 -140631
rect -75921 -140675 -75913 -140631
rect -75821 -140675 -75813 -140631
rect -75721 -140675 -75713 -140631
rect -83265 -140731 -83221 -140723
rect -83165 -140731 -83121 -140723
rect -83065 -140731 -83021 -140723
rect -82965 -140731 -82921 -140723
rect -82865 -140731 -82821 -140723
rect -82765 -140731 -82721 -140723
rect -82665 -140731 -82621 -140723
rect -82565 -140731 -82521 -140723
rect -82465 -140731 -82421 -140723
rect -82365 -140731 -82321 -140723
rect -82265 -140731 -82221 -140723
rect -82165 -140731 -82121 -140723
rect -82065 -140731 -82021 -140723
rect -81965 -140731 -81921 -140723
rect -81865 -140731 -81821 -140723
rect -81765 -140731 -81721 -140723
rect -81265 -140731 -81221 -140723
rect -81165 -140731 -81121 -140723
rect -81065 -140731 -81021 -140723
rect -80965 -140731 -80921 -140723
rect -80865 -140731 -80821 -140723
rect -80765 -140731 -80721 -140723
rect -80665 -140731 -80621 -140723
rect -80565 -140731 -80521 -140723
rect -80465 -140731 -80421 -140723
rect -80365 -140731 -80321 -140723
rect -80265 -140731 -80221 -140723
rect -80165 -140731 -80121 -140723
rect -80065 -140731 -80021 -140723
rect -79965 -140731 -79921 -140723
rect -79865 -140731 -79821 -140723
rect -79765 -140731 -79721 -140723
rect -79265 -140731 -79221 -140723
rect -79165 -140731 -79121 -140723
rect -79065 -140731 -79021 -140723
rect -78965 -140731 -78921 -140723
rect -78865 -140731 -78821 -140723
rect -78765 -140731 -78721 -140723
rect -78665 -140731 -78621 -140723
rect -78565 -140731 -78521 -140723
rect -78465 -140731 -78421 -140723
rect -78365 -140731 -78321 -140723
rect -78265 -140731 -78221 -140723
rect -78165 -140731 -78121 -140723
rect -78065 -140731 -78021 -140723
rect -77965 -140731 -77921 -140723
rect -77865 -140731 -77821 -140723
rect -77765 -140731 -77721 -140723
rect -77265 -140731 -77221 -140723
rect -77165 -140731 -77121 -140723
rect -77065 -140731 -77021 -140723
rect -76965 -140731 -76921 -140723
rect -76865 -140731 -76821 -140723
rect -76765 -140731 -76721 -140723
rect -76665 -140731 -76621 -140723
rect -76565 -140731 -76521 -140723
rect -76465 -140731 -76421 -140723
rect -76365 -140731 -76321 -140723
rect -76265 -140731 -76221 -140723
rect -76165 -140731 -76121 -140723
rect -76065 -140731 -76021 -140723
rect -75965 -140731 -75921 -140723
rect -75865 -140731 -75821 -140723
rect -75765 -140731 -75721 -140723
rect -83221 -140775 -83213 -140731
rect -83121 -140775 -83113 -140731
rect -83021 -140775 -83013 -140731
rect -82921 -140775 -82913 -140731
rect -82821 -140775 -82813 -140731
rect -82721 -140775 -82713 -140731
rect -82621 -140775 -82613 -140731
rect -82521 -140775 -82513 -140731
rect -82421 -140775 -82413 -140731
rect -82321 -140775 -82313 -140731
rect -82221 -140775 -82213 -140731
rect -82121 -140775 -82113 -140731
rect -82021 -140775 -82013 -140731
rect -81921 -140775 -81913 -140731
rect -81821 -140775 -81813 -140731
rect -81721 -140775 -81713 -140731
rect -81221 -140775 -81213 -140731
rect -81121 -140775 -81113 -140731
rect -81021 -140775 -81013 -140731
rect -80921 -140775 -80913 -140731
rect -80821 -140775 -80813 -140731
rect -80721 -140775 -80713 -140731
rect -80621 -140775 -80613 -140731
rect -80521 -140775 -80513 -140731
rect -80421 -140775 -80413 -140731
rect -80321 -140775 -80313 -140731
rect -80221 -140775 -80213 -140731
rect -80121 -140775 -80113 -140731
rect -80021 -140775 -80013 -140731
rect -79921 -140775 -79913 -140731
rect -79821 -140775 -79813 -140731
rect -79721 -140775 -79713 -140731
rect -79221 -140775 -79213 -140731
rect -79121 -140775 -79113 -140731
rect -79021 -140775 -79013 -140731
rect -78921 -140775 -78913 -140731
rect -78821 -140775 -78813 -140731
rect -78721 -140775 -78713 -140731
rect -78621 -140775 -78613 -140731
rect -78521 -140775 -78513 -140731
rect -78421 -140775 -78413 -140731
rect -78321 -140775 -78313 -140731
rect -78221 -140775 -78213 -140731
rect -78121 -140775 -78113 -140731
rect -78021 -140775 -78013 -140731
rect -77921 -140775 -77913 -140731
rect -77821 -140775 -77813 -140731
rect -77721 -140775 -77713 -140731
rect -77221 -140775 -77213 -140731
rect -77121 -140775 -77113 -140731
rect -77021 -140775 -77013 -140731
rect -76921 -140775 -76913 -140731
rect -76821 -140775 -76813 -140731
rect -76721 -140775 -76713 -140731
rect -76621 -140775 -76613 -140731
rect -76521 -140775 -76513 -140731
rect -76421 -140775 -76413 -140731
rect -76321 -140775 -76313 -140731
rect -76221 -140775 -76213 -140731
rect -76121 -140775 -76113 -140731
rect -76021 -140775 -76013 -140731
rect -75921 -140775 -75913 -140731
rect -75821 -140775 -75813 -140731
rect -75721 -140775 -75713 -140731
rect -83265 -140831 -83221 -140823
rect -83165 -140831 -83121 -140823
rect -83065 -140831 -83021 -140823
rect -82965 -140831 -82921 -140823
rect -82865 -140831 -82821 -140823
rect -82765 -140831 -82721 -140823
rect -82665 -140831 -82621 -140823
rect -82565 -140831 -82521 -140823
rect -82465 -140831 -82421 -140823
rect -82365 -140831 -82321 -140823
rect -82265 -140831 -82221 -140823
rect -82165 -140831 -82121 -140823
rect -82065 -140831 -82021 -140823
rect -81965 -140831 -81921 -140823
rect -81865 -140831 -81821 -140823
rect -81765 -140831 -81721 -140823
rect -81265 -140831 -81221 -140823
rect -81165 -140831 -81121 -140823
rect -81065 -140831 -81021 -140823
rect -80965 -140831 -80921 -140823
rect -80865 -140831 -80821 -140823
rect -80765 -140831 -80721 -140823
rect -80665 -140831 -80621 -140823
rect -80565 -140831 -80521 -140823
rect -80465 -140831 -80421 -140823
rect -80365 -140831 -80321 -140823
rect -80265 -140831 -80221 -140823
rect -80165 -140831 -80121 -140823
rect -80065 -140831 -80021 -140823
rect -79965 -140831 -79921 -140823
rect -79865 -140831 -79821 -140823
rect -79765 -140831 -79721 -140823
rect -79265 -140831 -79221 -140823
rect -79165 -140831 -79121 -140823
rect -79065 -140831 -79021 -140823
rect -78965 -140831 -78921 -140823
rect -78865 -140831 -78821 -140823
rect -78765 -140831 -78721 -140823
rect -78665 -140831 -78621 -140823
rect -78565 -140831 -78521 -140823
rect -78465 -140831 -78421 -140823
rect -78365 -140831 -78321 -140823
rect -78265 -140831 -78221 -140823
rect -78165 -140831 -78121 -140823
rect -78065 -140831 -78021 -140823
rect -77965 -140831 -77921 -140823
rect -77865 -140831 -77821 -140823
rect -77765 -140831 -77721 -140823
rect -77265 -140831 -77221 -140823
rect -77165 -140831 -77121 -140823
rect -77065 -140831 -77021 -140823
rect -76965 -140831 -76921 -140823
rect -76865 -140831 -76821 -140823
rect -76765 -140831 -76721 -140823
rect -76665 -140831 -76621 -140823
rect -76565 -140831 -76521 -140823
rect -76465 -140831 -76421 -140823
rect -76365 -140831 -76321 -140823
rect -76265 -140831 -76221 -140823
rect -76165 -140831 -76121 -140823
rect -76065 -140831 -76021 -140823
rect -75965 -140831 -75921 -140823
rect -75865 -140831 -75821 -140823
rect -75765 -140831 -75721 -140823
rect -83221 -140875 -83213 -140831
rect -83121 -140875 -83113 -140831
rect -83021 -140875 -83013 -140831
rect -82921 -140875 -82913 -140831
rect -82821 -140875 -82813 -140831
rect -82721 -140875 -82713 -140831
rect -82621 -140875 -82613 -140831
rect -82521 -140875 -82513 -140831
rect -82421 -140875 -82413 -140831
rect -82321 -140875 -82313 -140831
rect -82221 -140875 -82213 -140831
rect -82121 -140875 -82113 -140831
rect -82021 -140875 -82013 -140831
rect -81921 -140875 -81913 -140831
rect -81821 -140875 -81813 -140831
rect -81721 -140875 -81713 -140831
rect -81221 -140875 -81213 -140831
rect -81121 -140875 -81113 -140831
rect -81021 -140875 -81013 -140831
rect -80921 -140875 -80913 -140831
rect -80821 -140875 -80813 -140831
rect -80721 -140875 -80713 -140831
rect -80621 -140875 -80613 -140831
rect -80521 -140875 -80513 -140831
rect -80421 -140875 -80413 -140831
rect -80321 -140875 -80313 -140831
rect -80221 -140875 -80213 -140831
rect -80121 -140875 -80113 -140831
rect -80021 -140875 -80013 -140831
rect -79921 -140875 -79913 -140831
rect -79821 -140875 -79813 -140831
rect -79721 -140875 -79713 -140831
rect -79221 -140875 -79213 -140831
rect -79121 -140875 -79113 -140831
rect -79021 -140875 -79013 -140831
rect -78921 -140875 -78913 -140831
rect -78821 -140875 -78813 -140831
rect -78721 -140875 -78713 -140831
rect -78621 -140875 -78613 -140831
rect -78521 -140875 -78513 -140831
rect -78421 -140875 -78413 -140831
rect -78321 -140875 -78313 -140831
rect -78221 -140875 -78213 -140831
rect -78121 -140875 -78113 -140831
rect -78021 -140875 -78013 -140831
rect -77921 -140875 -77913 -140831
rect -77821 -140875 -77813 -140831
rect -77721 -140875 -77713 -140831
rect -77221 -140875 -77213 -140831
rect -77121 -140875 -77113 -140831
rect -77021 -140875 -77013 -140831
rect -76921 -140875 -76913 -140831
rect -76821 -140875 -76813 -140831
rect -76721 -140875 -76713 -140831
rect -76621 -140875 -76613 -140831
rect -76521 -140875 -76513 -140831
rect -76421 -140875 -76413 -140831
rect -76321 -140875 -76313 -140831
rect -76221 -140875 -76213 -140831
rect -76121 -140875 -76113 -140831
rect -76021 -140875 -76013 -140831
rect -75921 -140875 -75913 -140831
rect -75821 -140875 -75813 -140831
rect -75721 -140875 -75713 -140831
rect -83265 -140931 -83221 -140923
rect -83165 -140931 -83121 -140923
rect -83065 -140931 -83021 -140923
rect -82965 -140931 -82921 -140923
rect -82865 -140931 -82821 -140923
rect -82765 -140931 -82721 -140923
rect -82665 -140931 -82621 -140923
rect -82565 -140931 -82521 -140923
rect -82465 -140931 -82421 -140923
rect -82365 -140931 -82321 -140923
rect -82265 -140931 -82221 -140923
rect -82165 -140931 -82121 -140923
rect -82065 -140931 -82021 -140923
rect -81965 -140931 -81921 -140923
rect -81865 -140931 -81821 -140923
rect -81765 -140931 -81721 -140923
rect -81265 -140931 -81221 -140923
rect -81165 -140931 -81121 -140923
rect -81065 -140931 -81021 -140923
rect -80965 -140931 -80921 -140923
rect -80865 -140931 -80821 -140923
rect -80765 -140931 -80721 -140923
rect -80665 -140931 -80621 -140923
rect -80565 -140931 -80521 -140923
rect -80465 -140931 -80421 -140923
rect -80365 -140931 -80321 -140923
rect -80265 -140931 -80221 -140923
rect -80165 -140931 -80121 -140923
rect -80065 -140931 -80021 -140923
rect -79965 -140931 -79921 -140923
rect -79865 -140931 -79821 -140923
rect -79765 -140931 -79721 -140923
rect -79265 -140931 -79221 -140923
rect -79165 -140931 -79121 -140923
rect -79065 -140931 -79021 -140923
rect -78965 -140931 -78921 -140923
rect -78865 -140931 -78821 -140923
rect -78765 -140931 -78721 -140923
rect -78665 -140931 -78621 -140923
rect -78565 -140931 -78521 -140923
rect -78465 -140931 -78421 -140923
rect -78365 -140931 -78321 -140923
rect -78265 -140931 -78221 -140923
rect -78165 -140931 -78121 -140923
rect -78065 -140931 -78021 -140923
rect -77965 -140931 -77921 -140923
rect -77865 -140931 -77821 -140923
rect -77765 -140931 -77721 -140923
rect -77265 -140931 -77221 -140923
rect -77165 -140931 -77121 -140923
rect -77065 -140931 -77021 -140923
rect -76965 -140931 -76921 -140923
rect -76865 -140931 -76821 -140923
rect -76765 -140931 -76721 -140923
rect -76665 -140931 -76621 -140923
rect -76565 -140931 -76521 -140923
rect -76465 -140931 -76421 -140923
rect -76365 -140931 -76321 -140923
rect -76265 -140931 -76221 -140923
rect -76165 -140931 -76121 -140923
rect -76065 -140931 -76021 -140923
rect -75965 -140931 -75921 -140923
rect -75865 -140931 -75821 -140923
rect -75765 -140931 -75721 -140923
rect -83221 -140975 -83213 -140931
rect -83121 -140975 -83113 -140931
rect -83021 -140975 -83013 -140931
rect -82921 -140975 -82913 -140931
rect -82821 -140975 -82813 -140931
rect -82721 -140975 -82713 -140931
rect -82621 -140975 -82613 -140931
rect -82521 -140975 -82513 -140931
rect -82421 -140975 -82413 -140931
rect -82321 -140975 -82313 -140931
rect -82221 -140975 -82213 -140931
rect -82121 -140975 -82113 -140931
rect -82021 -140975 -82013 -140931
rect -81921 -140975 -81913 -140931
rect -81821 -140975 -81813 -140931
rect -81721 -140975 -81713 -140931
rect -81221 -140975 -81213 -140931
rect -81121 -140975 -81113 -140931
rect -81021 -140975 -81013 -140931
rect -80921 -140975 -80913 -140931
rect -80821 -140975 -80813 -140931
rect -80721 -140975 -80713 -140931
rect -80621 -140975 -80613 -140931
rect -80521 -140975 -80513 -140931
rect -80421 -140975 -80413 -140931
rect -80321 -140975 -80313 -140931
rect -80221 -140975 -80213 -140931
rect -80121 -140975 -80113 -140931
rect -80021 -140975 -80013 -140931
rect -79921 -140975 -79913 -140931
rect -79821 -140975 -79813 -140931
rect -79721 -140975 -79713 -140931
rect -79221 -140975 -79213 -140931
rect -79121 -140975 -79113 -140931
rect -79021 -140975 -79013 -140931
rect -78921 -140975 -78913 -140931
rect -78821 -140975 -78813 -140931
rect -78721 -140975 -78713 -140931
rect -78621 -140975 -78613 -140931
rect -78521 -140975 -78513 -140931
rect -78421 -140975 -78413 -140931
rect -78321 -140975 -78313 -140931
rect -78221 -140975 -78213 -140931
rect -78121 -140975 -78113 -140931
rect -78021 -140975 -78013 -140931
rect -77921 -140975 -77913 -140931
rect -77821 -140975 -77813 -140931
rect -77721 -140975 -77713 -140931
rect -77221 -140975 -77213 -140931
rect -77121 -140975 -77113 -140931
rect -77021 -140975 -77013 -140931
rect -76921 -140975 -76913 -140931
rect -76821 -140975 -76813 -140931
rect -76721 -140975 -76713 -140931
rect -76621 -140975 -76613 -140931
rect -76521 -140975 -76513 -140931
rect -76421 -140975 -76413 -140931
rect -76321 -140975 -76313 -140931
rect -76221 -140975 -76213 -140931
rect -76121 -140975 -76113 -140931
rect -76021 -140975 -76013 -140931
rect -75921 -140975 -75913 -140931
rect -75821 -140975 -75813 -140931
rect -75721 -140975 -75713 -140931
rect -83265 -141031 -83221 -141023
rect -83165 -141031 -83121 -141023
rect -83065 -141031 -83021 -141023
rect -82965 -141031 -82921 -141023
rect -82865 -141031 -82821 -141023
rect -82765 -141031 -82721 -141023
rect -82665 -141031 -82621 -141023
rect -82565 -141031 -82521 -141023
rect -82465 -141031 -82421 -141023
rect -82365 -141031 -82321 -141023
rect -82265 -141031 -82221 -141023
rect -82165 -141031 -82121 -141023
rect -82065 -141031 -82021 -141023
rect -81965 -141031 -81921 -141023
rect -81865 -141031 -81821 -141023
rect -81765 -141031 -81721 -141023
rect -81265 -141031 -81221 -141023
rect -81165 -141031 -81121 -141023
rect -81065 -141031 -81021 -141023
rect -80965 -141031 -80921 -141023
rect -80865 -141031 -80821 -141023
rect -80765 -141031 -80721 -141023
rect -80665 -141031 -80621 -141023
rect -80565 -141031 -80521 -141023
rect -80465 -141031 -80421 -141023
rect -80365 -141031 -80321 -141023
rect -80265 -141031 -80221 -141023
rect -80165 -141031 -80121 -141023
rect -80065 -141031 -80021 -141023
rect -79965 -141031 -79921 -141023
rect -79865 -141031 -79821 -141023
rect -79765 -141031 -79721 -141023
rect -79265 -141031 -79221 -141023
rect -79165 -141031 -79121 -141023
rect -79065 -141031 -79021 -141023
rect -78965 -141031 -78921 -141023
rect -78865 -141031 -78821 -141023
rect -78765 -141031 -78721 -141023
rect -78665 -141031 -78621 -141023
rect -78565 -141031 -78521 -141023
rect -78465 -141031 -78421 -141023
rect -78365 -141031 -78321 -141023
rect -78265 -141031 -78221 -141023
rect -78165 -141031 -78121 -141023
rect -78065 -141031 -78021 -141023
rect -77965 -141031 -77921 -141023
rect -77865 -141031 -77821 -141023
rect -77765 -141031 -77721 -141023
rect -77265 -141031 -77221 -141023
rect -77165 -141031 -77121 -141023
rect -77065 -141031 -77021 -141023
rect -76965 -141031 -76921 -141023
rect -76865 -141031 -76821 -141023
rect -76765 -141031 -76721 -141023
rect -76665 -141031 -76621 -141023
rect -76565 -141031 -76521 -141023
rect -76465 -141031 -76421 -141023
rect -76365 -141031 -76321 -141023
rect -76265 -141031 -76221 -141023
rect -76165 -141031 -76121 -141023
rect -76065 -141031 -76021 -141023
rect -75965 -141031 -75921 -141023
rect -75865 -141031 -75821 -141023
rect -75765 -141031 -75721 -141023
rect -83221 -141075 -83213 -141031
rect -83121 -141075 -83113 -141031
rect -83021 -141075 -83013 -141031
rect -82921 -141075 -82913 -141031
rect -82821 -141075 -82813 -141031
rect -82721 -141075 -82713 -141031
rect -82621 -141075 -82613 -141031
rect -82521 -141075 -82513 -141031
rect -82421 -141075 -82413 -141031
rect -82321 -141075 -82313 -141031
rect -82221 -141075 -82213 -141031
rect -82121 -141075 -82113 -141031
rect -82021 -141075 -82013 -141031
rect -81921 -141075 -81913 -141031
rect -81821 -141075 -81813 -141031
rect -81721 -141075 -81713 -141031
rect -81221 -141075 -81213 -141031
rect -81121 -141075 -81113 -141031
rect -81021 -141075 -81013 -141031
rect -80921 -141075 -80913 -141031
rect -80821 -141075 -80813 -141031
rect -80721 -141075 -80713 -141031
rect -80621 -141075 -80613 -141031
rect -80521 -141075 -80513 -141031
rect -80421 -141075 -80413 -141031
rect -80321 -141075 -80313 -141031
rect -80221 -141075 -80213 -141031
rect -80121 -141075 -80113 -141031
rect -80021 -141075 -80013 -141031
rect -79921 -141075 -79913 -141031
rect -79821 -141075 -79813 -141031
rect -79721 -141075 -79713 -141031
rect -79221 -141075 -79213 -141031
rect -79121 -141075 -79113 -141031
rect -79021 -141075 -79013 -141031
rect -78921 -141075 -78913 -141031
rect -78821 -141075 -78813 -141031
rect -78721 -141075 -78713 -141031
rect -78621 -141075 -78613 -141031
rect -78521 -141075 -78513 -141031
rect -78421 -141075 -78413 -141031
rect -78321 -141075 -78313 -141031
rect -78221 -141075 -78213 -141031
rect -78121 -141075 -78113 -141031
rect -78021 -141075 -78013 -141031
rect -77921 -141075 -77913 -141031
rect -77821 -141075 -77813 -141031
rect -77721 -141075 -77713 -141031
rect -77221 -141075 -77213 -141031
rect -77121 -141075 -77113 -141031
rect -77021 -141075 -77013 -141031
rect -76921 -141075 -76913 -141031
rect -76821 -141075 -76813 -141031
rect -76721 -141075 -76713 -141031
rect -76621 -141075 -76613 -141031
rect -76521 -141075 -76513 -141031
rect -76421 -141075 -76413 -141031
rect -76321 -141075 -76313 -141031
rect -76221 -141075 -76213 -141031
rect -76121 -141075 -76113 -141031
rect -76021 -141075 -76013 -141031
rect -75921 -141075 -75913 -141031
rect -75821 -141075 -75813 -141031
rect -75721 -141075 -75713 -141031
rect -83265 -141131 -83221 -141123
rect -83165 -141131 -83121 -141123
rect -83065 -141131 -83021 -141123
rect -82965 -141131 -82921 -141123
rect -82865 -141131 -82821 -141123
rect -82765 -141131 -82721 -141123
rect -82665 -141131 -82621 -141123
rect -82565 -141131 -82521 -141123
rect -82465 -141131 -82421 -141123
rect -82365 -141131 -82321 -141123
rect -82265 -141131 -82221 -141123
rect -82165 -141131 -82121 -141123
rect -82065 -141131 -82021 -141123
rect -81965 -141131 -81921 -141123
rect -81865 -141131 -81821 -141123
rect -81765 -141131 -81721 -141123
rect -81265 -141131 -81221 -141123
rect -81165 -141131 -81121 -141123
rect -81065 -141131 -81021 -141123
rect -80965 -141131 -80921 -141123
rect -80865 -141131 -80821 -141123
rect -80765 -141131 -80721 -141123
rect -80665 -141131 -80621 -141123
rect -80565 -141131 -80521 -141123
rect -80465 -141131 -80421 -141123
rect -80365 -141131 -80321 -141123
rect -80265 -141131 -80221 -141123
rect -80165 -141131 -80121 -141123
rect -80065 -141131 -80021 -141123
rect -79965 -141131 -79921 -141123
rect -79865 -141131 -79821 -141123
rect -79765 -141131 -79721 -141123
rect -79265 -141131 -79221 -141123
rect -79165 -141131 -79121 -141123
rect -79065 -141131 -79021 -141123
rect -78965 -141131 -78921 -141123
rect -78865 -141131 -78821 -141123
rect -78765 -141131 -78721 -141123
rect -78665 -141131 -78621 -141123
rect -78565 -141131 -78521 -141123
rect -78465 -141131 -78421 -141123
rect -78365 -141131 -78321 -141123
rect -78265 -141131 -78221 -141123
rect -78165 -141131 -78121 -141123
rect -78065 -141131 -78021 -141123
rect -77965 -141131 -77921 -141123
rect -77865 -141131 -77821 -141123
rect -77765 -141131 -77721 -141123
rect -77265 -141131 -77221 -141123
rect -77165 -141131 -77121 -141123
rect -77065 -141131 -77021 -141123
rect -76965 -141131 -76921 -141123
rect -76865 -141131 -76821 -141123
rect -76765 -141131 -76721 -141123
rect -76665 -141131 -76621 -141123
rect -76565 -141131 -76521 -141123
rect -76465 -141131 -76421 -141123
rect -76365 -141131 -76321 -141123
rect -76265 -141131 -76221 -141123
rect -76165 -141131 -76121 -141123
rect -76065 -141131 -76021 -141123
rect -75965 -141131 -75921 -141123
rect -75865 -141131 -75821 -141123
rect -75765 -141131 -75721 -141123
rect -83221 -141175 -83213 -141131
rect -83121 -141175 -83113 -141131
rect -83021 -141175 -83013 -141131
rect -82921 -141175 -82913 -141131
rect -82821 -141175 -82813 -141131
rect -82721 -141175 -82713 -141131
rect -82621 -141175 -82613 -141131
rect -82521 -141175 -82513 -141131
rect -82421 -141175 -82413 -141131
rect -82321 -141175 -82313 -141131
rect -82221 -141175 -82213 -141131
rect -82121 -141175 -82113 -141131
rect -82021 -141175 -82013 -141131
rect -81921 -141175 -81913 -141131
rect -81821 -141175 -81813 -141131
rect -81721 -141175 -81713 -141131
rect -81221 -141175 -81213 -141131
rect -81121 -141175 -81113 -141131
rect -81021 -141175 -81013 -141131
rect -80921 -141175 -80913 -141131
rect -80821 -141175 -80813 -141131
rect -80721 -141175 -80713 -141131
rect -80621 -141175 -80613 -141131
rect -80521 -141175 -80513 -141131
rect -80421 -141175 -80413 -141131
rect -80321 -141175 -80313 -141131
rect -80221 -141175 -80213 -141131
rect -80121 -141175 -80113 -141131
rect -80021 -141175 -80013 -141131
rect -79921 -141175 -79913 -141131
rect -79821 -141175 -79813 -141131
rect -79721 -141175 -79713 -141131
rect -79221 -141175 -79213 -141131
rect -79121 -141175 -79113 -141131
rect -79021 -141175 -79013 -141131
rect -78921 -141175 -78913 -141131
rect -78821 -141175 -78813 -141131
rect -78721 -141175 -78713 -141131
rect -78621 -141175 -78613 -141131
rect -78521 -141175 -78513 -141131
rect -78421 -141175 -78413 -141131
rect -78321 -141175 -78313 -141131
rect -78221 -141175 -78213 -141131
rect -78121 -141175 -78113 -141131
rect -78021 -141175 -78013 -141131
rect -77921 -141175 -77913 -141131
rect -77821 -141175 -77813 -141131
rect -77721 -141175 -77713 -141131
rect -77221 -141175 -77213 -141131
rect -77121 -141175 -77113 -141131
rect -77021 -141175 -77013 -141131
rect -76921 -141175 -76913 -141131
rect -76821 -141175 -76813 -141131
rect -76721 -141175 -76713 -141131
rect -76621 -141175 -76613 -141131
rect -76521 -141175 -76513 -141131
rect -76421 -141175 -76413 -141131
rect -76321 -141175 -76313 -141131
rect -76221 -141175 -76213 -141131
rect -76121 -141175 -76113 -141131
rect -76021 -141175 -76013 -141131
rect -75921 -141175 -75913 -141131
rect -75821 -141175 -75813 -141131
rect -75721 -141175 -75713 -141131
rect -83265 -141231 -83221 -141223
rect -83165 -141231 -83121 -141223
rect -83065 -141231 -83021 -141223
rect -82965 -141231 -82921 -141223
rect -82865 -141231 -82821 -141223
rect -82765 -141231 -82721 -141223
rect -82665 -141231 -82621 -141223
rect -82565 -141231 -82521 -141223
rect -82465 -141231 -82421 -141223
rect -82365 -141231 -82321 -141223
rect -82265 -141231 -82221 -141223
rect -82165 -141231 -82121 -141223
rect -82065 -141231 -82021 -141223
rect -81965 -141231 -81921 -141223
rect -81865 -141231 -81821 -141223
rect -81765 -141231 -81721 -141223
rect -81265 -141231 -81221 -141223
rect -81165 -141231 -81121 -141223
rect -81065 -141231 -81021 -141223
rect -80965 -141231 -80921 -141223
rect -80865 -141231 -80821 -141223
rect -80765 -141231 -80721 -141223
rect -80665 -141231 -80621 -141223
rect -80565 -141231 -80521 -141223
rect -80465 -141231 -80421 -141223
rect -80365 -141231 -80321 -141223
rect -80265 -141231 -80221 -141223
rect -80165 -141231 -80121 -141223
rect -80065 -141231 -80021 -141223
rect -79965 -141231 -79921 -141223
rect -79865 -141231 -79821 -141223
rect -79765 -141231 -79721 -141223
rect -79265 -141231 -79221 -141223
rect -79165 -141231 -79121 -141223
rect -79065 -141231 -79021 -141223
rect -78965 -141231 -78921 -141223
rect -78865 -141231 -78821 -141223
rect -78765 -141231 -78721 -141223
rect -78665 -141231 -78621 -141223
rect -78565 -141231 -78521 -141223
rect -78465 -141231 -78421 -141223
rect -78365 -141231 -78321 -141223
rect -78265 -141231 -78221 -141223
rect -78165 -141231 -78121 -141223
rect -78065 -141231 -78021 -141223
rect -77965 -141231 -77921 -141223
rect -77865 -141231 -77821 -141223
rect -77765 -141231 -77721 -141223
rect -77265 -141231 -77221 -141223
rect -77165 -141231 -77121 -141223
rect -77065 -141231 -77021 -141223
rect -76965 -141231 -76921 -141223
rect -76865 -141231 -76821 -141223
rect -76765 -141231 -76721 -141223
rect -76665 -141231 -76621 -141223
rect -76565 -141231 -76521 -141223
rect -76465 -141231 -76421 -141223
rect -76365 -141231 -76321 -141223
rect -76265 -141231 -76221 -141223
rect -76165 -141231 -76121 -141223
rect -76065 -141231 -76021 -141223
rect -75965 -141231 -75921 -141223
rect -75865 -141231 -75821 -141223
rect -75765 -141231 -75721 -141223
rect -83221 -141275 -83213 -141231
rect -83121 -141275 -83113 -141231
rect -83021 -141275 -83013 -141231
rect -82921 -141275 -82913 -141231
rect -82821 -141275 -82813 -141231
rect -82721 -141275 -82713 -141231
rect -82621 -141275 -82613 -141231
rect -82521 -141275 -82513 -141231
rect -82421 -141275 -82413 -141231
rect -82321 -141275 -82313 -141231
rect -82221 -141275 -82213 -141231
rect -82121 -141275 -82113 -141231
rect -82021 -141275 -82013 -141231
rect -81921 -141275 -81913 -141231
rect -81821 -141275 -81813 -141231
rect -81721 -141275 -81713 -141231
rect -81221 -141275 -81213 -141231
rect -81121 -141275 -81113 -141231
rect -81021 -141275 -81013 -141231
rect -80921 -141275 -80913 -141231
rect -80821 -141275 -80813 -141231
rect -80721 -141275 -80713 -141231
rect -80621 -141275 -80613 -141231
rect -80521 -141275 -80513 -141231
rect -80421 -141275 -80413 -141231
rect -80321 -141275 -80313 -141231
rect -80221 -141275 -80213 -141231
rect -80121 -141275 -80113 -141231
rect -80021 -141275 -80013 -141231
rect -79921 -141275 -79913 -141231
rect -79821 -141275 -79813 -141231
rect -79721 -141275 -79713 -141231
rect -79221 -141275 -79213 -141231
rect -79121 -141275 -79113 -141231
rect -79021 -141275 -79013 -141231
rect -78921 -141275 -78913 -141231
rect -78821 -141275 -78813 -141231
rect -78721 -141275 -78713 -141231
rect -78621 -141275 -78613 -141231
rect -78521 -141275 -78513 -141231
rect -78421 -141275 -78413 -141231
rect -78321 -141275 -78313 -141231
rect -78221 -141275 -78213 -141231
rect -78121 -141275 -78113 -141231
rect -78021 -141275 -78013 -141231
rect -77921 -141275 -77913 -141231
rect -77821 -141275 -77813 -141231
rect -77721 -141275 -77713 -141231
rect -77221 -141275 -77213 -141231
rect -77121 -141275 -77113 -141231
rect -77021 -141275 -77013 -141231
rect -76921 -141275 -76913 -141231
rect -76821 -141275 -76813 -141231
rect -76721 -141275 -76713 -141231
rect -76621 -141275 -76613 -141231
rect -76521 -141275 -76513 -141231
rect -76421 -141275 -76413 -141231
rect -76321 -141275 -76313 -141231
rect -76221 -141275 -76213 -141231
rect -76121 -141275 -76113 -141231
rect -76021 -141275 -76013 -141231
rect -75921 -141275 -75913 -141231
rect -75821 -141275 -75813 -141231
rect -75721 -141275 -75713 -141231
rect -83265 -141331 -83221 -141323
rect -83165 -141331 -83121 -141323
rect -83065 -141331 -83021 -141323
rect -82965 -141331 -82921 -141323
rect -82865 -141331 -82821 -141323
rect -82765 -141331 -82721 -141323
rect -82665 -141331 -82621 -141323
rect -82565 -141331 -82521 -141323
rect -82465 -141331 -82421 -141323
rect -82365 -141331 -82321 -141323
rect -82265 -141331 -82221 -141323
rect -82165 -141331 -82121 -141323
rect -82065 -141331 -82021 -141323
rect -81965 -141331 -81921 -141323
rect -81865 -141331 -81821 -141323
rect -81765 -141331 -81721 -141323
rect -81265 -141331 -81221 -141323
rect -81165 -141331 -81121 -141323
rect -81065 -141331 -81021 -141323
rect -80965 -141331 -80921 -141323
rect -80865 -141331 -80821 -141323
rect -80765 -141331 -80721 -141323
rect -80665 -141331 -80621 -141323
rect -80565 -141331 -80521 -141323
rect -80465 -141331 -80421 -141323
rect -80365 -141331 -80321 -141323
rect -80265 -141331 -80221 -141323
rect -80165 -141331 -80121 -141323
rect -80065 -141331 -80021 -141323
rect -79965 -141331 -79921 -141323
rect -79865 -141331 -79821 -141323
rect -79765 -141331 -79721 -141323
rect -79265 -141331 -79221 -141323
rect -79165 -141331 -79121 -141323
rect -79065 -141331 -79021 -141323
rect -78965 -141331 -78921 -141323
rect -78865 -141331 -78821 -141323
rect -78765 -141331 -78721 -141323
rect -78665 -141331 -78621 -141323
rect -78565 -141331 -78521 -141323
rect -78465 -141331 -78421 -141323
rect -78365 -141331 -78321 -141323
rect -78265 -141331 -78221 -141323
rect -78165 -141331 -78121 -141323
rect -78065 -141331 -78021 -141323
rect -77965 -141331 -77921 -141323
rect -77865 -141331 -77821 -141323
rect -77765 -141331 -77721 -141323
rect -77265 -141331 -77221 -141323
rect -77165 -141331 -77121 -141323
rect -77065 -141331 -77021 -141323
rect -76965 -141331 -76921 -141323
rect -76865 -141331 -76821 -141323
rect -76765 -141331 -76721 -141323
rect -76665 -141331 -76621 -141323
rect -76565 -141331 -76521 -141323
rect -76465 -141331 -76421 -141323
rect -76365 -141331 -76321 -141323
rect -76265 -141331 -76221 -141323
rect -76165 -141331 -76121 -141323
rect -76065 -141331 -76021 -141323
rect -75965 -141331 -75921 -141323
rect -75865 -141331 -75821 -141323
rect -75765 -141331 -75721 -141323
rect -83221 -141375 -83213 -141331
rect -83121 -141375 -83113 -141331
rect -83021 -141375 -83013 -141331
rect -82921 -141375 -82913 -141331
rect -82821 -141375 -82813 -141331
rect -82721 -141375 -82713 -141331
rect -82621 -141375 -82613 -141331
rect -82521 -141375 -82513 -141331
rect -82421 -141375 -82413 -141331
rect -82321 -141375 -82313 -141331
rect -82221 -141375 -82213 -141331
rect -82121 -141375 -82113 -141331
rect -82021 -141375 -82013 -141331
rect -81921 -141375 -81913 -141331
rect -81821 -141375 -81813 -141331
rect -81721 -141375 -81713 -141331
rect -81221 -141375 -81213 -141331
rect -81121 -141375 -81113 -141331
rect -81021 -141375 -81013 -141331
rect -80921 -141375 -80913 -141331
rect -80821 -141375 -80813 -141331
rect -80721 -141375 -80713 -141331
rect -80621 -141375 -80613 -141331
rect -80521 -141375 -80513 -141331
rect -80421 -141375 -80413 -141331
rect -80321 -141375 -80313 -141331
rect -80221 -141375 -80213 -141331
rect -80121 -141375 -80113 -141331
rect -80021 -141375 -80013 -141331
rect -79921 -141375 -79913 -141331
rect -79821 -141375 -79813 -141331
rect -79721 -141375 -79713 -141331
rect -79221 -141375 -79213 -141331
rect -79121 -141375 -79113 -141331
rect -79021 -141375 -79013 -141331
rect -78921 -141375 -78913 -141331
rect -78821 -141375 -78813 -141331
rect -78721 -141375 -78713 -141331
rect -78621 -141375 -78613 -141331
rect -78521 -141375 -78513 -141331
rect -78421 -141375 -78413 -141331
rect -78321 -141375 -78313 -141331
rect -78221 -141375 -78213 -141331
rect -78121 -141375 -78113 -141331
rect -78021 -141375 -78013 -141331
rect -77921 -141375 -77913 -141331
rect -77821 -141375 -77813 -141331
rect -77721 -141375 -77713 -141331
rect -77221 -141375 -77213 -141331
rect -77121 -141375 -77113 -141331
rect -77021 -141375 -77013 -141331
rect -76921 -141375 -76913 -141331
rect -76821 -141375 -76813 -141331
rect -76721 -141375 -76713 -141331
rect -76621 -141375 -76613 -141331
rect -76521 -141375 -76513 -141331
rect -76421 -141375 -76413 -141331
rect -76321 -141375 -76313 -141331
rect -76221 -141375 -76213 -141331
rect -76121 -141375 -76113 -141331
rect -76021 -141375 -76013 -141331
rect -75921 -141375 -75913 -141331
rect -75821 -141375 -75813 -141331
rect -75721 -141375 -75713 -141331
rect -83265 -141431 -83221 -141423
rect -83165 -141431 -83121 -141423
rect -83065 -141431 -83021 -141423
rect -82965 -141431 -82921 -141423
rect -82865 -141431 -82821 -141423
rect -82765 -141431 -82721 -141423
rect -82665 -141431 -82621 -141423
rect -82565 -141431 -82521 -141423
rect -82465 -141431 -82421 -141423
rect -82365 -141431 -82321 -141423
rect -82265 -141431 -82221 -141423
rect -82165 -141431 -82121 -141423
rect -82065 -141431 -82021 -141423
rect -81965 -141431 -81921 -141423
rect -81865 -141431 -81821 -141423
rect -81765 -141431 -81721 -141423
rect -81265 -141431 -81221 -141423
rect -81165 -141431 -81121 -141423
rect -81065 -141431 -81021 -141423
rect -80965 -141431 -80921 -141423
rect -80865 -141431 -80821 -141423
rect -80765 -141431 -80721 -141423
rect -80665 -141431 -80621 -141423
rect -80565 -141431 -80521 -141423
rect -80465 -141431 -80421 -141423
rect -80365 -141431 -80321 -141423
rect -80265 -141431 -80221 -141423
rect -80165 -141431 -80121 -141423
rect -80065 -141431 -80021 -141423
rect -79965 -141431 -79921 -141423
rect -79865 -141431 -79821 -141423
rect -79765 -141431 -79721 -141423
rect -79265 -141431 -79221 -141423
rect -79165 -141431 -79121 -141423
rect -79065 -141431 -79021 -141423
rect -78965 -141431 -78921 -141423
rect -78865 -141431 -78821 -141423
rect -78765 -141431 -78721 -141423
rect -78665 -141431 -78621 -141423
rect -78565 -141431 -78521 -141423
rect -78465 -141431 -78421 -141423
rect -78365 -141431 -78321 -141423
rect -78265 -141431 -78221 -141423
rect -78165 -141431 -78121 -141423
rect -78065 -141431 -78021 -141423
rect -77965 -141431 -77921 -141423
rect -77865 -141431 -77821 -141423
rect -77765 -141431 -77721 -141423
rect -77265 -141431 -77221 -141423
rect -77165 -141431 -77121 -141423
rect -77065 -141431 -77021 -141423
rect -76965 -141431 -76921 -141423
rect -76865 -141431 -76821 -141423
rect -76765 -141431 -76721 -141423
rect -76665 -141431 -76621 -141423
rect -76565 -141431 -76521 -141423
rect -76465 -141431 -76421 -141423
rect -76365 -141431 -76321 -141423
rect -76265 -141431 -76221 -141423
rect -76165 -141431 -76121 -141423
rect -76065 -141431 -76021 -141423
rect -75965 -141431 -75921 -141423
rect -75865 -141431 -75821 -141423
rect -75765 -141431 -75721 -141423
rect -83221 -141475 -83213 -141431
rect -83121 -141475 -83113 -141431
rect -83021 -141475 -83013 -141431
rect -82921 -141475 -82913 -141431
rect -82821 -141475 -82813 -141431
rect -82721 -141475 -82713 -141431
rect -82621 -141475 -82613 -141431
rect -82521 -141475 -82513 -141431
rect -82421 -141475 -82413 -141431
rect -82321 -141475 -82313 -141431
rect -82221 -141475 -82213 -141431
rect -82121 -141475 -82113 -141431
rect -82021 -141475 -82013 -141431
rect -81921 -141475 -81913 -141431
rect -81821 -141475 -81813 -141431
rect -81721 -141475 -81713 -141431
rect -81221 -141475 -81213 -141431
rect -81121 -141475 -81113 -141431
rect -81021 -141475 -81013 -141431
rect -80921 -141475 -80913 -141431
rect -80821 -141475 -80813 -141431
rect -80721 -141475 -80713 -141431
rect -80621 -141475 -80613 -141431
rect -80521 -141475 -80513 -141431
rect -80421 -141475 -80413 -141431
rect -80321 -141475 -80313 -141431
rect -80221 -141475 -80213 -141431
rect -80121 -141475 -80113 -141431
rect -80021 -141475 -80013 -141431
rect -79921 -141475 -79913 -141431
rect -79821 -141475 -79813 -141431
rect -79721 -141475 -79713 -141431
rect -79221 -141475 -79213 -141431
rect -79121 -141475 -79113 -141431
rect -79021 -141475 -79013 -141431
rect -78921 -141475 -78913 -141431
rect -78821 -141475 -78813 -141431
rect -78721 -141475 -78713 -141431
rect -78621 -141475 -78613 -141431
rect -78521 -141475 -78513 -141431
rect -78421 -141475 -78413 -141431
rect -78321 -141475 -78313 -141431
rect -78221 -141475 -78213 -141431
rect -78121 -141475 -78113 -141431
rect -78021 -141475 -78013 -141431
rect -77921 -141475 -77913 -141431
rect -77821 -141475 -77813 -141431
rect -77721 -141475 -77713 -141431
rect -77221 -141475 -77213 -141431
rect -77121 -141475 -77113 -141431
rect -77021 -141475 -77013 -141431
rect -76921 -141475 -76913 -141431
rect -76821 -141475 -76813 -141431
rect -76721 -141475 -76713 -141431
rect -76621 -141475 -76613 -141431
rect -76521 -141475 -76513 -141431
rect -76421 -141475 -76413 -141431
rect -76321 -141475 -76313 -141431
rect -76221 -141475 -76213 -141431
rect -76121 -141475 -76113 -141431
rect -76021 -141475 -76013 -141431
rect -75921 -141475 -75913 -141431
rect -75821 -141475 -75813 -141431
rect -75721 -141475 -75713 -141431
rect -83265 -141531 -83221 -141523
rect -83165 -141531 -83121 -141523
rect -83065 -141531 -83021 -141523
rect -82965 -141531 -82921 -141523
rect -82865 -141531 -82821 -141523
rect -82765 -141531 -82721 -141523
rect -82665 -141531 -82621 -141523
rect -82565 -141531 -82521 -141523
rect -82465 -141531 -82421 -141523
rect -82365 -141531 -82321 -141523
rect -82265 -141531 -82221 -141523
rect -82165 -141531 -82121 -141523
rect -82065 -141531 -82021 -141523
rect -81965 -141531 -81921 -141523
rect -81865 -141531 -81821 -141523
rect -81765 -141531 -81721 -141523
rect -81265 -141531 -81221 -141523
rect -81165 -141531 -81121 -141523
rect -81065 -141531 -81021 -141523
rect -80965 -141531 -80921 -141523
rect -80865 -141531 -80821 -141523
rect -80765 -141531 -80721 -141523
rect -80665 -141531 -80621 -141523
rect -80565 -141531 -80521 -141523
rect -80465 -141531 -80421 -141523
rect -80365 -141531 -80321 -141523
rect -80265 -141531 -80221 -141523
rect -80165 -141531 -80121 -141523
rect -80065 -141531 -80021 -141523
rect -79965 -141531 -79921 -141523
rect -79865 -141531 -79821 -141523
rect -79765 -141531 -79721 -141523
rect -79265 -141531 -79221 -141523
rect -79165 -141531 -79121 -141523
rect -79065 -141531 -79021 -141523
rect -78965 -141531 -78921 -141523
rect -78865 -141531 -78821 -141523
rect -78765 -141531 -78721 -141523
rect -78665 -141531 -78621 -141523
rect -78565 -141531 -78521 -141523
rect -78465 -141531 -78421 -141523
rect -78365 -141531 -78321 -141523
rect -78265 -141531 -78221 -141523
rect -78165 -141531 -78121 -141523
rect -78065 -141531 -78021 -141523
rect -77965 -141531 -77921 -141523
rect -77865 -141531 -77821 -141523
rect -77765 -141531 -77721 -141523
rect -77265 -141531 -77221 -141523
rect -77165 -141531 -77121 -141523
rect -77065 -141531 -77021 -141523
rect -76965 -141531 -76921 -141523
rect -76865 -141531 -76821 -141523
rect -76765 -141531 -76721 -141523
rect -76665 -141531 -76621 -141523
rect -76565 -141531 -76521 -141523
rect -76465 -141531 -76421 -141523
rect -76365 -141531 -76321 -141523
rect -76265 -141531 -76221 -141523
rect -76165 -141531 -76121 -141523
rect -76065 -141531 -76021 -141523
rect -75965 -141531 -75921 -141523
rect -75865 -141531 -75821 -141523
rect -75765 -141531 -75721 -141523
rect -83221 -141575 -83213 -141531
rect -83121 -141575 -83113 -141531
rect -83021 -141575 -83013 -141531
rect -82921 -141575 -82913 -141531
rect -82821 -141575 -82813 -141531
rect -82721 -141575 -82713 -141531
rect -82621 -141575 -82613 -141531
rect -82521 -141575 -82513 -141531
rect -82421 -141575 -82413 -141531
rect -82321 -141575 -82313 -141531
rect -82221 -141575 -82213 -141531
rect -82121 -141575 -82113 -141531
rect -82021 -141575 -82013 -141531
rect -81921 -141575 -81913 -141531
rect -81821 -141575 -81813 -141531
rect -81721 -141575 -81713 -141531
rect -81221 -141575 -81213 -141531
rect -81121 -141575 -81113 -141531
rect -81021 -141575 -81013 -141531
rect -80921 -141575 -80913 -141531
rect -80821 -141575 -80813 -141531
rect -80721 -141575 -80713 -141531
rect -80621 -141575 -80613 -141531
rect -80521 -141575 -80513 -141531
rect -80421 -141575 -80413 -141531
rect -80321 -141575 -80313 -141531
rect -80221 -141575 -80213 -141531
rect -80121 -141575 -80113 -141531
rect -80021 -141575 -80013 -141531
rect -79921 -141575 -79913 -141531
rect -79821 -141575 -79813 -141531
rect -79721 -141575 -79713 -141531
rect -79221 -141575 -79213 -141531
rect -79121 -141575 -79113 -141531
rect -79021 -141575 -79013 -141531
rect -78921 -141575 -78913 -141531
rect -78821 -141575 -78813 -141531
rect -78721 -141575 -78713 -141531
rect -78621 -141575 -78613 -141531
rect -78521 -141575 -78513 -141531
rect -78421 -141575 -78413 -141531
rect -78321 -141575 -78313 -141531
rect -78221 -141575 -78213 -141531
rect -78121 -141575 -78113 -141531
rect -78021 -141575 -78013 -141531
rect -77921 -141575 -77913 -141531
rect -77821 -141575 -77813 -141531
rect -77721 -141575 -77713 -141531
rect -77221 -141575 -77213 -141531
rect -77121 -141575 -77113 -141531
rect -77021 -141575 -77013 -141531
rect -76921 -141575 -76913 -141531
rect -76821 -141575 -76813 -141531
rect -76721 -141575 -76713 -141531
rect -76621 -141575 -76613 -141531
rect -76521 -141575 -76513 -141531
rect -76421 -141575 -76413 -141531
rect -76321 -141575 -76313 -141531
rect -76221 -141575 -76213 -141531
rect -76121 -141575 -76113 -141531
rect -76021 -141575 -76013 -141531
rect -75921 -141575 -75913 -141531
rect -75821 -141575 -75813 -141531
rect -75721 -141575 -75713 -141531
rect -83265 -141631 -83221 -141623
rect -83165 -141631 -83121 -141623
rect -83065 -141631 -83021 -141623
rect -82965 -141631 -82921 -141623
rect -82865 -141631 -82821 -141623
rect -82765 -141631 -82721 -141623
rect -82665 -141631 -82621 -141623
rect -82565 -141631 -82521 -141623
rect -82465 -141631 -82421 -141623
rect -82365 -141631 -82321 -141623
rect -82265 -141631 -82221 -141623
rect -82165 -141631 -82121 -141623
rect -82065 -141631 -82021 -141623
rect -81965 -141631 -81921 -141623
rect -81865 -141631 -81821 -141623
rect -81765 -141631 -81721 -141623
rect -81265 -141631 -81221 -141623
rect -81165 -141631 -81121 -141623
rect -81065 -141631 -81021 -141623
rect -80965 -141631 -80921 -141623
rect -80865 -141631 -80821 -141623
rect -80765 -141631 -80721 -141623
rect -80665 -141631 -80621 -141623
rect -80565 -141631 -80521 -141623
rect -80465 -141631 -80421 -141623
rect -80365 -141631 -80321 -141623
rect -80265 -141631 -80221 -141623
rect -80165 -141631 -80121 -141623
rect -80065 -141631 -80021 -141623
rect -79965 -141631 -79921 -141623
rect -79865 -141631 -79821 -141623
rect -79765 -141631 -79721 -141623
rect -79265 -141631 -79221 -141623
rect -79165 -141631 -79121 -141623
rect -79065 -141631 -79021 -141623
rect -78965 -141631 -78921 -141623
rect -78865 -141631 -78821 -141623
rect -78765 -141631 -78721 -141623
rect -78665 -141631 -78621 -141623
rect -78565 -141631 -78521 -141623
rect -78465 -141631 -78421 -141623
rect -78365 -141631 -78321 -141623
rect -78265 -141631 -78221 -141623
rect -78165 -141631 -78121 -141623
rect -78065 -141631 -78021 -141623
rect -77965 -141631 -77921 -141623
rect -77865 -141631 -77821 -141623
rect -77765 -141631 -77721 -141623
rect -77265 -141631 -77221 -141623
rect -77165 -141631 -77121 -141623
rect -77065 -141631 -77021 -141623
rect -76965 -141631 -76921 -141623
rect -76865 -141631 -76821 -141623
rect -76765 -141631 -76721 -141623
rect -76665 -141631 -76621 -141623
rect -76565 -141631 -76521 -141623
rect -76465 -141631 -76421 -141623
rect -76365 -141631 -76321 -141623
rect -76265 -141631 -76221 -141623
rect -76165 -141631 -76121 -141623
rect -76065 -141631 -76021 -141623
rect -75965 -141631 -75921 -141623
rect -75865 -141631 -75821 -141623
rect -75765 -141631 -75721 -141623
rect -83221 -141675 -83213 -141631
rect -83121 -141675 -83113 -141631
rect -83021 -141675 -83013 -141631
rect -82921 -141675 -82913 -141631
rect -82821 -141675 -82813 -141631
rect -82721 -141675 -82713 -141631
rect -82621 -141675 -82613 -141631
rect -82521 -141675 -82513 -141631
rect -82421 -141675 -82413 -141631
rect -82321 -141675 -82313 -141631
rect -82221 -141675 -82213 -141631
rect -82121 -141675 -82113 -141631
rect -82021 -141675 -82013 -141631
rect -81921 -141675 -81913 -141631
rect -81821 -141675 -81813 -141631
rect -81721 -141675 -81713 -141631
rect -81221 -141675 -81213 -141631
rect -81121 -141675 -81113 -141631
rect -81021 -141675 -81013 -141631
rect -80921 -141675 -80913 -141631
rect -80821 -141675 -80813 -141631
rect -80721 -141675 -80713 -141631
rect -80621 -141675 -80613 -141631
rect -80521 -141675 -80513 -141631
rect -80421 -141675 -80413 -141631
rect -80321 -141675 -80313 -141631
rect -80221 -141675 -80213 -141631
rect -80121 -141675 -80113 -141631
rect -80021 -141675 -80013 -141631
rect -79921 -141675 -79913 -141631
rect -79821 -141675 -79813 -141631
rect -79721 -141675 -79713 -141631
rect -79221 -141675 -79213 -141631
rect -79121 -141675 -79113 -141631
rect -79021 -141675 -79013 -141631
rect -78921 -141675 -78913 -141631
rect -78821 -141675 -78813 -141631
rect -78721 -141675 -78713 -141631
rect -78621 -141675 -78613 -141631
rect -78521 -141675 -78513 -141631
rect -78421 -141675 -78413 -141631
rect -78321 -141675 -78313 -141631
rect -78221 -141675 -78213 -141631
rect -78121 -141675 -78113 -141631
rect -78021 -141675 -78013 -141631
rect -77921 -141675 -77913 -141631
rect -77821 -141675 -77813 -141631
rect -77721 -141675 -77713 -141631
rect -77221 -141675 -77213 -141631
rect -77121 -141675 -77113 -141631
rect -77021 -141675 -77013 -141631
rect -76921 -141675 -76913 -141631
rect -76821 -141675 -76813 -141631
rect -76721 -141675 -76713 -141631
rect -76621 -141675 -76613 -141631
rect -76521 -141675 -76513 -141631
rect -76421 -141675 -76413 -141631
rect -76321 -141675 -76313 -141631
rect -76221 -141675 -76213 -141631
rect -76121 -141675 -76113 -141631
rect -76021 -141675 -76013 -141631
rect -75921 -141675 -75913 -141631
rect -75821 -141675 -75813 -141631
rect -75721 -141675 -75713 -141631
rect -83265 -141731 -83221 -141723
rect -83165 -141731 -83121 -141723
rect -83065 -141731 -83021 -141723
rect -82965 -141731 -82921 -141723
rect -82865 -141731 -82821 -141723
rect -82765 -141731 -82721 -141723
rect -82665 -141731 -82621 -141723
rect -82565 -141731 -82521 -141723
rect -82465 -141731 -82421 -141723
rect -82365 -141731 -82321 -141723
rect -82265 -141731 -82221 -141723
rect -82165 -141731 -82121 -141723
rect -82065 -141731 -82021 -141723
rect -81965 -141731 -81921 -141723
rect -81865 -141731 -81821 -141723
rect -81765 -141731 -81721 -141723
rect -81265 -141731 -81221 -141723
rect -81165 -141731 -81121 -141723
rect -81065 -141731 -81021 -141723
rect -80965 -141731 -80921 -141723
rect -80865 -141731 -80821 -141723
rect -80765 -141731 -80721 -141723
rect -80665 -141731 -80621 -141723
rect -80565 -141731 -80521 -141723
rect -80465 -141731 -80421 -141723
rect -80365 -141731 -80321 -141723
rect -80265 -141731 -80221 -141723
rect -80165 -141731 -80121 -141723
rect -80065 -141731 -80021 -141723
rect -79965 -141731 -79921 -141723
rect -79865 -141731 -79821 -141723
rect -79765 -141731 -79721 -141723
rect -79265 -141731 -79221 -141723
rect -79165 -141731 -79121 -141723
rect -79065 -141731 -79021 -141723
rect -78965 -141731 -78921 -141723
rect -78865 -141731 -78821 -141723
rect -78765 -141731 -78721 -141723
rect -78665 -141731 -78621 -141723
rect -78565 -141731 -78521 -141723
rect -78465 -141731 -78421 -141723
rect -78365 -141731 -78321 -141723
rect -78265 -141731 -78221 -141723
rect -78165 -141731 -78121 -141723
rect -78065 -141731 -78021 -141723
rect -77965 -141731 -77921 -141723
rect -77865 -141731 -77821 -141723
rect -77765 -141731 -77721 -141723
rect -77265 -141731 -77221 -141723
rect -77165 -141731 -77121 -141723
rect -77065 -141731 -77021 -141723
rect -76965 -141731 -76921 -141723
rect -76865 -141731 -76821 -141723
rect -76765 -141731 -76721 -141723
rect -76665 -141731 -76621 -141723
rect -76565 -141731 -76521 -141723
rect -76465 -141731 -76421 -141723
rect -76365 -141731 -76321 -141723
rect -76265 -141731 -76221 -141723
rect -76165 -141731 -76121 -141723
rect -76065 -141731 -76021 -141723
rect -75965 -141731 -75921 -141723
rect -75865 -141731 -75821 -141723
rect -75765 -141731 -75721 -141723
rect -83221 -141775 -83213 -141731
rect -83121 -141775 -83113 -141731
rect -83021 -141775 -83013 -141731
rect -82921 -141775 -82913 -141731
rect -82821 -141775 -82813 -141731
rect -82721 -141775 -82713 -141731
rect -82621 -141775 -82613 -141731
rect -82521 -141775 -82513 -141731
rect -82421 -141775 -82413 -141731
rect -82321 -141775 -82313 -141731
rect -82221 -141775 -82213 -141731
rect -82121 -141775 -82113 -141731
rect -82021 -141775 -82013 -141731
rect -81921 -141775 -81913 -141731
rect -81821 -141775 -81813 -141731
rect -81721 -141775 -81713 -141731
rect -81221 -141775 -81213 -141731
rect -81121 -141775 -81113 -141731
rect -81021 -141775 -81013 -141731
rect -80921 -141775 -80913 -141731
rect -80821 -141775 -80813 -141731
rect -80721 -141775 -80713 -141731
rect -80621 -141775 -80613 -141731
rect -80521 -141775 -80513 -141731
rect -80421 -141775 -80413 -141731
rect -80321 -141775 -80313 -141731
rect -80221 -141775 -80213 -141731
rect -80121 -141775 -80113 -141731
rect -80021 -141775 -80013 -141731
rect -79921 -141775 -79913 -141731
rect -79821 -141775 -79813 -141731
rect -79721 -141775 -79713 -141731
rect -79221 -141775 -79213 -141731
rect -79121 -141775 -79113 -141731
rect -79021 -141775 -79013 -141731
rect -78921 -141775 -78913 -141731
rect -78821 -141775 -78813 -141731
rect -78721 -141775 -78713 -141731
rect -78621 -141775 -78613 -141731
rect -78521 -141775 -78513 -141731
rect -78421 -141775 -78413 -141731
rect -78321 -141775 -78313 -141731
rect -78221 -141775 -78213 -141731
rect -78121 -141775 -78113 -141731
rect -78021 -141775 -78013 -141731
rect -77921 -141775 -77913 -141731
rect -77821 -141775 -77813 -141731
rect -77721 -141775 -77713 -141731
rect -77221 -141775 -77213 -141731
rect -77121 -141775 -77113 -141731
rect -77021 -141775 -77013 -141731
rect -76921 -141775 -76913 -141731
rect -76821 -141775 -76813 -141731
rect -76721 -141775 -76713 -141731
rect -76621 -141775 -76613 -141731
rect -76521 -141775 -76513 -141731
rect -76421 -141775 -76413 -141731
rect -76321 -141775 -76313 -141731
rect -76221 -141775 -76213 -141731
rect -76121 -141775 -76113 -141731
rect -76021 -141775 -76013 -141731
rect -75921 -141775 -75913 -141731
rect -75821 -141775 -75813 -141731
rect -75721 -141775 -75713 -141731
rect -98040 -162683 -98038 -150683
rect -97974 -162683 -97972 -150683
rect -60162 -162352 -60160 -142352
rect -60096 -162352 -60094 -142352
rect -26162 -162352 -26160 -142352
rect -26096 -162352 -26094 -142352
rect 7838 -162352 7840 -142352
rect 7904 -162352 7906 -142352
rect 41838 -162352 41840 -142352
rect 41904 -162352 41906 -142352
rect 75838 -162352 75840 -142352
rect 75904 -162352 75906 -142352
rect 109838 -162352 109840 -142352
rect 109904 -162352 109906 -142352
rect 143838 -162352 143840 -142352
rect 143904 -162352 143906 -142352
<< nwell >>
rect -14513 -14331 -4723 -6461
<< pwell >>
rect -109798 -48705 -78056 -27758
rect -77798 -48705 -46056 -27758
rect -45798 -48705 -14056 -27758
rect -13798 -48705 17944 -27758
rect 18202 -48705 49944 -27758
rect 50202 -48705 81944 -27758
rect 82202 -48705 113944 -27758
rect 114202 -48705 145944 -27758
rect 146202 -48705 177944 -27758
rect -109798 -74705 -78056 -53758
rect -77798 -74705 -46056 -53758
rect -45798 -74705 -14056 -53758
rect -13798 -74705 17944 -53758
rect 18202 -74705 49944 -53758
rect 50202 -74705 81944 -53758
rect 82202 -74705 113944 -53758
rect 114202 -74705 145944 -53758
rect 146202 -74705 177944 -53758
rect -109798 -103705 -78056 -82740
rect -77798 -103705 -46056 -82740
rect -45798 -103705 -14056 -82740
rect -13798 -103705 17944 -82740
rect 18202 -103705 49944 -82740
rect 50202 -103705 81944 -82740
rect 82202 -103705 113944 -82740
rect 114202 -103705 145944 -82740
rect 146202 -103705 177944 -82740
rect -109798 -129705 -78056 -108750
rect -77798 -129705 -46056 -108750
rect -45798 -129705 -14056 -108750
rect -13798 -129705 17944 -108750
rect 18202 -129705 49944 -108750
rect 50202 -129705 81944 -108750
rect 82202 -129705 113944 -108750
rect 114202 -129705 145944 -108750
rect 146202 -129705 177944 -108750
rect -106346 -143362 -104700 -138197
rect -98619 -163033 -79246 -150224
rect -60780 -162938 -29038 -142038
rect -26780 -162938 4962 -142038
rect 7220 -162938 38962 -142038
rect 41220 -162938 72962 -142038
rect 75220 -162938 106962 -142038
rect 109220 -162938 140962 -142038
rect 143220 -162938 174962 -142038
<< nsubdiff >>
rect -14393 -6941 -4843 -6581
rect -14393 -7230 -14033 -6941
rect -14393 -7452 -14324 -7230
rect -14102 -7452 -14033 -7230
rect -5203 -7230 -4843 -6941
rect -14393 -7700 -14033 -7452
rect -14393 -7922 -14324 -7700
rect -14102 -7922 -14033 -7700
rect -14393 -8170 -14033 -7922
rect -14393 -8392 -14324 -8170
rect -14102 -8392 -14033 -8170
rect -14393 -8640 -14033 -8392
rect -14393 -8862 -14324 -8640
rect -14102 -8862 -14033 -8640
rect -14393 -9110 -14033 -8862
rect -14393 -9332 -14324 -9110
rect -14102 -9332 -14033 -9110
rect -14393 -9580 -14033 -9332
rect -14393 -9802 -14324 -9580
rect -14102 -9802 -14033 -9580
rect -14393 -10050 -14033 -9802
rect -14393 -10272 -14324 -10050
rect -14102 -10272 -14033 -10050
rect -14393 -10520 -14033 -10272
rect -14393 -10742 -14324 -10520
rect -14102 -10742 -14033 -10520
rect -14393 -10990 -14033 -10742
rect -14393 -11212 -14324 -10990
rect -14102 -11212 -14033 -10990
rect -14393 -11460 -14033 -11212
rect -14393 -11682 -14324 -11460
rect -14102 -11682 -14033 -11460
rect -14393 -11930 -14033 -11682
rect -14393 -12152 -14324 -11930
rect -14102 -12152 -14033 -11930
rect -14393 -12400 -14033 -12152
rect -14393 -12622 -14324 -12400
rect -14102 -12622 -14033 -12400
rect -14393 -12870 -14033 -12622
rect -14393 -13092 -14324 -12870
rect -14102 -13092 -14033 -12870
rect -14393 -13340 -14033 -13092
rect -14393 -13562 -14324 -13340
rect -14102 -13562 -14033 -13340
rect -5203 -7452 -5134 -7230
rect -4912 -7452 -4843 -7230
rect -5203 -7700 -4843 -7452
rect -5203 -7922 -5134 -7700
rect -4912 -7922 -4843 -7700
rect -5203 -8170 -4843 -7922
rect -5203 -8392 -5134 -8170
rect -4912 -8392 -4843 -8170
rect -5203 -8640 -4843 -8392
rect -5203 -8862 -5134 -8640
rect -4912 -8862 -4843 -8640
rect -5203 -9110 -4843 -8862
rect -5203 -9332 -5134 -9110
rect -4912 -9332 -4843 -9110
rect -5203 -9580 -4843 -9332
rect -5203 -9802 -5134 -9580
rect -4912 -9802 -4843 -9580
rect -5203 -10050 -4843 -9802
rect -5203 -10272 -5134 -10050
rect -4912 -10272 -4843 -10050
rect -5203 -10520 -4843 -10272
rect -5203 -10742 -5134 -10520
rect -4912 -10742 -4843 -10520
rect -5203 -10990 -4843 -10742
rect -5203 -11212 -5134 -10990
rect -4912 -11212 -4843 -10990
rect -5203 -11460 -4843 -11212
rect -5203 -11682 -5134 -11460
rect -4912 -11682 -4843 -11460
rect -5203 -11930 -4843 -11682
rect -5203 -12152 -5134 -11930
rect -4912 -12152 -4843 -11930
rect -5203 -12400 -4843 -12152
rect -5203 -12622 -5134 -12400
rect -4912 -12622 -4843 -12400
rect -5203 -12870 -4843 -12622
rect -5203 -13092 -5134 -12870
rect -4912 -13092 -4843 -12870
rect -5203 -13340 -4843 -13092
rect -14393 -13851 -14033 -13562
rect -5203 -13562 -5134 -13340
rect -4912 -13562 -4843 -13340
rect -5203 -13851 -4843 -13562
rect -14393 -14211 -4843 -13851
<< nsubdiffcont >>
rect -14324 -7452 -14102 -7230
rect -14324 -7922 -14102 -7700
rect -14324 -8392 -14102 -8170
rect -14324 -8862 -14102 -8640
rect -14324 -9332 -14102 -9110
rect -14324 -9802 -14102 -9580
rect -14324 -10272 -14102 -10050
rect -14324 -10742 -14102 -10520
rect -14324 -11212 -14102 -10990
rect -14324 -11682 -14102 -11460
rect -14324 -12152 -14102 -11930
rect -14324 -12622 -14102 -12400
rect -14324 -13092 -14102 -12870
rect -14324 -13562 -14102 -13340
rect -5134 -7452 -4912 -7230
rect -5134 -7922 -4912 -7700
rect -5134 -8392 -4912 -8170
rect -5134 -8862 -4912 -8640
rect -5134 -9332 -4912 -9110
rect -5134 -9802 -4912 -9580
rect -5134 -10272 -4912 -10050
rect -5134 -10742 -4912 -10520
rect -5134 -11212 -4912 -10990
rect -5134 -11682 -4912 -11460
rect -5134 -12152 -4912 -11930
rect -5134 -12622 -4912 -12400
rect -5134 -13092 -4912 -12870
rect -5134 -13562 -4912 -13340
<< polysilicon >>
rect -36844 25369 -16844 27192
rect -36844 24319 -32735 25369
rect -31594 24319 -16844 25369
rect 58104 25351 109400 25613
rect -36844 7469 -16844 24319
rect -18 9998 53078 10300
rect -36844 7192 -6294 7469
rect -6694 6110 -6294 7192
rect 58104 3752 109400 5263
rect 55047 3509 109400 3752
rect 55047 2563 55404 3509
rect 55450 2563 109400 3509
rect 55047 2375 109400 2563
rect 58104 351 109400 2375
rect -18 -970 25078 -90
rect -18 -1016 2307 -970
rect 22253 -1016 25078 -970
rect -18 -1233 25078 -1016
rect -13593 -7450 -5643 -7381
rect -13593 -7672 -13489 -7450
rect -13267 -7672 -13019 -7450
rect -12797 -7672 -12549 -7450
rect -12327 -7672 -12079 -7450
rect -11857 -7672 -11609 -7450
rect -11387 -7672 -11139 -7450
rect -10917 -7672 -10669 -7450
rect -10447 -7672 -10199 -7450
rect -9977 -7672 -9729 -7450
rect -9507 -7672 -9259 -7450
rect -9037 -7672 -8789 -7450
rect -8567 -7672 -8319 -7450
rect -8097 -7672 -7849 -7450
rect -7627 -7672 -7379 -7450
rect -7157 -7672 -6909 -7450
rect -6687 -7672 -6439 -7450
rect -6217 -7672 -5969 -7450
rect -5747 -7672 -5643 -7450
rect -13593 -7896 -5643 -7672
rect -13593 -13120 -5643 -12896
rect -13593 -13342 -13489 -13120
rect -13267 -13342 -13019 -13120
rect -12797 -13342 -12549 -13120
rect -12327 -13342 -12079 -13120
rect -11857 -13342 -11609 -13120
rect -11387 -13342 -11139 -13120
rect -10917 -13342 -10669 -13120
rect -10447 -13342 -10199 -13120
rect -9977 -13342 -9729 -13120
rect -9507 -13342 -9259 -13120
rect -9037 -13342 -8789 -13120
rect -8567 -13342 -8319 -13120
rect -8097 -13342 -7849 -13120
rect -7627 -13342 -7379 -13120
rect -7157 -13342 -6909 -13120
rect -6687 -13342 -6439 -13120
rect -6217 -13342 -5969 -13120
rect -5747 -13342 -5643 -13120
rect -13593 -13411 -5643 -13342
rect -109026 -28075 -78730 -27418
rect -77026 -28075 -46730 -27418
rect -45026 -28075 -14730 -27418
rect -13026 -28075 17270 -27418
rect 18974 -28075 49270 -27418
rect 50974 -28075 81270 -27418
rect 82974 -28075 113270 -27418
rect 114974 -28075 145270 -27418
rect 146974 -28075 177270 -27418
rect -135098 -34142 -115098 -32005
rect -135098 -35301 -130077 -34142
rect -128909 -35301 -115098 -34142
rect -135098 -50407 -115098 -35301
rect -109026 -50407 177270 -48163
rect -135098 -52005 177270 -50407
rect -109026 -53418 177270 -52005
rect -109026 -54075 -78730 -53418
rect -77026 -54075 -46730 -53418
rect -45026 -54075 -14730 -53418
rect -13026 -54075 17270 -53418
rect 18974 -54075 49270 -53418
rect 50974 -54075 81270 -53418
rect 82974 -54075 113270 -53418
rect 114974 -54075 145270 -53418
rect 146974 -54075 177270 -53418
rect -109026 -83075 -78730 -82418
rect -77026 -83075 -46730 -82418
rect -45026 -83075 -14730 -82418
rect -13026 -83075 17270 -82418
rect 18974 -83075 49270 -82418
rect 50974 -83075 81270 -82418
rect 82974 -83075 113270 -82418
rect 114974 -83075 145270 -82418
rect 146974 -83075 177270 -82418
rect 179273 -95506 199273 -87181
rect 179273 -96423 185033 -95506
rect 185843 -96423 199273 -95506
rect -109026 -104817 177270 -103163
rect 179273 -104817 199273 -96423
rect -109026 -107181 199273 -104817
rect -109026 -108418 177270 -107181
rect -109026 -109075 -78730 -108418
rect -77026 -109075 -46730 -108418
rect -45026 -109075 -14730 -108418
rect -13026 -109075 17270 -108418
rect 18974 -109075 49270 -108418
rect 50974 -109075 81270 -108418
rect 82974 -109075 113270 -108418
rect 114974 -109075 145270 -108418
rect 146974 -109075 177270 -108418
rect -91201 -139838 -55139 -137922
rect -91201 -142398 -89852 -139838
rect -60008 -141877 -55139 -139838
rect -60008 -142308 174288 -141877
rect -103886 -142610 -79750 -142398
rect -105574 -145043 -105374 -142827
rect -103886 -143556 -103394 -142610
rect -102448 -143556 -79750 -142610
rect -103886 -143790 -79750 -143556
rect -97886 -145043 -79750 -143790
rect -105574 -145768 -79750 -145043
rect -97886 -150639 -79750 -145768
<< polycontact >>
rect -32735 24319 -31594 25369
rect 55404 2563 55450 3509
rect 2307 -1016 22253 -970
rect -13489 -7672 -13267 -7450
rect -13019 -7672 -12797 -7450
rect -12549 -7672 -12327 -7450
rect -12079 -7672 -11857 -7450
rect -11609 -7672 -11387 -7450
rect -11139 -7672 -10917 -7450
rect -10669 -7672 -10447 -7450
rect -10199 -7672 -9977 -7450
rect -9729 -7672 -9507 -7450
rect -9259 -7672 -9037 -7450
rect -8789 -7672 -8567 -7450
rect -8319 -7672 -8097 -7450
rect -7849 -7672 -7627 -7450
rect -7379 -7672 -7157 -7450
rect -6909 -7672 -6687 -7450
rect -6439 -7672 -6217 -7450
rect -5969 -7672 -5747 -7450
rect -13489 -13342 -13267 -13120
rect -13019 -13342 -12797 -13120
rect -12549 -13342 -12327 -13120
rect -12079 -13342 -11857 -13120
rect -11609 -13342 -11387 -13120
rect -11139 -13342 -10917 -13120
rect -10669 -13342 -10447 -13120
rect -10199 -13342 -9977 -13120
rect -9729 -13342 -9507 -13120
rect -9259 -13342 -9037 -13120
rect -8789 -13342 -8567 -13120
rect -8319 -13342 -8097 -13120
rect -7849 -13342 -7627 -13120
rect -7379 -13342 -7157 -13120
rect -6909 -13342 -6687 -13120
rect -6439 -13342 -6217 -13120
rect -5969 -13342 -5747 -13120
rect -130077 -35301 -128909 -34142
rect 185033 -96423 185843 -95506
rect -103394 -143556 -102448 -142610
<< ppolyres >>
rect -13593 -12896 -5643 -7896
<< metal1 >>
rect -13548 29110 109861 32249
rect -33873 25369 -23600 27192
rect -33873 24319 -32735 25369
rect -31594 24319 -23600 25369
rect -33873 20881 -23600 24319
rect -30138 3555 -17010 5889
rect -11550 4064 -6708 29110
rect -108 10678 25168 29110
rect -108 9956 -32 10678
rect 900 9956 976 10678
rect 1908 9956 1984 10678
rect 2916 9956 2992 10678
rect 3924 9956 4000 10678
rect 4932 9956 5008 10678
rect 5940 9956 6016 10678
rect 6948 9956 7024 10678
rect 7956 9956 8032 10678
rect 8964 9956 9040 10678
rect 9972 9956 10048 10678
rect 10980 9956 11056 10678
rect 11988 9956 12064 10678
rect 12996 9956 13072 10678
rect 14004 9956 14080 10678
rect 15012 9956 15088 10678
rect 16020 9956 16096 10678
rect 17028 9956 17104 10678
rect 18036 9956 18112 10678
rect 19044 9956 19120 10678
rect 20052 9956 20128 10678
rect 21060 9956 21136 10678
rect 22068 9956 22144 10678
rect 23076 9956 23152 10678
rect 24084 9956 24160 10678
rect 25092 9956 25168 10678
rect 27892 10678 53168 29110
rect 27892 9956 27968 10678
rect 28900 9956 28976 10678
rect 29908 9956 29984 10678
rect 30916 9956 30992 10678
rect 31924 9956 32000 10678
rect 32932 9956 33008 10678
rect 33940 9956 34016 10678
rect 34948 9956 35024 10678
rect 35956 9956 36032 10678
rect 36964 9956 37040 10678
rect 37972 9956 38048 10678
rect 38980 9956 39056 10678
rect 39988 9956 40064 10678
rect 40996 9956 41072 10678
rect 42004 9956 42080 10678
rect 43012 9956 43088 10678
rect 44020 9956 44096 10678
rect 45028 9956 45104 10678
rect 46036 9956 46112 10678
rect 47044 9956 47120 10678
rect 48052 9956 48128 10678
rect 49060 9956 49136 10678
rect 50068 9956 50144 10678
rect 51076 9956 51152 10678
rect 52084 9956 52160 10678
rect 53092 9956 53168 10678
rect 56492 25794 109490 29110
rect -30138 3511 -27407 3555
rect -27363 3511 -27307 3555
rect -27263 3511 -27207 3555
rect -27163 3511 -27107 3555
rect -27063 3511 -27007 3555
rect -26963 3511 -26907 3555
rect -26863 3511 -26807 3555
rect -26763 3511 -26707 3555
rect -26663 3511 -26607 3555
rect -26563 3511 -26507 3555
rect -26463 3511 -26407 3555
rect -26363 3511 -26307 3555
rect -26263 3511 -26207 3555
rect -26163 3511 -26107 3555
rect -26063 3511 -26007 3555
rect -25963 3511 -25907 3555
rect -25863 3511 -25407 3555
rect -25363 3511 -25307 3555
rect -25263 3511 -25207 3555
rect -25163 3511 -25107 3555
rect -25063 3511 -25007 3555
rect -24963 3511 -24907 3555
rect -24863 3511 -24807 3555
rect -24763 3511 -24707 3555
rect -24663 3511 -24607 3555
rect -24563 3511 -24507 3555
rect -24463 3511 -24407 3555
rect -24363 3511 -24307 3555
rect -24263 3511 -24207 3555
rect -24163 3511 -24107 3555
rect -24063 3511 -24007 3555
rect -23963 3511 -23907 3555
rect -23863 3511 -23407 3555
rect -23363 3511 -23307 3555
rect -23263 3511 -23207 3555
rect -23163 3511 -23107 3555
rect -23063 3511 -23007 3555
rect -22963 3511 -22907 3555
rect -22863 3511 -22807 3555
rect -22763 3511 -22707 3555
rect -22663 3511 -22607 3555
rect -22563 3511 -22507 3555
rect -22463 3511 -22407 3555
rect -22363 3511 -22307 3555
rect -22263 3511 -22207 3555
rect -22163 3511 -22107 3555
rect -22063 3511 -22007 3555
rect -21963 3511 -21907 3555
rect -21863 3511 -21407 3555
rect -21363 3511 -21307 3555
rect -21263 3511 -21207 3555
rect -21163 3511 -21107 3555
rect -21063 3511 -21007 3555
rect -20963 3511 -20907 3555
rect -20863 3511 -20807 3555
rect -20763 3511 -20707 3555
rect -20663 3511 -20607 3555
rect -20563 3511 -20507 3555
rect -20463 3511 -20407 3555
rect -20363 3511 -20307 3555
rect -20263 3511 -20207 3555
rect -20163 3511 -20107 3555
rect -20063 3511 -20007 3555
rect -19963 3511 -19907 3555
rect -19863 3511 -17010 3555
rect -30138 3455 -17010 3511
rect -30138 3411 -27407 3455
rect -27363 3411 -27307 3455
rect -27263 3411 -27207 3455
rect -27163 3411 -27107 3455
rect -27063 3411 -27007 3455
rect -26963 3411 -26907 3455
rect -26863 3411 -26807 3455
rect -26763 3411 -26707 3455
rect -26663 3411 -26607 3455
rect -26563 3411 -26507 3455
rect -26463 3411 -26407 3455
rect -26363 3411 -26307 3455
rect -26263 3411 -26207 3455
rect -26163 3411 -26107 3455
rect -26063 3411 -26007 3455
rect -25963 3411 -25907 3455
rect -25863 3411 -25407 3455
rect -25363 3411 -25307 3455
rect -25263 3411 -25207 3455
rect -25163 3411 -25107 3455
rect -25063 3411 -25007 3455
rect -24963 3411 -24907 3455
rect -24863 3411 -24807 3455
rect -24763 3411 -24707 3455
rect -24663 3411 -24607 3455
rect -24563 3411 -24507 3455
rect -24463 3411 -24407 3455
rect -24363 3411 -24307 3455
rect -24263 3411 -24207 3455
rect -24163 3411 -24107 3455
rect -24063 3411 -24007 3455
rect -23963 3411 -23907 3455
rect -23863 3411 -23407 3455
rect -23363 3411 -23307 3455
rect -23263 3411 -23207 3455
rect -23163 3411 -23107 3455
rect -23063 3411 -23007 3455
rect -22963 3411 -22907 3455
rect -22863 3411 -22807 3455
rect -22763 3411 -22707 3455
rect -22663 3411 -22607 3455
rect -22563 3411 -22507 3455
rect -22463 3411 -22407 3455
rect -22363 3411 -22307 3455
rect -22263 3411 -22207 3455
rect -22163 3411 -22107 3455
rect -22063 3411 -22007 3455
rect -21963 3411 -21907 3455
rect -21863 3411 -21407 3455
rect -21363 3411 -21307 3455
rect -21263 3411 -21207 3455
rect -21163 3411 -21107 3455
rect -21063 3411 -21007 3455
rect -20963 3411 -20907 3455
rect -20863 3411 -20807 3455
rect -20763 3411 -20707 3455
rect -20663 3411 -20607 3455
rect -20563 3411 -20507 3455
rect -20463 3411 -20407 3455
rect -20363 3411 -20307 3455
rect -20263 3411 -20207 3455
rect -20163 3411 -20107 3455
rect -20063 3411 -20007 3455
rect -19963 3411 -19907 3455
rect -19863 3411 -17010 3455
rect -30138 3355 -17010 3411
rect -30138 3311 -27407 3355
rect -27363 3311 -27307 3355
rect -27263 3311 -27207 3355
rect -27163 3311 -27107 3355
rect -27063 3311 -27007 3355
rect -26963 3311 -26907 3355
rect -26863 3311 -26807 3355
rect -26763 3311 -26707 3355
rect -26663 3311 -26607 3355
rect -26563 3311 -26507 3355
rect -26463 3311 -26407 3355
rect -26363 3311 -26307 3355
rect -26263 3311 -26207 3355
rect -26163 3311 -26107 3355
rect -26063 3311 -26007 3355
rect -25963 3311 -25907 3355
rect -25863 3311 -25407 3355
rect -25363 3311 -25307 3355
rect -25263 3311 -25207 3355
rect -25163 3311 -25107 3355
rect -25063 3311 -25007 3355
rect -24963 3311 -24907 3355
rect -24863 3311 -24807 3355
rect -24763 3311 -24707 3355
rect -24663 3311 -24607 3355
rect -24563 3311 -24507 3355
rect -24463 3311 -24407 3355
rect -24363 3311 -24307 3355
rect -24263 3311 -24207 3355
rect -24163 3311 -24107 3355
rect -24063 3311 -24007 3355
rect -23963 3311 -23907 3355
rect -23863 3311 -23407 3355
rect -23363 3311 -23307 3355
rect -23263 3311 -23207 3355
rect -23163 3311 -23107 3355
rect -23063 3311 -23007 3355
rect -22963 3311 -22907 3355
rect -22863 3311 -22807 3355
rect -22763 3311 -22707 3355
rect -22663 3311 -22607 3355
rect -22563 3311 -22507 3355
rect -22463 3311 -22407 3355
rect -22363 3311 -22307 3355
rect -22263 3311 -22207 3355
rect -22163 3311 -22107 3355
rect -22063 3311 -22007 3355
rect -21963 3311 -21907 3355
rect -21863 3311 -21407 3355
rect -21363 3311 -21307 3355
rect -21263 3311 -21207 3355
rect -21163 3311 -21107 3355
rect -21063 3311 -21007 3355
rect -20963 3311 -20907 3355
rect -20863 3311 -20807 3355
rect -20763 3311 -20707 3355
rect -20663 3311 -20607 3355
rect -20563 3311 -20507 3355
rect -20463 3311 -20407 3355
rect -20363 3311 -20307 3355
rect -20263 3311 -20207 3355
rect -20163 3311 -20107 3355
rect -20063 3311 -20007 3355
rect -19963 3311 -19907 3355
rect -19863 3311 -17010 3355
rect -30138 3255 -17010 3311
rect -30138 3211 -27407 3255
rect -27363 3211 -27307 3255
rect -27263 3211 -27207 3255
rect -27163 3211 -27107 3255
rect -27063 3211 -27007 3255
rect -26963 3211 -26907 3255
rect -26863 3211 -26807 3255
rect -26763 3211 -26707 3255
rect -26663 3211 -26607 3255
rect -26563 3211 -26507 3255
rect -26463 3211 -26407 3255
rect -26363 3211 -26307 3255
rect -26263 3211 -26207 3255
rect -26163 3211 -26107 3255
rect -26063 3211 -26007 3255
rect -25963 3211 -25907 3255
rect -25863 3211 -25407 3255
rect -25363 3211 -25307 3255
rect -25263 3211 -25207 3255
rect -25163 3211 -25107 3255
rect -25063 3211 -25007 3255
rect -24963 3211 -24907 3255
rect -24863 3211 -24807 3255
rect -24763 3211 -24707 3255
rect -24663 3211 -24607 3255
rect -24563 3211 -24507 3255
rect -24463 3211 -24407 3255
rect -24363 3211 -24307 3255
rect -24263 3211 -24207 3255
rect -24163 3211 -24107 3255
rect -24063 3211 -24007 3255
rect -23963 3211 -23907 3255
rect -23863 3211 -23407 3255
rect -23363 3211 -23307 3255
rect -23263 3211 -23207 3255
rect -23163 3211 -23107 3255
rect -23063 3211 -23007 3255
rect -22963 3211 -22907 3255
rect -22863 3211 -22807 3255
rect -22763 3211 -22707 3255
rect -22663 3211 -22607 3255
rect -22563 3211 -22507 3255
rect -22463 3211 -22407 3255
rect -22363 3211 -22307 3255
rect -22263 3211 -22207 3255
rect -22163 3211 -22107 3255
rect -22063 3211 -22007 3255
rect -21963 3211 -21907 3255
rect -21863 3211 -21407 3255
rect -21363 3211 -21307 3255
rect -21263 3211 -21207 3255
rect -21163 3211 -21107 3255
rect -21063 3211 -21007 3255
rect -20963 3211 -20907 3255
rect -20863 3211 -20807 3255
rect -20763 3211 -20707 3255
rect -20663 3211 -20607 3255
rect -20563 3211 -20507 3255
rect -20463 3211 -20407 3255
rect -20363 3211 -20307 3255
rect -20263 3211 -20207 3255
rect -20163 3211 -20107 3255
rect -20063 3211 -20007 3255
rect -19963 3211 -19907 3255
rect -19863 3211 -17010 3255
rect -30138 3155 -17010 3211
rect -30138 3111 -27407 3155
rect -27363 3111 -27307 3155
rect -27263 3111 -27207 3155
rect -27163 3111 -27107 3155
rect -27063 3111 -27007 3155
rect -26963 3111 -26907 3155
rect -26863 3111 -26807 3155
rect -26763 3111 -26707 3155
rect -26663 3111 -26607 3155
rect -26563 3111 -26507 3155
rect -26463 3111 -26407 3155
rect -26363 3111 -26307 3155
rect -26263 3111 -26207 3155
rect -26163 3111 -26107 3155
rect -26063 3111 -26007 3155
rect -25963 3111 -25907 3155
rect -25863 3111 -25407 3155
rect -25363 3111 -25307 3155
rect -25263 3111 -25207 3155
rect -25163 3111 -25107 3155
rect -25063 3111 -25007 3155
rect -24963 3111 -24907 3155
rect -24863 3111 -24807 3155
rect -24763 3111 -24707 3155
rect -24663 3111 -24607 3155
rect -24563 3111 -24507 3155
rect -24463 3111 -24407 3155
rect -24363 3111 -24307 3155
rect -24263 3111 -24207 3155
rect -24163 3111 -24107 3155
rect -24063 3111 -24007 3155
rect -23963 3111 -23907 3155
rect -23863 3111 -23407 3155
rect -23363 3111 -23307 3155
rect -23263 3111 -23207 3155
rect -23163 3111 -23107 3155
rect -23063 3111 -23007 3155
rect -22963 3111 -22907 3155
rect -22863 3111 -22807 3155
rect -22763 3111 -22707 3155
rect -22663 3111 -22607 3155
rect -22563 3111 -22507 3155
rect -22463 3111 -22407 3155
rect -22363 3111 -22307 3155
rect -22263 3111 -22207 3155
rect -22163 3111 -22107 3155
rect -22063 3111 -22007 3155
rect -21963 3111 -21907 3155
rect -21863 3111 -21407 3155
rect -21363 3111 -21307 3155
rect -21263 3111 -21207 3155
rect -21163 3111 -21107 3155
rect -21063 3111 -21007 3155
rect -20963 3111 -20907 3155
rect -20863 3111 -20807 3155
rect -20763 3111 -20707 3155
rect -20663 3111 -20607 3155
rect -20563 3111 -20507 3155
rect -20463 3111 -20407 3155
rect -20363 3111 -20307 3155
rect -20263 3111 -20207 3155
rect -20163 3111 -20107 3155
rect -20063 3111 -20007 3155
rect -19963 3111 -19907 3155
rect -19863 3111 -17010 3155
rect -30138 3055 -17010 3111
rect -30138 3011 -27407 3055
rect -27363 3011 -27307 3055
rect -27263 3011 -27207 3055
rect -27163 3011 -27107 3055
rect -27063 3011 -27007 3055
rect -26963 3011 -26907 3055
rect -26863 3011 -26807 3055
rect -26763 3011 -26707 3055
rect -26663 3011 -26607 3055
rect -26563 3011 -26507 3055
rect -26463 3011 -26407 3055
rect -26363 3011 -26307 3055
rect -26263 3011 -26207 3055
rect -26163 3011 -26107 3055
rect -26063 3011 -26007 3055
rect -25963 3011 -25907 3055
rect -25863 3011 -25407 3055
rect -25363 3011 -25307 3055
rect -25263 3011 -25207 3055
rect -25163 3011 -25107 3055
rect -25063 3011 -25007 3055
rect -24963 3011 -24907 3055
rect -24863 3011 -24807 3055
rect -24763 3011 -24707 3055
rect -24663 3011 -24607 3055
rect -24563 3011 -24507 3055
rect -24463 3011 -24407 3055
rect -24363 3011 -24307 3055
rect -24263 3011 -24207 3055
rect -24163 3011 -24107 3055
rect -24063 3011 -24007 3055
rect -23963 3011 -23907 3055
rect -23863 3011 -23407 3055
rect -23363 3011 -23307 3055
rect -23263 3011 -23207 3055
rect -23163 3011 -23107 3055
rect -23063 3011 -23007 3055
rect -22963 3011 -22907 3055
rect -22863 3011 -22807 3055
rect -22763 3011 -22707 3055
rect -22663 3011 -22607 3055
rect -22563 3011 -22507 3055
rect -22463 3011 -22407 3055
rect -22363 3011 -22307 3055
rect -22263 3011 -22207 3055
rect -22163 3011 -22107 3055
rect -22063 3011 -22007 3055
rect -21963 3011 -21907 3055
rect -21863 3011 -21407 3055
rect -21363 3011 -21307 3055
rect -21263 3011 -21207 3055
rect -21163 3011 -21107 3055
rect -21063 3011 -21007 3055
rect -20963 3011 -20907 3055
rect -20863 3011 -20807 3055
rect -20763 3011 -20707 3055
rect -20663 3011 -20607 3055
rect -20563 3011 -20507 3055
rect -20463 3011 -20407 3055
rect -20363 3011 -20307 3055
rect -20263 3011 -20207 3055
rect -20163 3011 -20107 3055
rect -20063 3011 -20007 3055
rect -19963 3011 -19907 3055
rect -19863 3011 -17010 3055
rect -30138 2955 -17010 3011
rect -30138 2911 -27407 2955
rect -27363 2911 -27307 2955
rect -27263 2911 -27207 2955
rect -27163 2911 -27107 2955
rect -27063 2911 -27007 2955
rect -26963 2911 -26907 2955
rect -26863 2911 -26807 2955
rect -26763 2911 -26707 2955
rect -26663 2911 -26607 2955
rect -26563 2911 -26507 2955
rect -26463 2911 -26407 2955
rect -26363 2911 -26307 2955
rect -26263 2911 -26207 2955
rect -26163 2911 -26107 2955
rect -26063 2911 -26007 2955
rect -25963 2911 -25907 2955
rect -25863 2911 -25407 2955
rect -25363 2911 -25307 2955
rect -25263 2911 -25207 2955
rect -25163 2911 -25107 2955
rect -25063 2911 -25007 2955
rect -24963 2911 -24907 2955
rect -24863 2911 -24807 2955
rect -24763 2911 -24707 2955
rect -24663 2911 -24607 2955
rect -24563 2911 -24507 2955
rect -24463 2911 -24407 2955
rect -24363 2911 -24307 2955
rect -24263 2911 -24207 2955
rect -24163 2911 -24107 2955
rect -24063 2911 -24007 2955
rect -23963 2911 -23907 2955
rect -23863 2911 -23407 2955
rect -23363 2911 -23307 2955
rect -23263 2911 -23207 2955
rect -23163 2911 -23107 2955
rect -23063 2911 -23007 2955
rect -22963 2911 -22907 2955
rect -22863 2911 -22807 2955
rect -22763 2911 -22707 2955
rect -22663 2911 -22607 2955
rect -22563 2911 -22507 2955
rect -22463 2911 -22407 2955
rect -22363 2911 -22307 2955
rect -22263 2911 -22207 2955
rect -22163 2911 -22107 2955
rect -22063 2911 -22007 2955
rect -21963 2911 -21907 2955
rect -21863 2911 -21407 2955
rect -21363 2911 -21307 2955
rect -21263 2911 -21207 2955
rect -21163 2911 -21107 2955
rect -21063 2911 -21007 2955
rect -20963 2911 -20907 2955
rect -20863 2911 -20807 2955
rect -20763 2911 -20707 2955
rect -20663 2911 -20607 2955
rect -20563 2911 -20507 2955
rect -20463 2911 -20407 2955
rect -20363 2911 -20307 2955
rect -20263 2911 -20207 2955
rect -20163 2911 -20107 2955
rect -20063 2911 -20007 2955
rect -19963 2911 -19907 2955
rect -19863 2911 -17010 2955
rect -30138 2855 -17010 2911
rect -30138 2811 -27407 2855
rect -27363 2811 -27307 2855
rect -27263 2811 -27207 2855
rect -27163 2811 -27107 2855
rect -27063 2811 -27007 2855
rect -26963 2811 -26907 2855
rect -26863 2811 -26807 2855
rect -26763 2811 -26707 2855
rect -26663 2811 -26607 2855
rect -26563 2811 -26507 2855
rect -26463 2811 -26407 2855
rect -26363 2811 -26307 2855
rect -26263 2811 -26207 2855
rect -26163 2811 -26107 2855
rect -26063 2811 -26007 2855
rect -25963 2811 -25907 2855
rect -25863 2811 -25407 2855
rect -25363 2811 -25307 2855
rect -25263 2811 -25207 2855
rect -25163 2811 -25107 2855
rect -25063 2811 -25007 2855
rect -24963 2811 -24907 2855
rect -24863 2811 -24807 2855
rect -24763 2811 -24707 2855
rect -24663 2811 -24607 2855
rect -24563 2811 -24507 2855
rect -24463 2811 -24407 2855
rect -24363 2811 -24307 2855
rect -24263 2811 -24207 2855
rect -24163 2811 -24107 2855
rect -24063 2811 -24007 2855
rect -23963 2811 -23907 2855
rect -23863 2811 -23407 2855
rect -23363 2811 -23307 2855
rect -23263 2811 -23207 2855
rect -23163 2811 -23107 2855
rect -23063 2811 -23007 2855
rect -22963 2811 -22907 2855
rect -22863 2811 -22807 2855
rect -22763 2811 -22707 2855
rect -22663 2811 -22607 2855
rect -22563 2811 -22507 2855
rect -22463 2811 -22407 2855
rect -22363 2811 -22307 2855
rect -22263 2811 -22207 2855
rect -22163 2811 -22107 2855
rect -22063 2811 -22007 2855
rect -21963 2811 -21907 2855
rect -21863 2811 -21407 2855
rect -21363 2811 -21307 2855
rect -21263 2811 -21207 2855
rect -21163 2811 -21107 2855
rect -21063 2811 -21007 2855
rect -20963 2811 -20907 2855
rect -20863 2811 -20807 2855
rect -20763 2811 -20707 2855
rect -20663 2811 -20607 2855
rect -20563 2811 -20507 2855
rect -20463 2811 -20407 2855
rect -20363 2811 -20307 2855
rect -20263 2811 -20207 2855
rect -20163 2811 -20107 2855
rect -20063 2811 -20007 2855
rect -19963 2811 -19907 2855
rect -19863 2811 -17010 2855
rect -30138 2755 -17010 2811
rect -30138 2711 -27407 2755
rect -27363 2711 -27307 2755
rect -27263 2711 -27207 2755
rect -27163 2711 -27107 2755
rect -27063 2711 -27007 2755
rect -26963 2711 -26907 2755
rect -26863 2711 -26807 2755
rect -26763 2711 -26707 2755
rect -26663 2711 -26607 2755
rect -26563 2711 -26507 2755
rect -26463 2711 -26407 2755
rect -26363 2711 -26307 2755
rect -26263 2711 -26207 2755
rect -26163 2711 -26107 2755
rect -26063 2711 -26007 2755
rect -25963 2711 -25907 2755
rect -25863 2711 -25407 2755
rect -25363 2711 -25307 2755
rect -25263 2711 -25207 2755
rect -25163 2711 -25107 2755
rect -25063 2711 -25007 2755
rect -24963 2711 -24907 2755
rect -24863 2711 -24807 2755
rect -24763 2711 -24707 2755
rect -24663 2711 -24607 2755
rect -24563 2711 -24507 2755
rect -24463 2711 -24407 2755
rect -24363 2711 -24307 2755
rect -24263 2711 -24207 2755
rect -24163 2711 -24107 2755
rect -24063 2711 -24007 2755
rect -23963 2711 -23907 2755
rect -23863 2711 -23407 2755
rect -23363 2711 -23307 2755
rect -23263 2711 -23207 2755
rect -23163 2711 -23107 2755
rect -23063 2711 -23007 2755
rect -22963 2711 -22907 2755
rect -22863 2711 -22807 2755
rect -22763 2711 -22707 2755
rect -22663 2711 -22607 2755
rect -22563 2711 -22507 2755
rect -22463 2711 -22407 2755
rect -22363 2711 -22307 2755
rect -22263 2711 -22207 2755
rect -22163 2711 -22107 2755
rect -22063 2711 -22007 2755
rect -21963 2711 -21907 2755
rect -21863 2711 -21407 2755
rect -21363 2711 -21307 2755
rect -21263 2711 -21207 2755
rect -21163 2711 -21107 2755
rect -21063 2711 -21007 2755
rect -20963 2711 -20907 2755
rect -20863 2711 -20807 2755
rect -20763 2711 -20707 2755
rect -20663 2711 -20607 2755
rect -20563 2711 -20507 2755
rect -20463 2711 -20407 2755
rect -20363 2711 -20307 2755
rect -20263 2711 -20207 2755
rect -20163 2711 -20107 2755
rect -20063 2711 -20007 2755
rect -19963 2711 -19907 2755
rect -19863 2711 -17010 2755
rect -30138 2655 -17010 2711
rect -6280 2655 -5369 6068
rect -30138 2611 -27407 2655
rect -27363 2611 -27307 2655
rect -27263 2611 -27207 2655
rect -27163 2611 -27107 2655
rect -27063 2611 -27007 2655
rect -26963 2611 -26907 2655
rect -26863 2611 -26807 2655
rect -26763 2611 -26707 2655
rect -26663 2611 -26607 2655
rect -26563 2611 -26507 2655
rect -26463 2611 -26407 2655
rect -26363 2611 -26307 2655
rect -26263 2611 -26207 2655
rect -26163 2611 -26107 2655
rect -26063 2611 -26007 2655
rect -25963 2611 -25907 2655
rect -25863 2611 -25407 2655
rect -25363 2611 -25307 2655
rect -25263 2611 -25207 2655
rect -25163 2611 -25107 2655
rect -25063 2611 -25007 2655
rect -24963 2611 -24907 2655
rect -24863 2611 -24807 2655
rect -24763 2611 -24707 2655
rect -24663 2611 -24607 2655
rect -24563 2611 -24507 2655
rect -24463 2611 -24407 2655
rect -24363 2611 -24307 2655
rect -24263 2611 -24207 2655
rect -24163 2611 -24107 2655
rect -24063 2611 -24007 2655
rect -23963 2611 -23907 2655
rect -23863 2611 -23407 2655
rect -23363 2611 -23307 2655
rect -23263 2611 -23207 2655
rect -23163 2611 -23107 2655
rect -23063 2611 -23007 2655
rect -22963 2611 -22907 2655
rect -22863 2611 -22807 2655
rect -22763 2611 -22707 2655
rect -22663 2611 -22607 2655
rect -22563 2611 -22507 2655
rect -22463 2611 -22407 2655
rect -22363 2611 -22307 2655
rect -22263 2611 -22207 2655
rect -22163 2611 -22107 2655
rect -22063 2611 -22007 2655
rect -21963 2611 -21907 2655
rect -21863 2611 -21407 2655
rect -21363 2611 -21307 2655
rect -21263 2611 -21207 2655
rect -21163 2611 -21107 2655
rect -21063 2611 -21007 2655
rect -20963 2611 -20907 2655
rect -20863 2611 -20807 2655
rect -20763 2611 -20707 2655
rect -20663 2611 -20607 2655
rect -20563 2611 -20507 2655
rect -20463 2611 -20407 2655
rect -20363 2611 -20307 2655
rect -20263 2611 -20207 2655
rect -20163 2611 -20107 2655
rect -20063 2611 -20007 2655
rect -19963 2611 -19907 2655
rect -19863 2611 -5369 2655
rect -30138 2555 -5369 2611
rect -30138 2511 -27407 2555
rect -27363 2511 -27307 2555
rect -27263 2511 -27207 2555
rect -27163 2511 -27107 2555
rect -27063 2511 -27007 2555
rect -26963 2511 -26907 2555
rect -26863 2511 -26807 2555
rect -26763 2511 -26707 2555
rect -26663 2511 -26607 2555
rect -26563 2511 -26507 2555
rect -26463 2511 -26407 2555
rect -26363 2511 -26307 2555
rect -26263 2511 -26207 2555
rect -26163 2511 -26107 2555
rect -26063 2511 -26007 2555
rect -25963 2511 -25907 2555
rect -25863 2511 -25407 2555
rect -25363 2511 -25307 2555
rect -25263 2511 -25207 2555
rect -25163 2511 -25107 2555
rect -25063 2511 -25007 2555
rect -24963 2511 -24907 2555
rect -24863 2511 -24807 2555
rect -24763 2511 -24707 2555
rect -24663 2511 -24607 2555
rect -24563 2511 -24507 2555
rect -24463 2511 -24407 2555
rect -24363 2511 -24307 2555
rect -24263 2511 -24207 2555
rect -24163 2511 -24107 2555
rect -24063 2511 -24007 2555
rect -23963 2511 -23907 2555
rect -23863 2511 -23407 2555
rect -23363 2511 -23307 2555
rect -23263 2511 -23207 2555
rect -23163 2511 -23107 2555
rect -23063 2511 -23007 2555
rect -22963 2511 -22907 2555
rect -22863 2511 -22807 2555
rect -22763 2511 -22707 2555
rect -22663 2511 -22607 2555
rect -22563 2511 -22507 2555
rect -22463 2511 -22407 2555
rect -22363 2511 -22307 2555
rect -22263 2511 -22207 2555
rect -22163 2511 -22107 2555
rect -22063 2511 -22007 2555
rect -21963 2511 -21907 2555
rect -21863 2511 -21407 2555
rect -21363 2511 -21307 2555
rect -21263 2511 -21207 2555
rect -21163 2511 -21107 2555
rect -21063 2511 -21007 2555
rect -20963 2511 -20907 2555
rect -20863 2511 -20807 2555
rect -20763 2511 -20707 2555
rect -20663 2511 -20607 2555
rect -20563 2511 -20507 2555
rect -20463 2511 -20407 2555
rect -20363 2511 -20307 2555
rect -20263 2511 -20207 2555
rect -20163 2511 -20107 2555
rect -20063 2511 -20007 2555
rect -19963 2511 -19907 2555
rect -19863 2511 -5369 2555
rect -30138 2455 -5369 2511
rect -30138 2411 -27407 2455
rect -27363 2411 -27307 2455
rect -27263 2411 -27207 2455
rect -27163 2411 -27107 2455
rect -27063 2411 -27007 2455
rect -26963 2411 -26907 2455
rect -26863 2411 -26807 2455
rect -26763 2411 -26707 2455
rect -26663 2411 -26607 2455
rect -26563 2411 -26507 2455
rect -26463 2411 -26407 2455
rect -26363 2411 -26307 2455
rect -26263 2411 -26207 2455
rect -26163 2411 -26107 2455
rect -26063 2411 -26007 2455
rect -25963 2411 -25907 2455
rect -25863 2411 -25407 2455
rect -25363 2411 -25307 2455
rect -25263 2411 -25207 2455
rect -25163 2411 -25107 2455
rect -25063 2411 -25007 2455
rect -24963 2411 -24907 2455
rect -24863 2411 -24807 2455
rect -24763 2411 -24707 2455
rect -24663 2411 -24607 2455
rect -24563 2411 -24507 2455
rect -24463 2411 -24407 2455
rect -24363 2411 -24307 2455
rect -24263 2411 -24207 2455
rect -24163 2411 -24107 2455
rect -24063 2411 -24007 2455
rect -23963 2411 -23907 2455
rect -23863 2411 -23407 2455
rect -23363 2411 -23307 2455
rect -23263 2411 -23207 2455
rect -23163 2411 -23107 2455
rect -23063 2411 -23007 2455
rect -22963 2411 -22907 2455
rect -22863 2411 -22807 2455
rect -22763 2411 -22707 2455
rect -22663 2411 -22607 2455
rect -22563 2411 -22507 2455
rect -22463 2411 -22407 2455
rect -22363 2411 -22307 2455
rect -22263 2411 -22207 2455
rect -22163 2411 -22107 2455
rect -22063 2411 -22007 2455
rect -21963 2411 -21907 2455
rect -21863 2411 -21407 2455
rect -21363 2411 -21307 2455
rect -21263 2411 -21207 2455
rect -21163 2411 -21107 2455
rect -21063 2411 -21007 2455
rect -20963 2411 -20907 2455
rect -20863 2411 -20807 2455
rect -20763 2411 -20707 2455
rect -20663 2411 -20607 2455
rect -20563 2411 -20507 2455
rect -20463 2411 -20407 2455
rect -20363 2411 -20307 2455
rect -20263 2411 -20207 2455
rect -20163 2411 -20107 2455
rect -20063 2411 -20007 2455
rect -19963 2411 -19907 2455
rect -19863 2411 -5369 2455
rect -30138 2355 -5369 2411
rect -30138 2311 -27407 2355
rect -27363 2311 -27307 2355
rect -27263 2311 -27207 2355
rect -27163 2311 -27107 2355
rect -27063 2311 -27007 2355
rect -26963 2311 -26907 2355
rect -26863 2311 -26807 2355
rect -26763 2311 -26707 2355
rect -26663 2311 -26607 2355
rect -26563 2311 -26507 2355
rect -26463 2311 -26407 2355
rect -26363 2311 -26307 2355
rect -26263 2311 -26207 2355
rect -26163 2311 -26107 2355
rect -26063 2311 -26007 2355
rect -25963 2311 -25907 2355
rect -25863 2311 -25407 2355
rect -25363 2311 -25307 2355
rect -25263 2311 -25207 2355
rect -25163 2311 -25107 2355
rect -25063 2311 -25007 2355
rect -24963 2311 -24907 2355
rect -24863 2311 -24807 2355
rect -24763 2311 -24707 2355
rect -24663 2311 -24607 2355
rect -24563 2311 -24507 2355
rect -24463 2311 -24407 2355
rect -24363 2311 -24307 2355
rect -24263 2311 -24207 2355
rect -24163 2311 -24107 2355
rect -24063 2311 -24007 2355
rect -23963 2311 -23907 2355
rect -23863 2311 -23407 2355
rect -23363 2311 -23307 2355
rect -23263 2311 -23207 2355
rect -23163 2311 -23107 2355
rect -23063 2311 -23007 2355
rect -22963 2311 -22907 2355
rect -22863 2311 -22807 2355
rect -22763 2311 -22707 2355
rect -22663 2311 -22607 2355
rect -22563 2311 -22507 2355
rect -22463 2311 -22407 2355
rect -22363 2311 -22307 2355
rect -22263 2311 -22207 2355
rect -22163 2311 -22107 2355
rect -22063 2311 -22007 2355
rect -21963 2311 -21907 2355
rect -21863 2311 -21407 2355
rect -21363 2311 -21307 2355
rect -21263 2311 -21207 2355
rect -21163 2311 -21107 2355
rect -21063 2311 -21007 2355
rect -20963 2311 -20907 2355
rect -20863 2311 -20807 2355
rect -20763 2311 -20707 2355
rect -20663 2311 -20607 2355
rect -20563 2311 -20507 2355
rect -20463 2311 -20407 2355
rect -20363 2311 -20307 2355
rect -20263 2311 -20207 2355
rect -20163 2311 -20107 2355
rect -20063 2311 -20007 2355
rect -19963 2311 -19907 2355
rect -19863 2311 -5369 2355
rect -30138 2255 -5369 2311
rect -30138 2211 -27407 2255
rect -27363 2211 -27307 2255
rect -27263 2211 -27207 2255
rect -27163 2211 -27107 2255
rect -27063 2211 -27007 2255
rect -26963 2211 -26907 2255
rect -26863 2211 -26807 2255
rect -26763 2211 -26707 2255
rect -26663 2211 -26607 2255
rect -26563 2211 -26507 2255
rect -26463 2211 -26407 2255
rect -26363 2211 -26307 2255
rect -26263 2211 -26207 2255
rect -26163 2211 -26107 2255
rect -26063 2211 -26007 2255
rect -25963 2211 -25907 2255
rect -25863 2211 -25407 2255
rect -25363 2211 -25307 2255
rect -25263 2211 -25207 2255
rect -25163 2211 -25107 2255
rect -25063 2211 -25007 2255
rect -24963 2211 -24907 2255
rect -24863 2211 -24807 2255
rect -24763 2211 -24707 2255
rect -24663 2211 -24607 2255
rect -24563 2211 -24507 2255
rect -24463 2211 -24407 2255
rect -24363 2211 -24307 2255
rect -24263 2211 -24207 2255
rect -24163 2211 -24107 2255
rect -24063 2211 -24007 2255
rect -23963 2211 -23907 2255
rect -23863 2211 -23407 2255
rect -23363 2211 -23307 2255
rect -23263 2211 -23207 2255
rect -23163 2211 -23107 2255
rect -23063 2211 -23007 2255
rect -22963 2211 -22907 2255
rect -22863 2211 -22807 2255
rect -22763 2211 -22707 2255
rect -22663 2211 -22607 2255
rect -22563 2211 -22507 2255
rect -22463 2211 -22407 2255
rect -22363 2211 -22307 2255
rect -22263 2211 -22207 2255
rect -22163 2211 -22107 2255
rect -22063 2211 -22007 2255
rect -21963 2211 -21907 2255
rect -21863 2211 -21407 2255
rect -21363 2211 -21307 2255
rect -21263 2211 -21207 2255
rect -21163 2211 -21107 2255
rect -21063 2211 -21007 2255
rect -20963 2211 -20907 2255
rect -20863 2211 -20807 2255
rect -20763 2211 -20707 2255
rect -20663 2211 -20607 2255
rect -20563 2211 -20507 2255
rect -20463 2211 -20407 2255
rect -20363 2211 -20307 2255
rect -20263 2211 -20207 2255
rect -20163 2211 -20107 2255
rect -20063 2211 -20007 2255
rect -19963 2211 -19907 2255
rect -19863 2211 -5369 2255
rect -30138 2155 -5369 2211
rect -30138 2111 -27407 2155
rect -27363 2111 -27307 2155
rect -27263 2111 -27207 2155
rect -27163 2111 -27107 2155
rect -27063 2111 -27007 2155
rect -26963 2111 -26907 2155
rect -26863 2111 -26807 2155
rect -26763 2111 -26707 2155
rect -26663 2111 -26607 2155
rect -26563 2111 -26507 2155
rect -26463 2111 -26407 2155
rect -26363 2111 -26307 2155
rect -26263 2111 -26207 2155
rect -26163 2111 -26107 2155
rect -26063 2111 -26007 2155
rect -25963 2111 -25907 2155
rect -25863 2111 -25407 2155
rect -25363 2111 -25307 2155
rect -25263 2111 -25207 2155
rect -25163 2111 -25107 2155
rect -25063 2111 -25007 2155
rect -24963 2111 -24907 2155
rect -24863 2111 -24807 2155
rect -24763 2111 -24707 2155
rect -24663 2111 -24607 2155
rect -24563 2111 -24507 2155
rect -24463 2111 -24407 2155
rect -24363 2111 -24307 2155
rect -24263 2111 -24207 2155
rect -24163 2111 -24107 2155
rect -24063 2111 -24007 2155
rect -23963 2111 -23907 2155
rect -23863 2111 -23407 2155
rect -23363 2111 -23307 2155
rect -23263 2111 -23207 2155
rect -23163 2111 -23107 2155
rect -23063 2111 -23007 2155
rect -22963 2111 -22907 2155
rect -22863 2111 -22807 2155
rect -22763 2111 -22707 2155
rect -22663 2111 -22607 2155
rect -22563 2111 -22507 2155
rect -22463 2111 -22407 2155
rect -22363 2111 -22307 2155
rect -22263 2111 -22207 2155
rect -22163 2111 -22107 2155
rect -22063 2111 -22007 2155
rect -21963 2111 -21907 2155
rect -21863 2111 -21407 2155
rect -21363 2111 -21307 2155
rect -21263 2111 -21207 2155
rect -21163 2111 -21107 2155
rect -21063 2111 -21007 2155
rect -20963 2111 -20907 2155
rect -20863 2111 -20807 2155
rect -20763 2111 -20707 2155
rect -20663 2111 -20607 2155
rect -20563 2111 -20507 2155
rect -20463 2111 -20407 2155
rect -20363 2111 -20307 2155
rect -20263 2111 -20207 2155
rect -20163 2111 -20107 2155
rect -20063 2111 -20007 2155
rect -19963 2111 -19907 2155
rect -19863 2111 -5369 2155
rect -30138 2055 -5369 2111
rect -30138 2011 -27407 2055
rect -27363 2011 -27307 2055
rect -27263 2011 -27207 2055
rect -27163 2011 -27107 2055
rect -27063 2011 -27007 2055
rect -26963 2011 -26907 2055
rect -26863 2011 -26807 2055
rect -26763 2011 -26707 2055
rect -26663 2011 -26607 2055
rect -26563 2011 -26507 2055
rect -26463 2011 -26407 2055
rect -26363 2011 -26307 2055
rect -26263 2011 -26207 2055
rect -26163 2011 -26107 2055
rect -26063 2011 -26007 2055
rect -25963 2011 -25907 2055
rect -25863 2011 -25407 2055
rect -25363 2011 -25307 2055
rect -25263 2011 -25207 2055
rect -25163 2011 -25107 2055
rect -25063 2011 -25007 2055
rect -24963 2011 -24907 2055
rect -24863 2011 -24807 2055
rect -24763 2011 -24707 2055
rect -24663 2011 -24607 2055
rect -24563 2011 -24507 2055
rect -24463 2011 -24407 2055
rect -24363 2011 -24307 2055
rect -24263 2011 -24207 2055
rect -24163 2011 -24107 2055
rect -24063 2011 -24007 2055
rect -23963 2011 -23907 2055
rect -23863 2011 -23407 2055
rect -23363 2011 -23307 2055
rect -23263 2011 -23207 2055
rect -23163 2011 -23107 2055
rect -23063 2011 -23007 2055
rect -22963 2011 -22907 2055
rect -22863 2011 -22807 2055
rect -22763 2011 -22707 2055
rect -22663 2011 -22607 2055
rect -22563 2011 -22507 2055
rect -22463 2011 -22407 2055
rect -22363 2011 -22307 2055
rect -22263 2011 -22207 2055
rect -22163 2011 -22107 2055
rect -22063 2011 -22007 2055
rect -21963 2011 -21907 2055
rect -21863 2011 -21407 2055
rect -21363 2011 -21307 2055
rect -21263 2011 -21207 2055
rect -21163 2011 -21107 2055
rect -21063 2011 -21007 2055
rect -20963 2011 -20907 2055
rect -20863 2011 -20807 2055
rect -20763 2011 -20707 2055
rect -20663 2011 -20607 2055
rect -20563 2011 -20507 2055
rect -20463 2011 -20407 2055
rect -20363 2011 -20307 2055
rect -20263 2011 -20207 2055
rect -20163 2011 -20107 2055
rect -20063 2011 -20007 2055
rect -19963 2011 -19907 2055
rect -19863 2011 -5369 2055
rect -30138 878 -5369 2011
rect -30138 -263 -17010 878
rect -266 -48 -32 9954
rect 27734 -48 27968 9954
rect 53672 3509 55820 3752
rect 53672 2563 55404 3509
rect 55450 2563 55820 3509
rect 396 -770 472 -48
rect 1404 -770 1480 -48
rect 2412 -770 2488 -48
rect 3420 -770 3496 -48
rect 4428 -770 4504 -48
rect 5436 -770 5512 -48
rect 6444 -770 6520 -48
rect 7452 -770 7528 -48
rect 8460 -770 8536 -48
rect 9468 -770 9544 -48
rect 10476 -770 10552 -48
rect 11484 -770 11560 -48
rect 12492 -770 12568 -48
rect 13500 -770 13576 -48
rect 14508 -770 14584 -48
rect 15516 -770 15592 -48
rect 16524 -770 16600 -48
rect 17532 -770 17608 -48
rect 18540 -770 18616 -48
rect 19548 -770 19624 -48
rect 20556 -770 20632 -48
rect 21564 -770 21640 -48
rect 22572 -770 22648 -48
rect 23580 -770 23656 -48
rect 24588 -770 24664 -48
rect 28396 -770 28472 -48
rect 29404 -770 29480 -48
rect 30412 -770 30488 -48
rect 31420 -770 31496 -48
rect 32428 -770 32504 -48
rect 33436 -770 33512 -48
rect 34444 -770 34520 -48
rect 35452 -770 35528 -48
rect 36460 -770 36536 -48
rect 37468 -770 37544 -48
rect 38476 -770 38552 -48
rect 39484 -770 39560 -48
rect 40492 -770 40568 -48
rect 41500 -770 41576 -48
rect 42508 -770 42584 -48
rect 43516 -770 43592 -48
rect 44524 -770 44600 -48
rect 45532 -770 45608 -48
rect 46540 -770 46616 -48
rect 47548 -770 47624 -48
rect 48556 -770 48632 -48
rect 49564 -770 49640 -48
rect 50572 -770 50648 -48
rect 51580 -770 51656 -48
rect 52588 -770 52664 -48
rect 53672 -770 55820 2563
rect 396 -970 25672 -770
rect 396 -1016 2307 -970
rect 22253 -1016 25672 -970
rect -14328 -6876 -4908 -6646
rect -14328 -7230 -14098 -6876
rect -14328 -7452 -14324 -7230
rect -14102 -7452 -14098 -7230
rect -14328 -7700 -14098 -7452
rect -13583 -7154 -5653 -7078
rect -13583 -7374 -12772 -7154
rect -12552 -7374 -12302 -7154
rect -12082 -7374 -11832 -7154
rect -11612 -7374 -11362 -7154
rect -11142 -7374 -10892 -7154
rect -10672 -7374 -10422 -7154
rect -10202 -7374 -9952 -7154
rect -9732 -7374 -9482 -7154
rect -9262 -7374 -9012 -7154
rect -8792 -7374 -8542 -7154
rect -8322 -7374 -8072 -7154
rect -7852 -7374 -7602 -7154
rect -7382 -7374 -7132 -7154
rect -6912 -7374 -6662 -7154
rect -6442 -7374 -5653 -7154
rect -13583 -7450 -5653 -7374
rect -13583 -7672 -13489 -7450
rect -13267 -7672 -13019 -7450
rect -12797 -7672 -12549 -7450
rect -12327 -7672 -12079 -7450
rect -11857 -7672 -11609 -7450
rect -11387 -7672 -11139 -7450
rect -10917 -7672 -10669 -7450
rect -10447 -7672 -10199 -7450
rect -9977 -7672 -9729 -7450
rect -9507 -7672 -9259 -7450
rect -9037 -7672 -8789 -7450
rect -8567 -7672 -8319 -7450
rect -8097 -7672 -7849 -7450
rect -7627 -7672 -7379 -7450
rect -7157 -7672 -6909 -7450
rect -6687 -7672 -6439 -7450
rect -6217 -7672 -5969 -7450
rect -5747 -7672 -5653 -7450
rect -13583 -7676 -5653 -7672
rect -5138 -7230 -4908 -6876
rect -5138 -7452 -5134 -7230
rect -4912 -7452 -4908 -7230
rect -14328 -7922 -14324 -7700
rect -14102 -7922 -14098 -7700
rect -14328 -8170 -14098 -7922
rect -14328 -8392 -14324 -8170
rect -14102 -8392 -14098 -8170
rect -14328 -8640 -14098 -8392
rect -14328 -8862 -14324 -8640
rect -14102 -8862 -14098 -8640
rect -14328 -9110 -14098 -8862
rect -14328 -9332 -14324 -9110
rect -14102 -9332 -14098 -9110
rect -14328 -9580 -14098 -9332
rect -14328 -9802 -14324 -9580
rect -14102 -9802 -14098 -9580
rect -14328 -10050 -14098 -9802
rect -14328 -10272 -14324 -10050
rect -14102 -10272 -14098 -10050
rect -14328 -10520 -14098 -10272
rect -14328 -10742 -14324 -10520
rect -14102 -10742 -14098 -10520
rect -14328 -10990 -14098 -10742
rect -14328 -11212 -14324 -10990
rect -14102 -11212 -14098 -10990
rect -14328 -11460 -14098 -11212
rect -14328 -11682 -14324 -11460
rect -14102 -11682 -14098 -11460
rect -14328 -11930 -14098 -11682
rect -14328 -12152 -14324 -11930
rect -14102 -12152 -14098 -11930
rect -14328 -12400 -14098 -12152
rect -14328 -12622 -14324 -12400
rect -14102 -12622 -14098 -12400
rect -14328 -12870 -14098 -12622
rect -14328 -13092 -14324 -12870
rect -14102 -13092 -14098 -12870
rect -14328 -13340 -14098 -13092
rect -5138 -7700 -4908 -7452
rect -5138 -7922 -5134 -7700
rect -4912 -7922 -4908 -7700
rect -5138 -8170 -4908 -7922
rect -5138 -8392 -5134 -8170
rect -4912 -8392 -4908 -8170
rect -5138 -8640 -4908 -8392
rect -5138 -8862 -5134 -8640
rect -4912 -8862 -4908 -8640
rect -5138 -9110 -4908 -8862
rect -5138 -9332 -5134 -9110
rect -4912 -9332 -4908 -9110
rect -5138 -9580 -4908 -9332
rect -5138 -9802 -5134 -9580
rect -4912 -9802 -4908 -9580
rect -5138 -10050 -4908 -9802
rect -5138 -10272 -5134 -10050
rect -4912 -10272 -4908 -10050
rect -5138 -10520 -4908 -10272
rect -5138 -10742 -5134 -10520
rect -4912 -10742 -4908 -10520
rect -5138 -10990 -4908 -10742
rect -5138 -11212 -5134 -10990
rect -4912 -11212 -4908 -10990
rect -5138 -11460 -4908 -11212
rect -5138 -11682 -5134 -11460
rect -4912 -11682 -4908 -11460
rect -5138 -11930 -4908 -11682
rect -5138 -12152 -5134 -11930
rect -4912 -12152 -4908 -11930
rect -5138 -12400 -4908 -12152
rect -5138 -12622 -5134 -12400
rect -4912 -12622 -4908 -12400
rect -5138 -12870 -4908 -12622
rect -5138 -13092 -5134 -12870
rect -4912 -13092 -4908 -12870
rect -14328 -13562 -14324 -13340
rect -14102 -13562 -14098 -13340
rect -14328 -13916 -14098 -13562
rect -13583 -13120 -5653 -13116
rect -13583 -13342 -13489 -13120
rect -13267 -13342 -13019 -13120
rect -12797 -13342 -12549 -13120
rect -12327 -13342 -12079 -13120
rect -11857 -13342 -11609 -13120
rect -11387 -13342 -11139 -13120
rect -10917 -13342 -10669 -13120
rect -10447 -13342 -10199 -13120
rect -9977 -13342 -9729 -13120
rect -9507 -13342 -9259 -13120
rect -9037 -13342 -8789 -13120
rect -8567 -13342 -8319 -13120
rect -8097 -13342 -7849 -13120
rect -7627 -13342 -7379 -13120
rect -7157 -13342 -6909 -13120
rect -6687 -13342 -6439 -13120
rect -6217 -13342 -5969 -13120
rect -5747 -13342 -5653 -13120
rect -13583 -13436 -5653 -13342
rect -13583 -13656 -12784 -13436
rect -12564 -13656 -12314 -13436
rect -12094 -13656 -11844 -13436
rect -11624 -13656 -11374 -13436
rect -11154 -13656 -10904 -13436
rect -10684 -13656 -10434 -13436
rect -10214 -13656 -9964 -13436
rect -9744 -13656 -9494 -13436
rect -9274 -13656 -9024 -13436
rect -8804 -13656 -8554 -13436
rect -8334 -13656 -8084 -13436
rect -7864 -13656 -7614 -13436
rect -7394 -13656 -7144 -13436
rect -6924 -13656 -6674 -13436
rect -6454 -13656 -5653 -13436
rect -13583 -13714 -5653 -13656
rect -5138 -13340 -4908 -13092
rect -5138 -13562 -5134 -13340
rect -4912 -13562 -4908 -13340
rect -5138 -13916 -4908 -13562
rect -14328 -14146 -4908 -13916
rect 396 -9756 25672 -1016
rect 28396 -1785 55820 -770
rect 56492 1489 58090 25794
rect 58502 25309 58578 25794
rect 58990 25309 59066 25794
rect 59478 25309 59554 25794
rect 59966 25309 60042 25794
rect 60454 25309 60530 25794
rect 60942 25309 61018 25794
rect 61430 25309 61506 25794
rect 61918 25309 61994 25794
rect 62406 25309 62482 25794
rect 62894 25309 62970 25794
rect 63382 25309 63458 25794
rect 63870 25309 63946 25794
rect 64358 25309 64434 25794
rect 64846 25309 64922 25794
rect 65334 25309 65410 25794
rect 65822 25309 65898 25794
rect 66310 25309 66386 25794
rect 66798 25309 66874 25794
rect 67286 25309 67362 25794
rect 67774 25309 67850 25794
rect 68262 25309 68338 25794
rect 68750 25309 68826 25794
rect 69238 25309 69314 25794
rect 69726 25309 69802 25794
rect 70214 25309 70290 25794
rect 70702 25309 70778 25794
rect 71190 25309 71266 25794
rect 71678 25309 71754 25794
rect 72166 25309 72242 25794
rect 72654 25309 72730 25794
rect 73142 25309 73218 25794
rect 73630 25309 73706 25794
rect 74118 25309 74194 25794
rect 74606 25309 74682 25794
rect 75094 25309 75170 25794
rect 75582 25309 75658 25794
rect 76070 25309 76146 25794
rect 76558 25309 76634 25794
rect 77046 25309 77122 25794
rect 77534 25309 77610 25794
rect 78022 25309 78098 25794
rect 78510 25309 78586 25794
rect 78998 25309 79074 25794
rect 79486 25309 79562 25794
rect 79974 25309 80050 25794
rect 80462 25309 80538 25794
rect 80950 25309 81026 25794
rect 81438 25309 81514 25794
rect 81926 25309 82002 25794
rect 82414 25309 82490 25794
rect 85014 25309 85090 25794
rect 85502 25309 85578 25794
rect 85990 25309 86066 25794
rect 86478 25309 86554 25794
rect 86966 25309 87042 25794
rect 87454 25309 87530 25794
rect 87942 25309 88018 25794
rect 88430 25309 88506 25794
rect 88918 25309 88994 25794
rect 89406 25309 89482 25794
rect 89894 25309 89970 25794
rect 90382 25309 90458 25794
rect 90870 25309 90946 25794
rect 91358 25309 91434 25794
rect 91846 25309 91922 25794
rect 92334 25309 92410 25794
rect 92822 25309 92898 25794
rect 93310 25309 93386 25794
rect 93798 25309 93874 25794
rect 94286 25309 94362 25794
rect 94774 25309 94850 25794
rect 95262 25309 95338 25794
rect 95750 25309 95826 25794
rect 96238 25309 96314 25794
rect 96726 25309 96802 25794
rect 97214 25309 97290 25794
rect 97702 25309 97778 25794
rect 98190 25309 98266 25794
rect 98678 25309 98754 25794
rect 99166 25309 99242 25794
rect 99654 25309 99730 25794
rect 100142 25309 100218 25794
rect 100630 25309 100706 25794
rect 101118 25309 101194 25794
rect 101606 25309 101682 25794
rect 102094 25309 102170 25794
rect 102582 25309 102658 25794
rect 103070 25309 103146 25794
rect 103558 25309 103634 25794
rect 104046 25309 104122 25794
rect 104534 25309 104610 25794
rect 105022 25309 105098 25794
rect 105510 25309 105586 25794
rect 105998 25309 106074 25794
rect 106486 25309 106562 25794
rect 106974 25309 107050 25794
rect 107462 25309 107538 25794
rect 107950 25309 108026 25794
rect 108438 25309 108514 25794
rect 108926 25309 109002 25794
rect 109414 25309 109490 25794
rect 84856 5305 85090 25307
rect 58258 4820 58334 5305
rect 58746 4820 58822 5305
rect 59234 4820 59310 5305
rect 59722 4820 59798 5305
rect 60210 4820 60286 5305
rect 60698 4820 60774 5305
rect 61186 4820 61262 5305
rect 61674 4820 61750 5305
rect 62162 4820 62238 5305
rect 62650 4820 62726 5305
rect 63138 4820 63214 5305
rect 63626 4820 63702 5305
rect 64114 4820 64190 5305
rect 64602 4820 64678 5305
rect 65090 4820 65166 5305
rect 65578 4820 65654 5305
rect 66066 4820 66142 5305
rect 66554 4820 66630 5305
rect 67042 4820 67118 5305
rect 67530 4820 67606 5305
rect 68018 4820 68094 5305
rect 68506 4820 68582 5305
rect 68994 4820 69070 5305
rect 69482 4820 69558 5305
rect 69970 4820 70046 5305
rect 70458 4820 70534 5305
rect 70946 4820 71022 5305
rect 71434 4820 71510 5305
rect 71922 4820 71998 5305
rect 72410 4820 72486 5305
rect 72898 4820 72974 5305
rect 73386 4820 73462 5305
rect 73874 4820 73950 5305
rect 74362 4820 74438 5305
rect 74850 4820 74926 5305
rect 75338 4820 75414 5305
rect 75826 4820 75902 5305
rect 76314 4820 76390 5305
rect 76802 4820 76878 5305
rect 77290 4820 77366 5305
rect 77778 4820 77854 5305
rect 78266 4820 78342 5305
rect 78754 4820 78830 5305
rect 79242 4820 79318 5305
rect 79730 4820 79806 5305
rect 80218 4820 80294 5305
rect 80706 4820 80782 5305
rect 81194 4820 81270 5305
rect 81682 4820 81758 5305
rect 82170 4820 82246 5305
rect 85258 4820 85334 5305
rect 85746 4820 85822 5305
rect 86234 4820 86310 5305
rect 86722 4820 86798 5305
rect 87210 4820 87286 5305
rect 87698 4820 87774 5305
rect 88186 4820 88262 5305
rect 88674 4820 88750 5305
rect 89162 4820 89238 5305
rect 89650 4820 89726 5305
rect 90138 4820 90214 5305
rect 90626 4820 90702 5305
rect 91114 4820 91190 5305
rect 91602 4820 91678 5305
rect 92090 4820 92166 5305
rect 92578 4820 92654 5305
rect 93066 4820 93142 5305
rect 93554 4820 93630 5305
rect 94042 4820 94118 5305
rect 94530 4820 94606 5305
rect 95018 4820 95094 5305
rect 95506 4820 95582 5305
rect 95994 4820 96070 5305
rect 96482 4820 96558 5305
rect 96970 4820 97046 5305
rect 97458 4820 97534 5305
rect 97946 4820 98022 5305
rect 98434 4820 98510 5305
rect 98922 4820 98998 5305
rect 99410 4820 99486 5305
rect 99898 4820 99974 5305
rect 100386 4820 100462 5305
rect 100874 4820 100950 5305
rect 101362 4820 101438 5305
rect 101850 4820 101926 5305
rect 102338 4820 102414 5305
rect 102826 4820 102902 5305
rect 103314 4820 103390 5305
rect 103802 4820 103878 5305
rect 104290 4820 104366 5305
rect 104778 4820 104854 5305
rect 105266 4820 105342 5305
rect 105754 4820 105830 5305
rect 106242 4820 106318 5305
rect 106730 4820 106806 5305
rect 107218 4820 107294 5305
rect 107706 4820 107782 5305
rect 108194 4820 108270 5305
rect 108682 4820 108758 5305
rect 109170 4820 109246 5305
rect 58258 4125 111646 4820
rect 56492 794 109490 1489
rect 396 -9800 9195 -9756
rect 9239 -9800 9295 -9756
rect 9339 -9800 9395 -9756
rect 9439 -9800 9495 -9756
rect 9539 -9800 9595 -9756
rect 9639 -9800 9695 -9756
rect 9739 -9800 9795 -9756
rect 9839 -9800 9895 -9756
rect 9939 -9800 9995 -9756
rect 10039 -9800 10095 -9756
rect 10139 -9800 10195 -9756
rect 10239 -9800 10295 -9756
rect 10339 -9800 10395 -9756
rect 10439 -9800 10495 -9756
rect 10539 -9800 10595 -9756
rect 10639 -9800 10695 -9756
rect 10739 -9800 11195 -9756
rect 11239 -9800 11295 -9756
rect 11339 -9800 11395 -9756
rect 11439 -9800 11495 -9756
rect 11539 -9800 11595 -9756
rect 11639 -9800 11695 -9756
rect 11739 -9800 11795 -9756
rect 11839 -9800 11895 -9756
rect 11939 -9800 11995 -9756
rect 12039 -9800 12095 -9756
rect 12139 -9800 12195 -9756
rect 12239 -9800 12295 -9756
rect 12339 -9800 12395 -9756
rect 12439 -9800 12495 -9756
rect 12539 -9800 12595 -9756
rect 12639 -9800 12695 -9756
rect 12739 -9800 13195 -9756
rect 13239 -9800 13295 -9756
rect 13339 -9800 13395 -9756
rect 13439 -9800 13495 -9756
rect 13539 -9800 13595 -9756
rect 13639 -9800 13695 -9756
rect 13739 -9800 13795 -9756
rect 13839 -9800 13895 -9756
rect 13939 -9800 13995 -9756
rect 14039 -9800 14095 -9756
rect 14139 -9800 14195 -9756
rect 14239 -9800 14295 -9756
rect 14339 -9800 14395 -9756
rect 14439 -9800 14495 -9756
rect 14539 -9800 14595 -9756
rect 14639 -9800 14695 -9756
rect 14739 -9800 15195 -9756
rect 15239 -9800 15295 -9756
rect 15339 -9800 15395 -9756
rect 15439 -9800 15495 -9756
rect 15539 -9800 15595 -9756
rect 15639 -9800 15695 -9756
rect 15739 -9800 15795 -9756
rect 15839 -9800 15895 -9756
rect 15939 -9800 15995 -9756
rect 16039 -9800 16095 -9756
rect 16139 -9800 16195 -9756
rect 16239 -9800 16295 -9756
rect 16339 -9800 16395 -9756
rect 16439 -9800 16495 -9756
rect 16539 -9800 16595 -9756
rect 16639 -9800 16695 -9756
rect 16739 -9800 25672 -9756
rect 396 -9856 25672 -9800
rect 396 -9900 9195 -9856
rect 9239 -9900 9295 -9856
rect 9339 -9900 9395 -9856
rect 9439 -9900 9495 -9856
rect 9539 -9900 9595 -9856
rect 9639 -9900 9695 -9856
rect 9739 -9900 9795 -9856
rect 9839 -9900 9895 -9856
rect 9939 -9900 9995 -9856
rect 10039 -9900 10095 -9856
rect 10139 -9900 10195 -9856
rect 10239 -9900 10295 -9856
rect 10339 -9900 10395 -9856
rect 10439 -9900 10495 -9856
rect 10539 -9900 10595 -9856
rect 10639 -9900 10695 -9856
rect 10739 -9900 11195 -9856
rect 11239 -9900 11295 -9856
rect 11339 -9900 11395 -9856
rect 11439 -9900 11495 -9856
rect 11539 -9900 11595 -9856
rect 11639 -9900 11695 -9856
rect 11739 -9900 11795 -9856
rect 11839 -9900 11895 -9856
rect 11939 -9900 11995 -9856
rect 12039 -9900 12095 -9856
rect 12139 -9900 12195 -9856
rect 12239 -9900 12295 -9856
rect 12339 -9900 12395 -9856
rect 12439 -9900 12495 -9856
rect 12539 -9900 12595 -9856
rect 12639 -9900 12695 -9856
rect 12739 -9900 13195 -9856
rect 13239 -9900 13295 -9856
rect 13339 -9900 13395 -9856
rect 13439 -9900 13495 -9856
rect 13539 -9900 13595 -9856
rect 13639 -9900 13695 -9856
rect 13739 -9900 13795 -9856
rect 13839 -9900 13895 -9856
rect 13939 -9900 13995 -9856
rect 14039 -9900 14095 -9856
rect 14139 -9900 14195 -9856
rect 14239 -9900 14295 -9856
rect 14339 -9900 14395 -9856
rect 14439 -9900 14495 -9856
rect 14539 -9900 14595 -9856
rect 14639 -9900 14695 -9856
rect 14739 -9900 15195 -9856
rect 15239 -9900 15295 -9856
rect 15339 -9900 15395 -9856
rect 15439 -9900 15495 -9856
rect 15539 -9900 15595 -9856
rect 15639 -9900 15695 -9856
rect 15739 -9900 15795 -9856
rect 15839 -9900 15895 -9856
rect 15939 -9900 15995 -9856
rect 16039 -9900 16095 -9856
rect 16139 -9900 16195 -9856
rect 16239 -9900 16295 -9856
rect 16339 -9900 16395 -9856
rect 16439 -9900 16495 -9856
rect 16539 -9900 16595 -9856
rect 16639 -9900 16695 -9856
rect 16739 -9900 25672 -9856
rect 396 -9956 25672 -9900
rect 396 -10000 9195 -9956
rect 9239 -10000 9295 -9956
rect 9339 -10000 9395 -9956
rect 9439 -10000 9495 -9956
rect 9539 -10000 9595 -9956
rect 9639 -10000 9695 -9956
rect 9739 -10000 9795 -9956
rect 9839 -10000 9895 -9956
rect 9939 -10000 9995 -9956
rect 10039 -10000 10095 -9956
rect 10139 -10000 10195 -9956
rect 10239 -10000 10295 -9956
rect 10339 -10000 10395 -9956
rect 10439 -10000 10495 -9956
rect 10539 -10000 10595 -9956
rect 10639 -10000 10695 -9956
rect 10739 -10000 11195 -9956
rect 11239 -10000 11295 -9956
rect 11339 -10000 11395 -9956
rect 11439 -10000 11495 -9956
rect 11539 -10000 11595 -9956
rect 11639 -10000 11695 -9956
rect 11739 -10000 11795 -9956
rect 11839 -10000 11895 -9956
rect 11939 -10000 11995 -9956
rect 12039 -10000 12095 -9956
rect 12139 -10000 12195 -9956
rect 12239 -10000 12295 -9956
rect 12339 -10000 12395 -9956
rect 12439 -10000 12495 -9956
rect 12539 -10000 12595 -9956
rect 12639 -10000 12695 -9956
rect 12739 -10000 13195 -9956
rect 13239 -10000 13295 -9956
rect 13339 -10000 13395 -9956
rect 13439 -10000 13495 -9956
rect 13539 -10000 13595 -9956
rect 13639 -10000 13695 -9956
rect 13739 -10000 13795 -9956
rect 13839 -10000 13895 -9956
rect 13939 -10000 13995 -9956
rect 14039 -10000 14095 -9956
rect 14139 -10000 14195 -9956
rect 14239 -10000 14295 -9956
rect 14339 -10000 14395 -9956
rect 14439 -10000 14495 -9956
rect 14539 -10000 14595 -9956
rect 14639 -10000 14695 -9956
rect 14739 -10000 15195 -9956
rect 15239 -10000 15295 -9956
rect 15339 -10000 15395 -9956
rect 15439 -10000 15495 -9956
rect 15539 -10000 15595 -9956
rect 15639 -10000 15695 -9956
rect 15739 -10000 15795 -9956
rect 15839 -10000 15895 -9956
rect 15939 -10000 15995 -9956
rect 16039 -10000 16095 -9956
rect 16139 -10000 16195 -9956
rect 16239 -10000 16295 -9956
rect 16339 -10000 16395 -9956
rect 16439 -10000 16495 -9956
rect 16539 -10000 16595 -9956
rect 16639 -10000 16695 -9956
rect 16739 -10000 25672 -9956
rect 396 -10056 25672 -10000
rect 396 -10100 9195 -10056
rect 9239 -10100 9295 -10056
rect 9339 -10100 9395 -10056
rect 9439 -10100 9495 -10056
rect 9539 -10100 9595 -10056
rect 9639 -10100 9695 -10056
rect 9739 -10100 9795 -10056
rect 9839 -10100 9895 -10056
rect 9939 -10100 9995 -10056
rect 10039 -10100 10095 -10056
rect 10139 -10100 10195 -10056
rect 10239 -10100 10295 -10056
rect 10339 -10100 10395 -10056
rect 10439 -10100 10495 -10056
rect 10539 -10100 10595 -10056
rect 10639 -10100 10695 -10056
rect 10739 -10100 11195 -10056
rect 11239 -10100 11295 -10056
rect 11339 -10100 11395 -10056
rect 11439 -10100 11495 -10056
rect 11539 -10100 11595 -10056
rect 11639 -10100 11695 -10056
rect 11739 -10100 11795 -10056
rect 11839 -10100 11895 -10056
rect 11939 -10100 11995 -10056
rect 12039 -10100 12095 -10056
rect 12139 -10100 12195 -10056
rect 12239 -10100 12295 -10056
rect 12339 -10100 12395 -10056
rect 12439 -10100 12495 -10056
rect 12539 -10100 12595 -10056
rect 12639 -10100 12695 -10056
rect 12739 -10100 13195 -10056
rect 13239 -10100 13295 -10056
rect 13339 -10100 13395 -10056
rect 13439 -10100 13495 -10056
rect 13539 -10100 13595 -10056
rect 13639 -10100 13695 -10056
rect 13739 -10100 13795 -10056
rect 13839 -10100 13895 -10056
rect 13939 -10100 13995 -10056
rect 14039 -10100 14095 -10056
rect 14139 -10100 14195 -10056
rect 14239 -10100 14295 -10056
rect 14339 -10100 14395 -10056
rect 14439 -10100 14495 -10056
rect 14539 -10100 14595 -10056
rect 14639 -10100 14695 -10056
rect 14739 -10100 15195 -10056
rect 15239 -10100 15295 -10056
rect 15339 -10100 15395 -10056
rect 15439 -10100 15495 -10056
rect 15539 -10100 15595 -10056
rect 15639 -10100 15695 -10056
rect 15739 -10100 15795 -10056
rect 15839 -10100 15895 -10056
rect 15939 -10100 15995 -10056
rect 16039 -10100 16095 -10056
rect 16139 -10100 16195 -10056
rect 16239 -10100 16295 -10056
rect 16339 -10100 16395 -10056
rect 16439 -10100 16495 -10056
rect 16539 -10100 16595 -10056
rect 16639 -10100 16695 -10056
rect 16739 -10100 25672 -10056
rect 396 -10156 25672 -10100
rect 396 -10200 9195 -10156
rect 9239 -10200 9295 -10156
rect 9339 -10200 9395 -10156
rect 9439 -10200 9495 -10156
rect 9539 -10200 9595 -10156
rect 9639 -10200 9695 -10156
rect 9739 -10200 9795 -10156
rect 9839 -10200 9895 -10156
rect 9939 -10200 9995 -10156
rect 10039 -10200 10095 -10156
rect 10139 -10200 10195 -10156
rect 10239 -10200 10295 -10156
rect 10339 -10200 10395 -10156
rect 10439 -10200 10495 -10156
rect 10539 -10200 10595 -10156
rect 10639 -10200 10695 -10156
rect 10739 -10200 11195 -10156
rect 11239 -10200 11295 -10156
rect 11339 -10200 11395 -10156
rect 11439 -10200 11495 -10156
rect 11539 -10200 11595 -10156
rect 11639 -10200 11695 -10156
rect 11739 -10200 11795 -10156
rect 11839 -10200 11895 -10156
rect 11939 -10200 11995 -10156
rect 12039 -10200 12095 -10156
rect 12139 -10200 12195 -10156
rect 12239 -10200 12295 -10156
rect 12339 -10200 12395 -10156
rect 12439 -10200 12495 -10156
rect 12539 -10200 12595 -10156
rect 12639 -10200 12695 -10156
rect 12739 -10200 13195 -10156
rect 13239 -10200 13295 -10156
rect 13339 -10200 13395 -10156
rect 13439 -10200 13495 -10156
rect 13539 -10200 13595 -10156
rect 13639 -10200 13695 -10156
rect 13739 -10200 13795 -10156
rect 13839 -10200 13895 -10156
rect 13939 -10200 13995 -10156
rect 14039 -10200 14095 -10156
rect 14139 -10200 14195 -10156
rect 14239 -10200 14295 -10156
rect 14339 -10200 14395 -10156
rect 14439 -10200 14495 -10156
rect 14539 -10200 14595 -10156
rect 14639 -10200 14695 -10156
rect 14739 -10200 15195 -10156
rect 15239 -10200 15295 -10156
rect 15339 -10200 15395 -10156
rect 15439 -10200 15495 -10156
rect 15539 -10200 15595 -10156
rect 15639 -10200 15695 -10156
rect 15739 -10200 15795 -10156
rect 15839 -10200 15895 -10156
rect 15939 -10200 15995 -10156
rect 16039 -10200 16095 -10156
rect 16139 -10200 16195 -10156
rect 16239 -10200 16295 -10156
rect 16339 -10200 16395 -10156
rect 16439 -10200 16495 -10156
rect 16539 -10200 16595 -10156
rect 16639 -10200 16695 -10156
rect 16739 -10200 25672 -10156
rect 396 -10256 25672 -10200
rect 396 -10300 9195 -10256
rect 9239 -10300 9295 -10256
rect 9339 -10300 9395 -10256
rect 9439 -10300 9495 -10256
rect 9539 -10300 9595 -10256
rect 9639 -10300 9695 -10256
rect 9739 -10300 9795 -10256
rect 9839 -10300 9895 -10256
rect 9939 -10300 9995 -10256
rect 10039 -10300 10095 -10256
rect 10139 -10300 10195 -10256
rect 10239 -10300 10295 -10256
rect 10339 -10300 10395 -10256
rect 10439 -10300 10495 -10256
rect 10539 -10300 10595 -10256
rect 10639 -10300 10695 -10256
rect 10739 -10300 11195 -10256
rect 11239 -10300 11295 -10256
rect 11339 -10300 11395 -10256
rect 11439 -10300 11495 -10256
rect 11539 -10300 11595 -10256
rect 11639 -10300 11695 -10256
rect 11739 -10300 11795 -10256
rect 11839 -10300 11895 -10256
rect 11939 -10300 11995 -10256
rect 12039 -10300 12095 -10256
rect 12139 -10300 12195 -10256
rect 12239 -10300 12295 -10256
rect 12339 -10300 12395 -10256
rect 12439 -10300 12495 -10256
rect 12539 -10300 12595 -10256
rect 12639 -10300 12695 -10256
rect 12739 -10300 13195 -10256
rect 13239 -10300 13295 -10256
rect 13339 -10300 13395 -10256
rect 13439 -10300 13495 -10256
rect 13539 -10300 13595 -10256
rect 13639 -10300 13695 -10256
rect 13739 -10300 13795 -10256
rect 13839 -10300 13895 -10256
rect 13939 -10300 13995 -10256
rect 14039 -10300 14095 -10256
rect 14139 -10300 14195 -10256
rect 14239 -10300 14295 -10256
rect 14339 -10300 14395 -10256
rect 14439 -10300 14495 -10256
rect 14539 -10300 14595 -10256
rect 14639 -10300 14695 -10256
rect 14739 -10300 15195 -10256
rect 15239 -10300 15295 -10256
rect 15339 -10300 15395 -10256
rect 15439 -10300 15495 -10256
rect 15539 -10300 15595 -10256
rect 15639 -10300 15695 -10256
rect 15739 -10300 15795 -10256
rect 15839 -10300 15895 -10256
rect 15939 -10300 15995 -10256
rect 16039 -10300 16095 -10256
rect 16139 -10300 16195 -10256
rect 16239 -10300 16295 -10256
rect 16339 -10300 16395 -10256
rect 16439 -10300 16495 -10256
rect 16539 -10300 16595 -10256
rect 16639 -10300 16695 -10256
rect 16739 -10300 25672 -10256
rect 396 -10356 25672 -10300
rect 396 -10400 9195 -10356
rect 9239 -10400 9295 -10356
rect 9339 -10400 9395 -10356
rect 9439 -10400 9495 -10356
rect 9539 -10400 9595 -10356
rect 9639 -10400 9695 -10356
rect 9739 -10400 9795 -10356
rect 9839 -10400 9895 -10356
rect 9939 -10400 9995 -10356
rect 10039 -10400 10095 -10356
rect 10139 -10400 10195 -10356
rect 10239 -10400 10295 -10356
rect 10339 -10400 10395 -10356
rect 10439 -10400 10495 -10356
rect 10539 -10400 10595 -10356
rect 10639 -10400 10695 -10356
rect 10739 -10400 11195 -10356
rect 11239 -10400 11295 -10356
rect 11339 -10400 11395 -10356
rect 11439 -10400 11495 -10356
rect 11539 -10400 11595 -10356
rect 11639 -10400 11695 -10356
rect 11739 -10400 11795 -10356
rect 11839 -10400 11895 -10356
rect 11939 -10400 11995 -10356
rect 12039 -10400 12095 -10356
rect 12139 -10400 12195 -10356
rect 12239 -10400 12295 -10356
rect 12339 -10400 12395 -10356
rect 12439 -10400 12495 -10356
rect 12539 -10400 12595 -10356
rect 12639 -10400 12695 -10356
rect 12739 -10400 13195 -10356
rect 13239 -10400 13295 -10356
rect 13339 -10400 13395 -10356
rect 13439 -10400 13495 -10356
rect 13539 -10400 13595 -10356
rect 13639 -10400 13695 -10356
rect 13739 -10400 13795 -10356
rect 13839 -10400 13895 -10356
rect 13939 -10400 13995 -10356
rect 14039 -10400 14095 -10356
rect 14139 -10400 14195 -10356
rect 14239 -10400 14295 -10356
rect 14339 -10400 14395 -10356
rect 14439 -10400 14495 -10356
rect 14539 -10400 14595 -10356
rect 14639 -10400 14695 -10356
rect 14739 -10400 15195 -10356
rect 15239 -10400 15295 -10356
rect 15339 -10400 15395 -10356
rect 15439 -10400 15495 -10356
rect 15539 -10400 15595 -10356
rect 15639 -10400 15695 -10356
rect 15739 -10400 15795 -10356
rect 15839 -10400 15895 -10356
rect 15939 -10400 15995 -10356
rect 16039 -10400 16095 -10356
rect 16139 -10400 16195 -10356
rect 16239 -10400 16295 -10356
rect 16339 -10400 16395 -10356
rect 16439 -10400 16495 -10356
rect 16539 -10400 16595 -10356
rect 16639 -10400 16695 -10356
rect 16739 -10400 25672 -10356
rect 396 -10456 25672 -10400
rect 396 -10500 9195 -10456
rect 9239 -10500 9295 -10456
rect 9339 -10500 9395 -10456
rect 9439 -10500 9495 -10456
rect 9539 -10500 9595 -10456
rect 9639 -10500 9695 -10456
rect 9739 -10500 9795 -10456
rect 9839 -10500 9895 -10456
rect 9939 -10500 9995 -10456
rect 10039 -10500 10095 -10456
rect 10139 -10500 10195 -10456
rect 10239 -10500 10295 -10456
rect 10339 -10500 10395 -10456
rect 10439 -10500 10495 -10456
rect 10539 -10500 10595 -10456
rect 10639 -10500 10695 -10456
rect 10739 -10500 11195 -10456
rect 11239 -10500 11295 -10456
rect 11339 -10500 11395 -10456
rect 11439 -10500 11495 -10456
rect 11539 -10500 11595 -10456
rect 11639 -10500 11695 -10456
rect 11739 -10500 11795 -10456
rect 11839 -10500 11895 -10456
rect 11939 -10500 11995 -10456
rect 12039 -10500 12095 -10456
rect 12139 -10500 12195 -10456
rect 12239 -10500 12295 -10456
rect 12339 -10500 12395 -10456
rect 12439 -10500 12495 -10456
rect 12539 -10500 12595 -10456
rect 12639 -10500 12695 -10456
rect 12739 -10500 13195 -10456
rect 13239 -10500 13295 -10456
rect 13339 -10500 13395 -10456
rect 13439 -10500 13495 -10456
rect 13539 -10500 13595 -10456
rect 13639 -10500 13695 -10456
rect 13739 -10500 13795 -10456
rect 13839 -10500 13895 -10456
rect 13939 -10500 13995 -10456
rect 14039 -10500 14095 -10456
rect 14139 -10500 14195 -10456
rect 14239 -10500 14295 -10456
rect 14339 -10500 14395 -10456
rect 14439 -10500 14495 -10456
rect 14539 -10500 14595 -10456
rect 14639 -10500 14695 -10456
rect 14739 -10500 15195 -10456
rect 15239 -10500 15295 -10456
rect 15339 -10500 15395 -10456
rect 15439 -10500 15495 -10456
rect 15539 -10500 15595 -10456
rect 15639 -10500 15695 -10456
rect 15739 -10500 15795 -10456
rect 15839 -10500 15895 -10456
rect 15939 -10500 15995 -10456
rect 16039 -10500 16095 -10456
rect 16139 -10500 16195 -10456
rect 16239 -10500 16295 -10456
rect 16339 -10500 16395 -10456
rect 16439 -10500 16495 -10456
rect 16539 -10500 16595 -10456
rect 16639 -10500 16695 -10456
rect 16739 -10500 25672 -10456
rect 396 -10556 25672 -10500
rect 396 -10600 9195 -10556
rect 9239 -10600 9295 -10556
rect 9339 -10600 9395 -10556
rect 9439 -10600 9495 -10556
rect 9539 -10600 9595 -10556
rect 9639 -10600 9695 -10556
rect 9739 -10600 9795 -10556
rect 9839 -10600 9895 -10556
rect 9939 -10600 9995 -10556
rect 10039 -10600 10095 -10556
rect 10139 -10600 10195 -10556
rect 10239 -10600 10295 -10556
rect 10339 -10600 10395 -10556
rect 10439 -10600 10495 -10556
rect 10539 -10600 10595 -10556
rect 10639 -10600 10695 -10556
rect 10739 -10600 11195 -10556
rect 11239 -10600 11295 -10556
rect 11339 -10600 11395 -10556
rect 11439 -10600 11495 -10556
rect 11539 -10600 11595 -10556
rect 11639 -10600 11695 -10556
rect 11739 -10600 11795 -10556
rect 11839 -10600 11895 -10556
rect 11939 -10600 11995 -10556
rect 12039 -10600 12095 -10556
rect 12139 -10600 12195 -10556
rect 12239 -10600 12295 -10556
rect 12339 -10600 12395 -10556
rect 12439 -10600 12495 -10556
rect 12539 -10600 12595 -10556
rect 12639 -10600 12695 -10556
rect 12739 -10600 13195 -10556
rect 13239 -10600 13295 -10556
rect 13339 -10600 13395 -10556
rect 13439 -10600 13495 -10556
rect 13539 -10600 13595 -10556
rect 13639 -10600 13695 -10556
rect 13739 -10600 13795 -10556
rect 13839 -10600 13895 -10556
rect 13939 -10600 13995 -10556
rect 14039 -10600 14095 -10556
rect 14139 -10600 14195 -10556
rect 14239 -10600 14295 -10556
rect 14339 -10600 14395 -10556
rect 14439 -10600 14495 -10556
rect 14539 -10600 14595 -10556
rect 14639 -10600 14695 -10556
rect 14739 -10600 15195 -10556
rect 15239 -10600 15295 -10556
rect 15339 -10600 15395 -10556
rect 15439 -10600 15495 -10556
rect 15539 -10600 15595 -10556
rect 15639 -10600 15695 -10556
rect 15739 -10600 15795 -10556
rect 15839 -10600 15895 -10556
rect 15939 -10600 15995 -10556
rect 16039 -10600 16095 -10556
rect 16139 -10600 16195 -10556
rect 16239 -10600 16295 -10556
rect 16339 -10600 16395 -10556
rect 16439 -10600 16495 -10556
rect 16539 -10600 16595 -10556
rect 16639 -10600 16695 -10556
rect 16739 -10600 25672 -10556
rect 396 -10656 25672 -10600
rect 396 -10700 9195 -10656
rect 9239 -10700 9295 -10656
rect 9339 -10700 9395 -10656
rect 9439 -10700 9495 -10656
rect 9539 -10700 9595 -10656
rect 9639 -10700 9695 -10656
rect 9739 -10700 9795 -10656
rect 9839 -10700 9895 -10656
rect 9939 -10700 9995 -10656
rect 10039 -10700 10095 -10656
rect 10139 -10700 10195 -10656
rect 10239 -10700 10295 -10656
rect 10339 -10700 10395 -10656
rect 10439 -10700 10495 -10656
rect 10539 -10700 10595 -10656
rect 10639 -10700 10695 -10656
rect 10739 -10700 11195 -10656
rect 11239 -10700 11295 -10656
rect 11339 -10700 11395 -10656
rect 11439 -10700 11495 -10656
rect 11539 -10700 11595 -10656
rect 11639 -10700 11695 -10656
rect 11739 -10700 11795 -10656
rect 11839 -10700 11895 -10656
rect 11939 -10700 11995 -10656
rect 12039 -10700 12095 -10656
rect 12139 -10700 12195 -10656
rect 12239 -10700 12295 -10656
rect 12339 -10700 12395 -10656
rect 12439 -10700 12495 -10656
rect 12539 -10700 12595 -10656
rect 12639 -10700 12695 -10656
rect 12739 -10700 13195 -10656
rect 13239 -10700 13295 -10656
rect 13339 -10700 13395 -10656
rect 13439 -10700 13495 -10656
rect 13539 -10700 13595 -10656
rect 13639 -10700 13695 -10656
rect 13739 -10700 13795 -10656
rect 13839 -10700 13895 -10656
rect 13939 -10700 13995 -10656
rect 14039 -10700 14095 -10656
rect 14139 -10700 14195 -10656
rect 14239 -10700 14295 -10656
rect 14339 -10700 14395 -10656
rect 14439 -10700 14495 -10656
rect 14539 -10700 14595 -10656
rect 14639 -10700 14695 -10656
rect 14739 -10700 15195 -10656
rect 15239 -10700 15295 -10656
rect 15339 -10700 15395 -10656
rect 15439 -10700 15495 -10656
rect 15539 -10700 15595 -10656
rect 15639 -10700 15695 -10656
rect 15739 -10700 15795 -10656
rect 15839 -10700 15895 -10656
rect 15939 -10700 15995 -10656
rect 16039 -10700 16095 -10656
rect 16139 -10700 16195 -10656
rect 16239 -10700 16295 -10656
rect 16339 -10700 16395 -10656
rect 16439 -10700 16495 -10656
rect 16539 -10700 16595 -10656
rect 16639 -10700 16695 -10656
rect 16739 -10700 25672 -10656
rect 396 -10756 25672 -10700
rect 396 -10800 9195 -10756
rect 9239 -10800 9295 -10756
rect 9339 -10800 9395 -10756
rect 9439 -10800 9495 -10756
rect 9539 -10800 9595 -10756
rect 9639 -10800 9695 -10756
rect 9739 -10800 9795 -10756
rect 9839 -10800 9895 -10756
rect 9939 -10800 9995 -10756
rect 10039 -10800 10095 -10756
rect 10139 -10800 10195 -10756
rect 10239 -10800 10295 -10756
rect 10339 -10800 10395 -10756
rect 10439 -10800 10495 -10756
rect 10539 -10800 10595 -10756
rect 10639 -10800 10695 -10756
rect 10739 -10800 11195 -10756
rect 11239 -10800 11295 -10756
rect 11339 -10800 11395 -10756
rect 11439 -10800 11495 -10756
rect 11539 -10800 11595 -10756
rect 11639 -10800 11695 -10756
rect 11739 -10800 11795 -10756
rect 11839 -10800 11895 -10756
rect 11939 -10800 11995 -10756
rect 12039 -10800 12095 -10756
rect 12139 -10800 12195 -10756
rect 12239 -10800 12295 -10756
rect 12339 -10800 12395 -10756
rect 12439 -10800 12495 -10756
rect 12539 -10800 12595 -10756
rect 12639 -10800 12695 -10756
rect 12739 -10800 13195 -10756
rect 13239 -10800 13295 -10756
rect 13339 -10800 13395 -10756
rect 13439 -10800 13495 -10756
rect 13539 -10800 13595 -10756
rect 13639 -10800 13695 -10756
rect 13739 -10800 13795 -10756
rect 13839 -10800 13895 -10756
rect 13939 -10800 13995 -10756
rect 14039 -10800 14095 -10756
rect 14139 -10800 14195 -10756
rect 14239 -10800 14295 -10756
rect 14339 -10800 14395 -10756
rect 14439 -10800 14495 -10756
rect 14539 -10800 14595 -10756
rect 14639 -10800 14695 -10756
rect 14739 -10800 15195 -10756
rect 15239 -10800 15295 -10756
rect 15339 -10800 15395 -10756
rect 15439 -10800 15495 -10756
rect 15539 -10800 15595 -10756
rect 15639 -10800 15695 -10756
rect 15739 -10800 15795 -10756
rect 15839 -10800 15895 -10756
rect 15939 -10800 15995 -10756
rect 16039 -10800 16095 -10756
rect 16139 -10800 16195 -10756
rect 16239 -10800 16295 -10756
rect 16339 -10800 16395 -10756
rect 16439 -10800 16495 -10756
rect 16539 -10800 16595 -10756
rect 16639 -10800 16695 -10756
rect 16739 -10800 25672 -10756
rect 396 -10856 25672 -10800
rect 396 -10900 9195 -10856
rect 9239 -10900 9295 -10856
rect 9339 -10900 9395 -10856
rect 9439 -10900 9495 -10856
rect 9539 -10900 9595 -10856
rect 9639 -10900 9695 -10856
rect 9739 -10900 9795 -10856
rect 9839 -10900 9895 -10856
rect 9939 -10900 9995 -10856
rect 10039 -10900 10095 -10856
rect 10139 -10900 10195 -10856
rect 10239 -10900 10295 -10856
rect 10339 -10900 10395 -10856
rect 10439 -10900 10495 -10856
rect 10539 -10900 10595 -10856
rect 10639 -10900 10695 -10856
rect 10739 -10900 11195 -10856
rect 11239 -10900 11295 -10856
rect 11339 -10900 11395 -10856
rect 11439 -10900 11495 -10856
rect 11539 -10900 11595 -10856
rect 11639 -10900 11695 -10856
rect 11739 -10900 11795 -10856
rect 11839 -10900 11895 -10856
rect 11939 -10900 11995 -10856
rect 12039 -10900 12095 -10856
rect 12139 -10900 12195 -10856
rect 12239 -10900 12295 -10856
rect 12339 -10900 12395 -10856
rect 12439 -10900 12495 -10856
rect 12539 -10900 12595 -10856
rect 12639 -10900 12695 -10856
rect 12739 -10900 13195 -10856
rect 13239 -10900 13295 -10856
rect 13339 -10900 13395 -10856
rect 13439 -10900 13495 -10856
rect 13539 -10900 13595 -10856
rect 13639 -10900 13695 -10856
rect 13739 -10900 13795 -10856
rect 13839 -10900 13895 -10856
rect 13939 -10900 13995 -10856
rect 14039 -10900 14095 -10856
rect 14139 -10900 14195 -10856
rect 14239 -10900 14295 -10856
rect 14339 -10900 14395 -10856
rect 14439 -10900 14495 -10856
rect 14539 -10900 14595 -10856
rect 14639 -10900 14695 -10856
rect 14739 -10900 15195 -10856
rect 15239 -10900 15295 -10856
rect 15339 -10900 15395 -10856
rect 15439 -10900 15495 -10856
rect 15539 -10900 15595 -10856
rect 15639 -10900 15695 -10856
rect 15739 -10900 15795 -10856
rect 15839 -10900 15895 -10856
rect 15939 -10900 15995 -10856
rect 16039 -10900 16095 -10856
rect 16139 -10900 16195 -10856
rect 16239 -10900 16295 -10856
rect 16339 -10900 16395 -10856
rect 16439 -10900 16495 -10856
rect 16539 -10900 16595 -10856
rect 16639 -10900 16695 -10856
rect 16739 -10900 25672 -10856
rect 396 -10956 25672 -10900
rect 396 -11000 9195 -10956
rect 9239 -11000 9295 -10956
rect 9339 -11000 9395 -10956
rect 9439 -11000 9495 -10956
rect 9539 -11000 9595 -10956
rect 9639 -11000 9695 -10956
rect 9739 -11000 9795 -10956
rect 9839 -11000 9895 -10956
rect 9939 -11000 9995 -10956
rect 10039 -11000 10095 -10956
rect 10139 -11000 10195 -10956
rect 10239 -11000 10295 -10956
rect 10339 -11000 10395 -10956
rect 10439 -11000 10495 -10956
rect 10539 -11000 10595 -10956
rect 10639 -11000 10695 -10956
rect 10739 -11000 11195 -10956
rect 11239 -11000 11295 -10956
rect 11339 -11000 11395 -10956
rect 11439 -11000 11495 -10956
rect 11539 -11000 11595 -10956
rect 11639 -11000 11695 -10956
rect 11739 -11000 11795 -10956
rect 11839 -11000 11895 -10956
rect 11939 -11000 11995 -10956
rect 12039 -11000 12095 -10956
rect 12139 -11000 12195 -10956
rect 12239 -11000 12295 -10956
rect 12339 -11000 12395 -10956
rect 12439 -11000 12495 -10956
rect 12539 -11000 12595 -10956
rect 12639 -11000 12695 -10956
rect 12739 -11000 13195 -10956
rect 13239 -11000 13295 -10956
rect 13339 -11000 13395 -10956
rect 13439 -11000 13495 -10956
rect 13539 -11000 13595 -10956
rect 13639 -11000 13695 -10956
rect 13739 -11000 13795 -10956
rect 13839 -11000 13895 -10956
rect 13939 -11000 13995 -10956
rect 14039 -11000 14095 -10956
rect 14139 -11000 14195 -10956
rect 14239 -11000 14295 -10956
rect 14339 -11000 14395 -10956
rect 14439 -11000 14495 -10956
rect 14539 -11000 14595 -10956
rect 14639 -11000 14695 -10956
rect 14739 -11000 15195 -10956
rect 15239 -11000 15295 -10956
rect 15339 -11000 15395 -10956
rect 15439 -11000 15495 -10956
rect 15539 -11000 15595 -10956
rect 15639 -11000 15695 -10956
rect 15739 -11000 15795 -10956
rect 15839 -11000 15895 -10956
rect 15939 -11000 15995 -10956
rect 16039 -11000 16095 -10956
rect 16139 -11000 16195 -10956
rect 16239 -11000 16295 -10956
rect 16339 -11000 16395 -10956
rect 16439 -11000 16495 -10956
rect 16539 -11000 16595 -10956
rect 16639 -11000 16695 -10956
rect 16739 -11000 25672 -10956
rect 396 -11056 25672 -11000
rect 396 -11100 9195 -11056
rect 9239 -11100 9295 -11056
rect 9339 -11100 9395 -11056
rect 9439 -11100 9495 -11056
rect 9539 -11100 9595 -11056
rect 9639 -11100 9695 -11056
rect 9739 -11100 9795 -11056
rect 9839 -11100 9895 -11056
rect 9939 -11100 9995 -11056
rect 10039 -11100 10095 -11056
rect 10139 -11100 10195 -11056
rect 10239 -11100 10295 -11056
rect 10339 -11100 10395 -11056
rect 10439 -11100 10495 -11056
rect 10539 -11100 10595 -11056
rect 10639 -11100 10695 -11056
rect 10739 -11100 11195 -11056
rect 11239 -11100 11295 -11056
rect 11339 -11100 11395 -11056
rect 11439 -11100 11495 -11056
rect 11539 -11100 11595 -11056
rect 11639 -11100 11695 -11056
rect 11739 -11100 11795 -11056
rect 11839 -11100 11895 -11056
rect 11939 -11100 11995 -11056
rect 12039 -11100 12095 -11056
rect 12139 -11100 12195 -11056
rect 12239 -11100 12295 -11056
rect 12339 -11100 12395 -11056
rect 12439 -11100 12495 -11056
rect 12539 -11100 12595 -11056
rect 12639 -11100 12695 -11056
rect 12739 -11100 13195 -11056
rect 13239 -11100 13295 -11056
rect 13339 -11100 13395 -11056
rect 13439 -11100 13495 -11056
rect 13539 -11100 13595 -11056
rect 13639 -11100 13695 -11056
rect 13739 -11100 13795 -11056
rect 13839 -11100 13895 -11056
rect 13939 -11100 13995 -11056
rect 14039 -11100 14095 -11056
rect 14139 -11100 14195 -11056
rect 14239 -11100 14295 -11056
rect 14339 -11100 14395 -11056
rect 14439 -11100 14495 -11056
rect 14539 -11100 14595 -11056
rect 14639 -11100 14695 -11056
rect 14739 -11100 15195 -11056
rect 15239 -11100 15295 -11056
rect 15339 -11100 15395 -11056
rect 15439 -11100 15495 -11056
rect 15539 -11100 15595 -11056
rect 15639 -11100 15695 -11056
rect 15739 -11100 15795 -11056
rect 15839 -11100 15895 -11056
rect 15939 -11100 15995 -11056
rect 16039 -11100 16095 -11056
rect 16139 -11100 16195 -11056
rect 16239 -11100 16295 -11056
rect 16339 -11100 16395 -11056
rect 16439 -11100 16495 -11056
rect 16539 -11100 16595 -11056
rect 16639 -11100 16695 -11056
rect 16739 -11100 25672 -11056
rect 396 -11156 25672 -11100
rect 396 -11200 9195 -11156
rect 9239 -11200 9295 -11156
rect 9339 -11200 9395 -11156
rect 9439 -11200 9495 -11156
rect 9539 -11200 9595 -11156
rect 9639 -11200 9695 -11156
rect 9739 -11200 9795 -11156
rect 9839 -11200 9895 -11156
rect 9939 -11200 9995 -11156
rect 10039 -11200 10095 -11156
rect 10139 -11200 10195 -11156
rect 10239 -11200 10295 -11156
rect 10339 -11200 10395 -11156
rect 10439 -11200 10495 -11156
rect 10539 -11200 10595 -11156
rect 10639 -11200 10695 -11156
rect 10739 -11200 11195 -11156
rect 11239 -11200 11295 -11156
rect 11339 -11200 11395 -11156
rect 11439 -11200 11495 -11156
rect 11539 -11200 11595 -11156
rect 11639 -11200 11695 -11156
rect 11739 -11200 11795 -11156
rect 11839 -11200 11895 -11156
rect 11939 -11200 11995 -11156
rect 12039 -11200 12095 -11156
rect 12139 -11200 12195 -11156
rect 12239 -11200 12295 -11156
rect 12339 -11200 12395 -11156
rect 12439 -11200 12495 -11156
rect 12539 -11200 12595 -11156
rect 12639 -11200 12695 -11156
rect 12739 -11200 13195 -11156
rect 13239 -11200 13295 -11156
rect 13339 -11200 13395 -11156
rect 13439 -11200 13495 -11156
rect 13539 -11200 13595 -11156
rect 13639 -11200 13695 -11156
rect 13739 -11200 13795 -11156
rect 13839 -11200 13895 -11156
rect 13939 -11200 13995 -11156
rect 14039 -11200 14095 -11156
rect 14139 -11200 14195 -11156
rect 14239 -11200 14295 -11156
rect 14339 -11200 14395 -11156
rect 14439 -11200 14495 -11156
rect 14539 -11200 14595 -11156
rect 14639 -11200 14695 -11156
rect 14739 -11200 15195 -11156
rect 15239 -11200 15295 -11156
rect 15339 -11200 15395 -11156
rect 15439 -11200 15495 -11156
rect 15539 -11200 15595 -11156
rect 15639 -11200 15695 -11156
rect 15739 -11200 15795 -11156
rect 15839 -11200 15895 -11156
rect 15939 -11200 15995 -11156
rect 16039 -11200 16095 -11156
rect 16139 -11200 16195 -11156
rect 16239 -11200 16295 -11156
rect 16339 -11200 16395 -11156
rect 16439 -11200 16495 -11156
rect 16539 -11200 16595 -11156
rect 16639 -11200 16695 -11156
rect 16739 -11200 25672 -11156
rect 396 -11256 25672 -11200
rect 396 -11300 9195 -11256
rect 9239 -11300 9295 -11256
rect 9339 -11300 9395 -11256
rect 9439 -11300 9495 -11256
rect 9539 -11300 9595 -11256
rect 9639 -11300 9695 -11256
rect 9739 -11300 9795 -11256
rect 9839 -11300 9895 -11256
rect 9939 -11300 9995 -11256
rect 10039 -11300 10095 -11256
rect 10139 -11300 10195 -11256
rect 10239 -11300 10295 -11256
rect 10339 -11300 10395 -11256
rect 10439 -11300 10495 -11256
rect 10539 -11300 10595 -11256
rect 10639 -11300 10695 -11256
rect 10739 -11300 11195 -11256
rect 11239 -11300 11295 -11256
rect 11339 -11300 11395 -11256
rect 11439 -11300 11495 -11256
rect 11539 -11300 11595 -11256
rect 11639 -11300 11695 -11256
rect 11739 -11300 11795 -11256
rect 11839 -11300 11895 -11256
rect 11939 -11300 11995 -11256
rect 12039 -11300 12095 -11256
rect 12139 -11300 12195 -11256
rect 12239 -11300 12295 -11256
rect 12339 -11300 12395 -11256
rect 12439 -11300 12495 -11256
rect 12539 -11300 12595 -11256
rect 12639 -11300 12695 -11256
rect 12739 -11300 13195 -11256
rect 13239 -11300 13295 -11256
rect 13339 -11300 13395 -11256
rect 13439 -11300 13495 -11256
rect 13539 -11300 13595 -11256
rect 13639 -11300 13695 -11256
rect 13739 -11300 13795 -11256
rect 13839 -11300 13895 -11256
rect 13939 -11300 13995 -11256
rect 14039 -11300 14095 -11256
rect 14139 -11300 14195 -11256
rect 14239 -11300 14295 -11256
rect 14339 -11300 14395 -11256
rect 14439 -11300 14495 -11256
rect 14539 -11300 14595 -11256
rect 14639 -11300 14695 -11256
rect 14739 -11300 15195 -11256
rect 15239 -11300 15295 -11256
rect 15339 -11300 15395 -11256
rect 15439 -11300 15495 -11256
rect 15539 -11300 15595 -11256
rect 15639 -11300 15695 -11256
rect 15739 -11300 15795 -11256
rect 15839 -11300 15895 -11256
rect 15939 -11300 15995 -11256
rect 16039 -11300 16095 -11256
rect 16139 -11300 16195 -11256
rect 16239 -11300 16295 -11256
rect 16339 -11300 16395 -11256
rect 16439 -11300 16495 -11256
rect 16539 -11300 16595 -11256
rect 16639 -11300 16695 -11256
rect 16739 -11300 25672 -11256
rect 396 -19035 25672 -11300
rect 34207 -9638 50994 -1785
rect 34207 -9682 37223 -9638
rect 37267 -9682 37323 -9638
rect 37367 -9682 37423 -9638
rect 37467 -9682 37523 -9638
rect 37567 -9682 37623 -9638
rect 37667 -9682 37723 -9638
rect 37767 -9682 37823 -9638
rect 37867 -9682 37923 -9638
rect 37967 -9682 38023 -9638
rect 38067 -9682 38123 -9638
rect 38167 -9682 38223 -9638
rect 38267 -9682 38323 -9638
rect 38367 -9682 38423 -9638
rect 38467 -9682 38523 -9638
rect 38567 -9682 38623 -9638
rect 38667 -9682 38723 -9638
rect 38767 -9682 39223 -9638
rect 39267 -9682 39323 -9638
rect 39367 -9682 39423 -9638
rect 39467 -9682 39523 -9638
rect 39567 -9682 39623 -9638
rect 39667 -9682 39723 -9638
rect 39767 -9682 39823 -9638
rect 39867 -9682 39923 -9638
rect 39967 -9682 40023 -9638
rect 40067 -9682 40123 -9638
rect 40167 -9682 40223 -9638
rect 40267 -9682 40323 -9638
rect 40367 -9682 40423 -9638
rect 40467 -9682 40523 -9638
rect 40567 -9682 40623 -9638
rect 40667 -9682 40723 -9638
rect 40767 -9682 41223 -9638
rect 41267 -9682 41323 -9638
rect 41367 -9682 41423 -9638
rect 41467 -9682 41523 -9638
rect 41567 -9682 41623 -9638
rect 41667 -9682 41723 -9638
rect 41767 -9682 41823 -9638
rect 41867 -9682 41923 -9638
rect 41967 -9682 42023 -9638
rect 42067 -9682 42123 -9638
rect 42167 -9682 42223 -9638
rect 42267 -9682 42323 -9638
rect 42367 -9682 42423 -9638
rect 42467 -9682 42523 -9638
rect 42567 -9682 42623 -9638
rect 42667 -9682 42723 -9638
rect 42767 -9682 43223 -9638
rect 43267 -9682 43323 -9638
rect 43367 -9682 43423 -9638
rect 43467 -9682 43523 -9638
rect 43567 -9682 43623 -9638
rect 43667 -9682 43723 -9638
rect 43767 -9682 43823 -9638
rect 43867 -9682 43923 -9638
rect 43967 -9682 44023 -9638
rect 44067 -9682 44123 -9638
rect 44167 -9682 44223 -9638
rect 44267 -9682 44323 -9638
rect 44367 -9682 44423 -9638
rect 44467 -9682 44523 -9638
rect 44567 -9682 44623 -9638
rect 44667 -9682 44723 -9638
rect 44767 -9682 50994 -9638
rect 34207 -9738 50994 -9682
rect 34207 -9782 37223 -9738
rect 37267 -9782 37323 -9738
rect 37367 -9782 37423 -9738
rect 37467 -9782 37523 -9738
rect 37567 -9782 37623 -9738
rect 37667 -9782 37723 -9738
rect 37767 -9782 37823 -9738
rect 37867 -9782 37923 -9738
rect 37967 -9782 38023 -9738
rect 38067 -9782 38123 -9738
rect 38167 -9782 38223 -9738
rect 38267 -9782 38323 -9738
rect 38367 -9782 38423 -9738
rect 38467 -9782 38523 -9738
rect 38567 -9782 38623 -9738
rect 38667 -9782 38723 -9738
rect 38767 -9782 39223 -9738
rect 39267 -9782 39323 -9738
rect 39367 -9782 39423 -9738
rect 39467 -9782 39523 -9738
rect 39567 -9782 39623 -9738
rect 39667 -9782 39723 -9738
rect 39767 -9782 39823 -9738
rect 39867 -9782 39923 -9738
rect 39967 -9782 40023 -9738
rect 40067 -9782 40123 -9738
rect 40167 -9782 40223 -9738
rect 40267 -9782 40323 -9738
rect 40367 -9782 40423 -9738
rect 40467 -9782 40523 -9738
rect 40567 -9782 40623 -9738
rect 40667 -9782 40723 -9738
rect 40767 -9782 41223 -9738
rect 41267 -9782 41323 -9738
rect 41367 -9782 41423 -9738
rect 41467 -9782 41523 -9738
rect 41567 -9782 41623 -9738
rect 41667 -9782 41723 -9738
rect 41767 -9782 41823 -9738
rect 41867 -9782 41923 -9738
rect 41967 -9782 42023 -9738
rect 42067 -9782 42123 -9738
rect 42167 -9782 42223 -9738
rect 42267 -9782 42323 -9738
rect 42367 -9782 42423 -9738
rect 42467 -9782 42523 -9738
rect 42567 -9782 42623 -9738
rect 42667 -9782 42723 -9738
rect 42767 -9782 43223 -9738
rect 43267 -9782 43323 -9738
rect 43367 -9782 43423 -9738
rect 43467 -9782 43523 -9738
rect 43567 -9782 43623 -9738
rect 43667 -9782 43723 -9738
rect 43767 -9782 43823 -9738
rect 43867 -9782 43923 -9738
rect 43967 -9782 44023 -9738
rect 44067 -9782 44123 -9738
rect 44167 -9782 44223 -9738
rect 44267 -9782 44323 -9738
rect 44367 -9782 44423 -9738
rect 44467 -9782 44523 -9738
rect 44567 -9782 44623 -9738
rect 44667 -9782 44723 -9738
rect 44767 -9782 50994 -9738
rect 34207 -9838 50994 -9782
rect 34207 -9882 37223 -9838
rect 37267 -9882 37323 -9838
rect 37367 -9882 37423 -9838
rect 37467 -9882 37523 -9838
rect 37567 -9882 37623 -9838
rect 37667 -9882 37723 -9838
rect 37767 -9882 37823 -9838
rect 37867 -9882 37923 -9838
rect 37967 -9882 38023 -9838
rect 38067 -9882 38123 -9838
rect 38167 -9882 38223 -9838
rect 38267 -9882 38323 -9838
rect 38367 -9882 38423 -9838
rect 38467 -9882 38523 -9838
rect 38567 -9882 38623 -9838
rect 38667 -9882 38723 -9838
rect 38767 -9882 39223 -9838
rect 39267 -9882 39323 -9838
rect 39367 -9882 39423 -9838
rect 39467 -9882 39523 -9838
rect 39567 -9882 39623 -9838
rect 39667 -9882 39723 -9838
rect 39767 -9882 39823 -9838
rect 39867 -9882 39923 -9838
rect 39967 -9882 40023 -9838
rect 40067 -9882 40123 -9838
rect 40167 -9882 40223 -9838
rect 40267 -9882 40323 -9838
rect 40367 -9882 40423 -9838
rect 40467 -9882 40523 -9838
rect 40567 -9882 40623 -9838
rect 40667 -9882 40723 -9838
rect 40767 -9882 41223 -9838
rect 41267 -9882 41323 -9838
rect 41367 -9882 41423 -9838
rect 41467 -9882 41523 -9838
rect 41567 -9882 41623 -9838
rect 41667 -9882 41723 -9838
rect 41767 -9882 41823 -9838
rect 41867 -9882 41923 -9838
rect 41967 -9882 42023 -9838
rect 42067 -9882 42123 -9838
rect 42167 -9882 42223 -9838
rect 42267 -9882 42323 -9838
rect 42367 -9882 42423 -9838
rect 42467 -9882 42523 -9838
rect 42567 -9882 42623 -9838
rect 42667 -9882 42723 -9838
rect 42767 -9882 43223 -9838
rect 43267 -9882 43323 -9838
rect 43367 -9882 43423 -9838
rect 43467 -9882 43523 -9838
rect 43567 -9882 43623 -9838
rect 43667 -9882 43723 -9838
rect 43767 -9882 43823 -9838
rect 43867 -9882 43923 -9838
rect 43967 -9882 44023 -9838
rect 44067 -9882 44123 -9838
rect 44167 -9882 44223 -9838
rect 44267 -9882 44323 -9838
rect 44367 -9882 44423 -9838
rect 44467 -9882 44523 -9838
rect 44567 -9882 44623 -9838
rect 44667 -9882 44723 -9838
rect 44767 -9882 50994 -9838
rect 34207 -9938 50994 -9882
rect 34207 -9982 37223 -9938
rect 37267 -9982 37323 -9938
rect 37367 -9982 37423 -9938
rect 37467 -9982 37523 -9938
rect 37567 -9982 37623 -9938
rect 37667 -9982 37723 -9938
rect 37767 -9982 37823 -9938
rect 37867 -9982 37923 -9938
rect 37967 -9982 38023 -9938
rect 38067 -9982 38123 -9938
rect 38167 -9982 38223 -9938
rect 38267 -9982 38323 -9938
rect 38367 -9982 38423 -9938
rect 38467 -9982 38523 -9938
rect 38567 -9982 38623 -9938
rect 38667 -9982 38723 -9938
rect 38767 -9982 39223 -9938
rect 39267 -9982 39323 -9938
rect 39367 -9982 39423 -9938
rect 39467 -9982 39523 -9938
rect 39567 -9982 39623 -9938
rect 39667 -9982 39723 -9938
rect 39767 -9982 39823 -9938
rect 39867 -9982 39923 -9938
rect 39967 -9982 40023 -9938
rect 40067 -9982 40123 -9938
rect 40167 -9982 40223 -9938
rect 40267 -9982 40323 -9938
rect 40367 -9982 40423 -9938
rect 40467 -9982 40523 -9938
rect 40567 -9982 40623 -9938
rect 40667 -9982 40723 -9938
rect 40767 -9982 41223 -9938
rect 41267 -9982 41323 -9938
rect 41367 -9982 41423 -9938
rect 41467 -9982 41523 -9938
rect 41567 -9982 41623 -9938
rect 41667 -9982 41723 -9938
rect 41767 -9982 41823 -9938
rect 41867 -9982 41923 -9938
rect 41967 -9982 42023 -9938
rect 42067 -9982 42123 -9938
rect 42167 -9982 42223 -9938
rect 42267 -9982 42323 -9938
rect 42367 -9982 42423 -9938
rect 42467 -9982 42523 -9938
rect 42567 -9982 42623 -9938
rect 42667 -9982 42723 -9938
rect 42767 -9982 43223 -9938
rect 43267 -9982 43323 -9938
rect 43367 -9982 43423 -9938
rect 43467 -9982 43523 -9938
rect 43567 -9982 43623 -9938
rect 43667 -9982 43723 -9938
rect 43767 -9982 43823 -9938
rect 43867 -9982 43923 -9938
rect 43967 -9982 44023 -9938
rect 44067 -9982 44123 -9938
rect 44167 -9982 44223 -9938
rect 44267 -9982 44323 -9938
rect 44367 -9982 44423 -9938
rect 44467 -9982 44523 -9938
rect 44567 -9982 44623 -9938
rect 44667 -9982 44723 -9938
rect 44767 -9982 50994 -9938
rect 34207 -10038 50994 -9982
rect 34207 -10082 37223 -10038
rect 37267 -10082 37323 -10038
rect 37367 -10082 37423 -10038
rect 37467 -10082 37523 -10038
rect 37567 -10082 37623 -10038
rect 37667 -10082 37723 -10038
rect 37767 -10082 37823 -10038
rect 37867 -10082 37923 -10038
rect 37967 -10082 38023 -10038
rect 38067 -10082 38123 -10038
rect 38167 -10082 38223 -10038
rect 38267 -10082 38323 -10038
rect 38367 -10082 38423 -10038
rect 38467 -10082 38523 -10038
rect 38567 -10082 38623 -10038
rect 38667 -10082 38723 -10038
rect 38767 -10082 39223 -10038
rect 39267 -10082 39323 -10038
rect 39367 -10082 39423 -10038
rect 39467 -10082 39523 -10038
rect 39567 -10082 39623 -10038
rect 39667 -10082 39723 -10038
rect 39767 -10082 39823 -10038
rect 39867 -10082 39923 -10038
rect 39967 -10082 40023 -10038
rect 40067 -10082 40123 -10038
rect 40167 -10082 40223 -10038
rect 40267 -10082 40323 -10038
rect 40367 -10082 40423 -10038
rect 40467 -10082 40523 -10038
rect 40567 -10082 40623 -10038
rect 40667 -10082 40723 -10038
rect 40767 -10082 41223 -10038
rect 41267 -10082 41323 -10038
rect 41367 -10082 41423 -10038
rect 41467 -10082 41523 -10038
rect 41567 -10082 41623 -10038
rect 41667 -10082 41723 -10038
rect 41767 -10082 41823 -10038
rect 41867 -10082 41923 -10038
rect 41967 -10082 42023 -10038
rect 42067 -10082 42123 -10038
rect 42167 -10082 42223 -10038
rect 42267 -10082 42323 -10038
rect 42367 -10082 42423 -10038
rect 42467 -10082 42523 -10038
rect 42567 -10082 42623 -10038
rect 42667 -10082 42723 -10038
rect 42767 -10082 43223 -10038
rect 43267 -10082 43323 -10038
rect 43367 -10082 43423 -10038
rect 43467 -10082 43523 -10038
rect 43567 -10082 43623 -10038
rect 43667 -10082 43723 -10038
rect 43767 -10082 43823 -10038
rect 43867 -10082 43923 -10038
rect 43967 -10082 44023 -10038
rect 44067 -10082 44123 -10038
rect 44167 -10082 44223 -10038
rect 44267 -10082 44323 -10038
rect 44367 -10082 44423 -10038
rect 44467 -10082 44523 -10038
rect 44567 -10082 44623 -10038
rect 44667 -10082 44723 -10038
rect 44767 -10082 50994 -10038
rect 34207 -10138 50994 -10082
rect 34207 -10182 37223 -10138
rect 37267 -10182 37323 -10138
rect 37367 -10182 37423 -10138
rect 37467 -10182 37523 -10138
rect 37567 -10182 37623 -10138
rect 37667 -10182 37723 -10138
rect 37767 -10182 37823 -10138
rect 37867 -10182 37923 -10138
rect 37967 -10182 38023 -10138
rect 38067 -10182 38123 -10138
rect 38167 -10182 38223 -10138
rect 38267 -10182 38323 -10138
rect 38367 -10182 38423 -10138
rect 38467 -10182 38523 -10138
rect 38567 -10182 38623 -10138
rect 38667 -10182 38723 -10138
rect 38767 -10182 39223 -10138
rect 39267 -10182 39323 -10138
rect 39367 -10182 39423 -10138
rect 39467 -10182 39523 -10138
rect 39567 -10182 39623 -10138
rect 39667 -10182 39723 -10138
rect 39767 -10182 39823 -10138
rect 39867 -10182 39923 -10138
rect 39967 -10182 40023 -10138
rect 40067 -10182 40123 -10138
rect 40167 -10182 40223 -10138
rect 40267 -10182 40323 -10138
rect 40367 -10182 40423 -10138
rect 40467 -10182 40523 -10138
rect 40567 -10182 40623 -10138
rect 40667 -10182 40723 -10138
rect 40767 -10182 41223 -10138
rect 41267 -10182 41323 -10138
rect 41367 -10182 41423 -10138
rect 41467 -10182 41523 -10138
rect 41567 -10182 41623 -10138
rect 41667 -10182 41723 -10138
rect 41767 -10182 41823 -10138
rect 41867 -10182 41923 -10138
rect 41967 -10182 42023 -10138
rect 42067 -10182 42123 -10138
rect 42167 -10182 42223 -10138
rect 42267 -10182 42323 -10138
rect 42367 -10182 42423 -10138
rect 42467 -10182 42523 -10138
rect 42567 -10182 42623 -10138
rect 42667 -10182 42723 -10138
rect 42767 -10182 43223 -10138
rect 43267 -10182 43323 -10138
rect 43367 -10182 43423 -10138
rect 43467 -10182 43523 -10138
rect 43567 -10182 43623 -10138
rect 43667 -10182 43723 -10138
rect 43767 -10182 43823 -10138
rect 43867 -10182 43923 -10138
rect 43967 -10182 44023 -10138
rect 44067 -10182 44123 -10138
rect 44167 -10182 44223 -10138
rect 44267 -10182 44323 -10138
rect 44367 -10182 44423 -10138
rect 44467 -10182 44523 -10138
rect 44567 -10182 44623 -10138
rect 44667 -10182 44723 -10138
rect 44767 -10182 50994 -10138
rect 34207 -10238 50994 -10182
rect 34207 -10282 37223 -10238
rect 37267 -10282 37323 -10238
rect 37367 -10282 37423 -10238
rect 37467 -10282 37523 -10238
rect 37567 -10282 37623 -10238
rect 37667 -10282 37723 -10238
rect 37767 -10282 37823 -10238
rect 37867 -10282 37923 -10238
rect 37967 -10282 38023 -10238
rect 38067 -10282 38123 -10238
rect 38167 -10282 38223 -10238
rect 38267 -10282 38323 -10238
rect 38367 -10282 38423 -10238
rect 38467 -10282 38523 -10238
rect 38567 -10282 38623 -10238
rect 38667 -10282 38723 -10238
rect 38767 -10282 39223 -10238
rect 39267 -10282 39323 -10238
rect 39367 -10282 39423 -10238
rect 39467 -10282 39523 -10238
rect 39567 -10282 39623 -10238
rect 39667 -10282 39723 -10238
rect 39767 -10282 39823 -10238
rect 39867 -10282 39923 -10238
rect 39967 -10282 40023 -10238
rect 40067 -10282 40123 -10238
rect 40167 -10282 40223 -10238
rect 40267 -10282 40323 -10238
rect 40367 -10282 40423 -10238
rect 40467 -10282 40523 -10238
rect 40567 -10282 40623 -10238
rect 40667 -10282 40723 -10238
rect 40767 -10282 41223 -10238
rect 41267 -10282 41323 -10238
rect 41367 -10282 41423 -10238
rect 41467 -10282 41523 -10238
rect 41567 -10282 41623 -10238
rect 41667 -10282 41723 -10238
rect 41767 -10282 41823 -10238
rect 41867 -10282 41923 -10238
rect 41967 -10282 42023 -10238
rect 42067 -10282 42123 -10238
rect 42167 -10282 42223 -10238
rect 42267 -10282 42323 -10238
rect 42367 -10282 42423 -10238
rect 42467 -10282 42523 -10238
rect 42567 -10282 42623 -10238
rect 42667 -10282 42723 -10238
rect 42767 -10282 43223 -10238
rect 43267 -10282 43323 -10238
rect 43367 -10282 43423 -10238
rect 43467 -10282 43523 -10238
rect 43567 -10282 43623 -10238
rect 43667 -10282 43723 -10238
rect 43767 -10282 43823 -10238
rect 43867 -10282 43923 -10238
rect 43967 -10282 44023 -10238
rect 44067 -10282 44123 -10238
rect 44167 -10282 44223 -10238
rect 44267 -10282 44323 -10238
rect 44367 -10282 44423 -10238
rect 44467 -10282 44523 -10238
rect 44567 -10282 44623 -10238
rect 44667 -10282 44723 -10238
rect 44767 -10282 50994 -10238
rect 34207 -10338 50994 -10282
rect 34207 -10382 37223 -10338
rect 37267 -10382 37323 -10338
rect 37367 -10382 37423 -10338
rect 37467 -10382 37523 -10338
rect 37567 -10382 37623 -10338
rect 37667 -10382 37723 -10338
rect 37767 -10382 37823 -10338
rect 37867 -10382 37923 -10338
rect 37967 -10382 38023 -10338
rect 38067 -10382 38123 -10338
rect 38167 -10382 38223 -10338
rect 38267 -10382 38323 -10338
rect 38367 -10382 38423 -10338
rect 38467 -10382 38523 -10338
rect 38567 -10382 38623 -10338
rect 38667 -10382 38723 -10338
rect 38767 -10382 39223 -10338
rect 39267 -10382 39323 -10338
rect 39367 -10382 39423 -10338
rect 39467 -10382 39523 -10338
rect 39567 -10382 39623 -10338
rect 39667 -10382 39723 -10338
rect 39767 -10382 39823 -10338
rect 39867 -10382 39923 -10338
rect 39967 -10382 40023 -10338
rect 40067 -10382 40123 -10338
rect 40167 -10382 40223 -10338
rect 40267 -10382 40323 -10338
rect 40367 -10382 40423 -10338
rect 40467 -10382 40523 -10338
rect 40567 -10382 40623 -10338
rect 40667 -10382 40723 -10338
rect 40767 -10382 41223 -10338
rect 41267 -10382 41323 -10338
rect 41367 -10382 41423 -10338
rect 41467 -10382 41523 -10338
rect 41567 -10382 41623 -10338
rect 41667 -10382 41723 -10338
rect 41767 -10382 41823 -10338
rect 41867 -10382 41923 -10338
rect 41967 -10382 42023 -10338
rect 42067 -10382 42123 -10338
rect 42167 -10382 42223 -10338
rect 42267 -10382 42323 -10338
rect 42367 -10382 42423 -10338
rect 42467 -10382 42523 -10338
rect 42567 -10382 42623 -10338
rect 42667 -10382 42723 -10338
rect 42767 -10382 43223 -10338
rect 43267 -10382 43323 -10338
rect 43367 -10382 43423 -10338
rect 43467 -10382 43523 -10338
rect 43567 -10382 43623 -10338
rect 43667 -10382 43723 -10338
rect 43767 -10382 43823 -10338
rect 43867 -10382 43923 -10338
rect 43967 -10382 44023 -10338
rect 44067 -10382 44123 -10338
rect 44167 -10382 44223 -10338
rect 44267 -10382 44323 -10338
rect 44367 -10382 44423 -10338
rect 44467 -10382 44523 -10338
rect 44567 -10382 44623 -10338
rect 44667 -10382 44723 -10338
rect 44767 -10382 50994 -10338
rect 34207 -10438 50994 -10382
rect 34207 -10482 37223 -10438
rect 37267 -10482 37323 -10438
rect 37367 -10482 37423 -10438
rect 37467 -10482 37523 -10438
rect 37567 -10482 37623 -10438
rect 37667 -10482 37723 -10438
rect 37767 -10482 37823 -10438
rect 37867 -10482 37923 -10438
rect 37967 -10482 38023 -10438
rect 38067 -10482 38123 -10438
rect 38167 -10482 38223 -10438
rect 38267 -10482 38323 -10438
rect 38367 -10482 38423 -10438
rect 38467 -10482 38523 -10438
rect 38567 -10482 38623 -10438
rect 38667 -10482 38723 -10438
rect 38767 -10482 39223 -10438
rect 39267 -10482 39323 -10438
rect 39367 -10482 39423 -10438
rect 39467 -10482 39523 -10438
rect 39567 -10482 39623 -10438
rect 39667 -10482 39723 -10438
rect 39767 -10482 39823 -10438
rect 39867 -10482 39923 -10438
rect 39967 -10482 40023 -10438
rect 40067 -10482 40123 -10438
rect 40167 -10482 40223 -10438
rect 40267 -10482 40323 -10438
rect 40367 -10482 40423 -10438
rect 40467 -10482 40523 -10438
rect 40567 -10482 40623 -10438
rect 40667 -10482 40723 -10438
rect 40767 -10482 41223 -10438
rect 41267 -10482 41323 -10438
rect 41367 -10482 41423 -10438
rect 41467 -10482 41523 -10438
rect 41567 -10482 41623 -10438
rect 41667 -10482 41723 -10438
rect 41767 -10482 41823 -10438
rect 41867 -10482 41923 -10438
rect 41967 -10482 42023 -10438
rect 42067 -10482 42123 -10438
rect 42167 -10482 42223 -10438
rect 42267 -10482 42323 -10438
rect 42367 -10482 42423 -10438
rect 42467 -10482 42523 -10438
rect 42567 -10482 42623 -10438
rect 42667 -10482 42723 -10438
rect 42767 -10482 43223 -10438
rect 43267 -10482 43323 -10438
rect 43367 -10482 43423 -10438
rect 43467 -10482 43523 -10438
rect 43567 -10482 43623 -10438
rect 43667 -10482 43723 -10438
rect 43767 -10482 43823 -10438
rect 43867 -10482 43923 -10438
rect 43967 -10482 44023 -10438
rect 44067 -10482 44123 -10438
rect 44167 -10482 44223 -10438
rect 44267 -10482 44323 -10438
rect 44367 -10482 44423 -10438
rect 44467 -10482 44523 -10438
rect 44567 -10482 44623 -10438
rect 44667 -10482 44723 -10438
rect 44767 -10482 50994 -10438
rect 34207 -10538 50994 -10482
rect 34207 -10582 37223 -10538
rect 37267 -10582 37323 -10538
rect 37367 -10582 37423 -10538
rect 37467 -10582 37523 -10538
rect 37567 -10582 37623 -10538
rect 37667 -10582 37723 -10538
rect 37767 -10582 37823 -10538
rect 37867 -10582 37923 -10538
rect 37967 -10582 38023 -10538
rect 38067 -10582 38123 -10538
rect 38167 -10582 38223 -10538
rect 38267 -10582 38323 -10538
rect 38367 -10582 38423 -10538
rect 38467 -10582 38523 -10538
rect 38567 -10582 38623 -10538
rect 38667 -10582 38723 -10538
rect 38767 -10582 39223 -10538
rect 39267 -10582 39323 -10538
rect 39367 -10582 39423 -10538
rect 39467 -10582 39523 -10538
rect 39567 -10582 39623 -10538
rect 39667 -10582 39723 -10538
rect 39767 -10582 39823 -10538
rect 39867 -10582 39923 -10538
rect 39967 -10582 40023 -10538
rect 40067 -10582 40123 -10538
rect 40167 -10582 40223 -10538
rect 40267 -10582 40323 -10538
rect 40367 -10582 40423 -10538
rect 40467 -10582 40523 -10538
rect 40567 -10582 40623 -10538
rect 40667 -10582 40723 -10538
rect 40767 -10582 41223 -10538
rect 41267 -10582 41323 -10538
rect 41367 -10582 41423 -10538
rect 41467 -10582 41523 -10538
rect 41567 -10582 41623 -10538
rect 41667 -10582 41723 -10538
rect 41767 -10582 41823 -10538
rect 41867 -10582 41923 -10538
rect 41967 -10582 42023 -10538
rect 42067 -10582 42123 -10538
rect 42167 -10582 42223 -10538
rect 42267 -10582 42323 -10538
rect 42367 -10582 42423 -10538
rect 42467 -10582 42523 -10538
rect 42567 -10582 42623 -10538
rect 42667 -10582 42723 -10538
rect 42767 -10582 43223 -10538
rect 43267 -10582 43323 -10538
rect 43367 -10582 43423 -10538
rect 43467 -10582 43523 -10538
rect 43567 -10582 43623 -10538
rect 43667 -10582 43723 -10538
rect 43767 -10582 43823 -10538
rect 43867 -10582 43923 -10538
rect 43967 -10582 44023 -10538
rect 44067 -10582 44123 -10538
rect 44167 -10582 44223 -10538
rect 44267 -10582 44323 -10538
rect 44367 -10582 44423 -10538
rect 44467 -10582 44523 -10538
rect 44567 -10582 44623 -10538
rect 44667 -10582 44723 -10538
rect 44767 -10582 50994 -10538
rect 34207 -10638 50994 -10582
rect 34207 -10682 37223 -10638
rect 37267 -10682 37323 -10638
rect 37367 -10682 37423 -10638
rect 37467 -10682 37523 -10638
rect 37567 -10682 37623 -10638
rect 37667 -10682 37723 -10638
rect 37767 -10682 37823 -10638
rect 37867 -10682 37923 -10638
rect 37967 -10682 38023 -10638
rect 38067 -10682 38123 -10638
rect 38167 -10682 38223 -10638
rect 38267 -10682 38323 -10638
rect 38367 -10682 38423 -10638
rect 38467 -10682 38523 -10638
rect 38567 -10682 38623 -10638
rect 38667 -10682 38723 -10638
rect 38767 -10682 39223 -10638
rect 39267 -10682 39323 -10638
rect 39367 -10682 39423 -10638
rect 39467 -10682 39523 -10638
rect 39567 -10682 39623 -10638
rect 39667 -10682 39723 -10638
rect 39767 -10682 39823 -10638
rect 39867 -10682 39923 -10638
rect 39967 -10682 40023 -10638
rect 40067 -10682 40123 -10638
rect 40167 -10682 40223 -10638
rect 40267 -10682 40323 -10638
rect 40367 -10682 40423 -10638
rect 40467 -10682 40523 -10638
rect 40567 -10682 40623 -10638
rect 40667 -10682 40723 -10638
rect 40767 -10682 41223 -10638
rect 41267 -10682 41323 -10638
rect 41367 -10682 41423 -10638
rect 41467 -10682 41523 -10638
rect 41567 -10682 41623 -10638
rect 41667 -10682 41723 -10638
rect 41767 -10682 41823 -10638
rect 41867 -10682 41923 -10638
rect 41967 -10682 42023 -10638
rect 42067 -10682 42123 -10638
rect 42167 -10682 42223 -10638
rect 42267 -10682 42323 -10638
rect 42367 -10682 42423 -10638
rect 42467 -10682 42523 -10638
rect 42567 -10682 42623 -10638
rect 42667 -10682 42723 -10638
rect 42767 -10682 43223 -10638
rect 43267 -10682 43323 -10638
rect 43367 -10682 43423 -10638
rect 43467 -10682 43523 -10638
rect 43567 -10682 43623 -10638
rect 43667 -10682 43723 -10638
rect 43767 -10682 43823 -10638
rect 43867 -10682 43923 -10638
rect 43967 -10682 44023 -10638
rect 44067 -10682 44123 -10638
rect 44167 -10682 44223 -10638
rect 44267 -10682 44323 -10638
rect 44367 -10682 44423 -10638
rect 44467 -10682 44523 -10638
rect 44567 -10682 44623 -10638
rect 44667 -10682 44723 -10638
rect 44767 -10682 50994 -10638
rect 34207 -10738 50994 -10682
rect 34207 -10782 37223 -10738
rect 37267 -10782 37323 -10738
rect 37367 -10782 37423 -10738
rect 37467 -10782 37523 -10738
rect 37567 -10782 37623 -10738
rect 37667 -10782 37723 -10738
rect 37767 -10782 37823 -10738
rect 37867 -10782 37923 -10738
rect 37967 -10782 38023 -10738
rect 38067 -10782 38123 -10738
rect 38167 -10782 38223 -10738
rect 38267 -10782 38323 -10738
rect 38367 -10782 38423 -10738
rect 38467 -10782 38523 -10738
rect 38567 -10782 38623 -10738
rect 38667 -10782 38723 -10738
rect 38767 -10782 39223 -10738
rect 39267 -10782 39323 -10738
rect 39367 -10782 39423 -10738
rect 39467 -10782 39523 -10738
rect 39567 -10782 39623 -10738
rect 39667 -10782 39723 -10738
rect 39767 -10782 39823 -10738
rect 39867 -10782 39923 -10738
rect 39967 -10782 40023 -10738
rect 40067 -10782 40123 -10738
rect 40167 -10782 40223 -10738
rect 40267 -10782 40323 -10738
rect 40367 -10782 40423 -10738
rect 40467 -10782 40523 -10738
rect 40567 -10782 40623 -10738
rect 40667 -10782 40723 -10738
rect 40767 -10782 41223 -10738
rect 41267 -10782 41323 -10738
rect 41367 -10782 41423 -10738
rect 41467 -10782 41523 -10738
rect 41567 -10782 41623 -10738
rect 41667 -10782 41723 -10738
rect 41767 -10782 41823 -10738
rect 41867 -10782 41923 -10738
rect 41967 -10782 42023 -10738
rect 42067 -10782 42123 -10738
rect 42167 -10782 42223 -10738
rect 42267 -10782 42323 -10738
rect 42367 -10782 42423 -10738
rect 42467 -10782 42523 -10738
rect 42567 -10782 42623 -10738
rect 42667 -10782 42723 -10738
rect 42767 -10782 43223 -10738
rect 43267 -10782 43323 -10738
rect 43367 -10782 43423 -10738
rect 43467 -10782 43523 -10738
rect 43567 -10782 43623 -10738
rect 43667 -10782 43723 -10738
rect 43767 -10782 43823 -10738
rect 43867 -10782 43923 -10738
rect 43967 -10782 44023 -10738
rect 44067 -10782 44123 -10738
rect 44167 -10782 44223 -10738
rect 44267 -10782 44323 -10738
rect 44367 -10782 44423 -10738
rect 44467 -10782 44523 -10738
rect 44567 -10782 44623 -10738
rect 44667 -10782 44723 -10738
rect 44767 -10782 50994 -10738
rect 34207 -10838 50994 -10782
rect 34207 -10882 37223 -10838
rect 37267 -10882 37323 -10838
rect 37367 -10882 37423 -10838
rect 37467 -10882 37523 -10838
rect 37567 -10882 37623 -10838
rect 37667 -10882 37723 -10838
rect 37767 -10882 37823 -10838
rect 37867 -10882 37923 -10838
rect 37967 -10882 38023 -10838
rect 38067 -10882 38123 -10838
rect 38167 -10882 38223 -10838
rect 38267 -10882 38323 -10838
rect 38367 -10882 38423 -10838
rect 38467 -10882 38523 -10838
rect 38567 -10882 38623 -10838
rect 38667 -10882 38723 -10838
rect 38767 -10882 39223 -10838
rect 39267 -10882 39323 -10838
rect 39367 -10882 39423 -10838
rect 39467 -10882 39523 -10838
rect 39567 -10882 39623 -10838
rect 39667 -10882 39723 -10838
rect 39767 -10882 39823 -10838
rect 39867 -10882 39923 -10838
rect 39967 -10882 40023 -10838
rect 40067 -10882 40123 -10838
rect 40167 -10882 40223 -10838
rect 40267 -10882 40323 -10838
rect 40367 -10882 40423 -10838
rect 40467 -10882 40523 -10838
rect 40567 -10882 40623 -10838
rect 40667 -10882 40723 -10838
rect 40767 -10882 41223 -10838
rect 41267 -10882 41323 -10838
rect 41367 -10882 41423 -10838
rect 41467 -10882 41523 -10838
rect 41567 -10882 41623 -10838
rect 41667 -10882 41723 -10838
rect 41767 -10882 41823 -10838
rect 41867 -10882 41923 -10838
rect 41967 -10882 42023 -10838
rect 42067 -10882 42123 -10838
rect 42167 -10882 42223 -10838
rect 42267 -10882 42323 -10838
rect 42367 -10882 42423 -10838
rect 42467 -10882 42523 -10838
rect 42567 -10882 42623 -10838
rect 42667 -10882 42723 -10838
rect 42767 -10882 43223 -10838
rect 43267 -10882 43323 -10838
rect 43367 -10882 43423 -10838
rect 43467 -10882 43523 -10838
rect 43567 -10882 43623 -10838
rect 43667 -10882 43723 -10838
rect 43767 -10882 43823 -10838
rect 43867 -10882 43923 -10838
rect 43967 -10882 44023 -10838
rect 44067 -10882 44123 -10838
rect 44167 -10882 44223 -10838
rect 44267 -10882 44323 -10838
rect 44367 -10882 44423 -10838
rect 44467 -10882 44523 -10838
rect 44567 -10882 44623 -10838
rect 44667 -10882 44723 -10838
rect 44767 -10882 50994 -10838
rect 34207 -10938 50994 -10882
rect 34207 -10982 37223 -10938
rect 37267 -10982 37323 -10938
rect 37367 -10982 37423 -10938
rect 37467 -10982 37523 -10938
rect 37567 -10982 37623 -10938
rect 37667 -10982 37723 -10938
rect 37767 -10982 37823 -10938
rect 37867 -10982 37923 -10938
rect 37967 -10982 38023 -10938
rect 38067 -10982 38123 -10938
rect 38167 -10982 38223 -10938
rect 38267 -10982 38323 -10938
rect 38367 -10982 38423 -10938
rect 38467 -10982 38523 -10938
rect 38567 -10982 38623 -10938
rect 38667 -10982 38723 -10938
rect 38767 -10982 39223 -10938
rect 39267 -10982 39323 -10938
rect 39367 -10982 39423 -10938
rect 39467 -10982 39523 -10938
rect 39567 -10982 39623 -10938
rect 39667 -10982 39723 -10938
rect 39767 -10982 39823 -10938
rect 39867 -10982 39923 -10938
rect 39967 -10982 40023 -10938
rect 40067 -10982 40123 -10938
rect 40167 -10982 40223 -10938
rect 40267 -10982 40323 -10938
rect 40367 -10982 40423 -10938
rect 40467 -10982 40523 -10938
rect 40567 -10982 40623 -10938
rect 40667 -10982 40723 -10938
rect 40767 -10982 41223 -10938
rect 41267 -10982 41323 -10938
rect 41367 -10982 41423 -10938
rect 41467 -10982 41523 -10938
rect 41567 -10982 41623 -10938
rect 41667 -10982 41723 -10938
rect 41767 -10982 41823 -10938
rect 41867 -10982 41923 -10938
rect 41967 -10982 42023 -10938
rect 42067 -10982 42123 -10938
rect 42167 -10982 42223 -10938
rect 42267 -10982 42323 -10938
rect 42367 -10982 42423 -10938
rect 42467 -10982 42523 -10938
rect 42567 -10982 42623 -10938
rect 42667 -10982 42723 -10938
rect 42767 -10982 43223 -10938
rect 43267 -10982 43323 -10938
rect 43367 -10982 43423 -10938
rect 43467 -10982 43523 -10938
rect 43567 -10982 43623 -10938
rect 43667 -10982 43723 -10938
rect 43767 -10982 43823 -10938
rect 43867 -10982 43923 -10938
rect 43967 -10982 44023 -10938
rect 44067 -10982 44123 -10938
rect 44167 -10982 44223 -10938
rect 44267 -10982 44323 -10938
rect 44367 -10982 44423 -10938
rect 44467 -10982 44523 -10938
rect 44567 -10982 44623 -10938
rect 44667 -10982 44723 -10938
rect 44767 -10982 50994 -10938
rect 34207 -11038 50994 -10982
rect 34207 -11082 37223 -11038
rect 37267 -11082 37323 -11038
rect 37367 -11082 37423 -11038
rect 37467 -11082 37523 -11038
rect 37567 -11082 37623 -11038
rect 37667 -11082 37723 -11038
rect 37767 -11082 37823 -11038
rect 37867 -11082 37923 -11038
rect 37967 -11082 38023 -11038
rect 38067 -11082 38123 -11038
rect 38167 -11082 38223 -11038
rect 38267 -11082 38323 -11038
rect 38367 -11082 38423 -11038
rect 38467 -11082 38523 -11038
rect 38567 -11082 38623 -11038
rect 38667 -11082 38723 -11038
rect 38767 -11082 39223 -11038
rect 39267 -11082 39323 -11038
rect 39367 -11082 39423 -11038
rect 39467 -11082 39523 -11038
rect 39567 -11082 39623 -11038
rect 39667 -11082 39723 -11038
rect 39767 -11082 39823 -11038
rect 39867 -11082 39923 -11038
rect 39967 -11082 40023 -11038
rect 40067 -11082 40123 -11038
rect 40167 -11082 40223 -11038
rect 40267 -11082 40323 -11038
rect 40367 -11082 40423 -11038
rect 40467 -11082 40523 -11038
rect 40567 -11082 40623 -11038
rect 40667 -11082 40723 -11038
rect 40767 -11082 41223 -11038
rect 41267 -11082 41323 -11038
rect 41367 -11082 41423 -11038
rect 41467 -11082 41523 -11038
rect 41567 -11082 41623 -11038
rect 41667 -11082 41723 -11038
rect 41767 -11082 41823 -11038
rect 41867 -11082 41923 -11038
rect 41967 -11082 42023 -11038
rect 42067 -11082 42123 -11038
rect 42167 -11082 42223 -11038
rect 42267 -11082 42323 -11038
rect 42367 -11082 42423 -11038
rect 42467 -11082 42523 -11038
rect 42567 -11082 42623 -11038
rect 42667 -11082 42723 -11038
rect 42767 -11082 43223 -11038
rect 43267 -11082 43323 -11038
rect 43367 -11082 43423 -11038
rect 43467 -11082 43523 -11038
rect 43567 -11082 43623 -11038
rect 43667 -11082 43723 -11038
rect 43767 -11082 43823 -11038
rect 43867 -11082 43923 -11038
rect 43967 -11082 44023 -11038
rect 44067 -11082 44123 -11038
rect 44167 -11082 44223 -11038
rect 44267 -11082 44323 -11038
rect 44367 -11082 44423 -11038
rect 44467 -11082 44523 -11038
rect 44567 -11082 44623 -11038
rect 44667 -11082 44723 -11038
rect 44767 -11082 50994 -11038
rect 34207 -11138 50994 -11082
rect 34207 -11182 37223 -11138
rect 37267 -11182 37323 -11138
rect 37367 -11182 37423 -11138
rect 37467 -11182 37523 -11138
rect 37567 -11182 37623 -11138
rect 37667 -11182 37723 -11138
rect 37767 -11182 37823 -11138
rect 37867 -11182 37923 -11138
rect 37967 -11182 38023 -11138
rect 38067 -11182 38123 -11138
rect 38167 -11182 38223 -11138
rect 38267 -11182 38323 -11138
rect 38367 -11182 38423 -11138
rect 38467 -11182 38523 -11138
rect 38567 -11182 38623 -11138
rect 38667 -11182 38723 -11138
rect 38767 -11182 39223 -11138
rect 39267 -11182 39323 -11138
rect 39367 -11182 39423 -11138
rect 39467 -11182 39523 -11138
rect 39567 -11182 39623 -11138
rect 39667 -11182 39723 -11138
rect 39767 -11182 39823 -11138
rect 39867 -11182 39923 -11138
rect 39967 -11182 40023 -11138
rect 40067 -11182 40123 -11138
rect 40167 -11182 40223 -11138
rect 40267 -11182 40323 -11138
rect 40367 -11182 40423 -11138
rect 40467 -11182 40523 -11138
rect 40567 -11182 40623 -11138
rect 40667 -11182 40723 -11138
rect 40767 -11182 41223 -11138
rect 41267 -11182 41323 -11138
rect 41367 -11182 41423 -11138
rect 41467 -11182 41523 -11138
rect 41567 -11182 41623 -11138
rect 41667 -11182 41723 -11138
rect 41767 -11182 41823 -11138
rect 41867 -11182 41923 -11138
rect 41967 -11182 42023 -11138
rect 42067 -11182 42123 -11138
rect 42167 -11182 42223 -11138
rect 42267 -11182 42323 -11138
rect 42367 -11182 42423 -11138
rect 42467 -11182 42523 -11138
rect 42567 -11182 42623 -11138
rect 42667 -11182 42723 -11138
rect 42767 -11182 43223 -11138
rect 43267 -11182 43323 -11138
rect 43367 -11182 43423 -11138
rect 43467 -11182 43523 -11138
rect 43567 -11182 43623 -11138
rect 43667 -11182 43723 -11138
rect 43767 -11182 43823 -11138
rect 43867 -11182 43923 -11138
rect 43967 -11182 44023 -11138
rect 44067 -11182 44123 -11138
rect 44167 -11182 44223 -11138
rect 44267 -11182 44323 -11138
rect 44367 -11182 44423 -11138
rect 44467 -11182 44523 -11138
rect 44567 -11182 44623 -11138
rect 44667 -11182 44723 -11138
rect 44767 -11182 50994 -11138
rect 34207 -19129 50994 -11182
rect 56492 -19695 58090 794
rect 58502 309 58578 794
rect 58990 309 59066 794
rect 59478 309 59554 794
rect 59966 309 60042 794
rect 60454 309 60530 794
rect 60942 309 61018 794
rect 61430 309 61506 794
rect 61918 309 61994 794
rect 62406 309 62482 794
rect 62894 309 62970 794
rect 63382 309 63458 794
rect 63870 309 63946 794
rect 64358 309 64434 794
rect 64846 309 64922 794
rect 65334 309 65410 794
rect 65822 309 65898 794
rect 66310 309 66386 794
rect 66798 309 66874 794
rect 67286 309 67362 794
rect 67774 309 67850 794
rect 68262 309 68338 794
rect 68750 309 68826 794
rect 69238 309 69314 794
rect 69726 309 69802 794
rect 70214 309 70290 794
rect 70702 309 70778 794
rect 71190 309 71266 794
rect 71678 309 71754 794
rect 72166 309 72242 794
rect 72654 309 72730 794
rect 73142 309 73218 794
rect 73630 309 73706 794
rect 74118 309 74194 794
rect 74606 309 74682 794
rect 75094 309 75170 794
rect 75582 309 75658 794
rect 76070 309 76146 794
rect 76558 309 76634 794
rect 77046 309 77122 794
rect 77534 309 77610 794
rect 78022 309 78098 794
rect 78510 309 78586 794
rect 78998 309 79074 794
rect 79486 309 79562 794
rect 79974 309 80050 794
rect 80462 309 80538 794
rect 80950 309 81026 794
rect 81438 309 81514 794
rect 81926 309 82002 794
rect 82414 309 82490 794
rect 85014 309 85090 794
rect 85502 309 85578 794
rect 85990 309 86066 794
rect 86478 309 86554 794
rect 86966 309 87042 794
rect 87454 309 87530 794
rect 87942 309 88018 794
rect 88430 309 88506 794
rect 88918 309 88994 794
rect 89406 309 89482 794
rect 89894 309 89970 794
rect 90382 309 90458 794
rect 90870 309 90946 794
rect 91358 309 91434 794
rect 91846 309 91922 794
rect 92334 309 92410 794
rect 92822 309 92898 794
rect 93310 309 93386 794
rect 93798 309 93874 794
rect 94286 309 94362 794
rect 94774 309 94850 794
rect 95262 309 95338 794
rect 95750 309 95826 794
rect 96238 309 96314 794
rect 96726 309 96802 794
rect 97214 309 97290 794
rect 97702 309 97778 794
rect 98190 309 98266 794
rect 98678 309 98754 794
rect 99166 309 99242 794
rect 99654 309 99730 794
rect 100142 309 100218 794
rect 100630 309 100706 794
rect 101118 309 101194 794
rect 101606 309 101682 794
rect 102094 309 102170 794
rect 102582 309 102658 794
rect 103070 309 103146 794
rect 103558 309 103634 794
rect 104046 309 104122 794
rect 104534 309 104610 794
rect 105022 309 105098 794
rect 105510 309 105586 794
rect 105998 309 106074 794
rect 106486 309 106562 794
rect 106974 309 107050 794
rect 107462 309 107538 794
rect 107950 309 108026 794
rect 108438 309 108514 794
rect 108926 309 109002 794
rect 109414 309 109490 794
rect 84856 -19695 85090 307
rect 109734 -14975 111646 4125
rect 109734 -17214 178142 -14975
rect 109734 -17445 173611 -17214
rect 109734 -17489 144904 -17445
rect 144948 -17489 145004 -17445
rect 145048 -17489 145104 -17445
rect 145148 -17489 145204 -17445
rect 145248 -17489 145304 -17445
rect 145348 -17489 145404 -17445
rect 145448 -17489 145504 -17445
rect 145548 -17489 145604 -17445
rect 145648 -17489 145704 -17445
rect 145748 -17489 145804 -17445
rect 145848 -17489 145904 -17445
rect 145948 -17489 146004 -17445
rect 146048 -17489 146104 -17445
rect 146148 -17489 146204 -17445
rect 146248 -17489 146304 -17445
rect 146348 -17489 146404 -17445
rect 146448 -17489 146904 -17445
rect 146948 -17489 147004 -17445
rect 147048 -17489 147104 -17445
rect 147148 -17489 147204 -17445
rect 147248 -17489 147304 -17445
rect 147348 -17489 147404 -17445
rect 147448 -17489 147504 -17445
rect 147548 -17489 147604 -17445
rect 147648 -17489 147704 -17445
rect 147748 -17489 147804 -17445
rect 147848 -17489 147904 -17445
rect 147948 -17489 148004 -17445
rect 148048 -17489 148104 -17445
rect 148148 -17489 148204 -17445
rect 148248 -17489 148304 -17445
rect 148348 -17489 148404 -17445
rect 148448 -17489 148904 -17445
rect 148948 -17489 149004 -17445
rect 149048 -17489 149104 -17445
rect 149148 -17489 149204 -17445
rect 149248 -17489 149304 -17445
rect 149348 -17489 149404 -17445
rect 149448 -17489 149504 -17445
rect 149548 -17489 149604 -17445
rect 149648 -17489 149704 -17445
rect 149748 -17489 149804 -17445
rect 149848 -17489 149904 -17445
rect 149948 -17489 150004 -17445
rect 150048 -17489 150104 -17445
rect 150148 -17489 150204 -17445
rect 150248 -17489 150304 -17445
rect 150348 -17489 150404 -17445
rect 150448 -17489 150904 -17445
rect 150948 -17489 151004 -17445
rect 151048 -17489 151104 -17445
rect 151148 -17489 151204 -17445
rect 151248 -17489 151304 -17445
rect 151348 -17489 151404 -17445
rect 151448 -17489 151504 -17445
rect 151548 -17489 151604 -17445
rect 151648 -17489 151704 -17445
rect 151748 -17489 151804 -17445
rect 151848 -17489 151904 -17445
rect 151948 -17489 152004 -17445
rect 152048 -17489 152104 -17445
rect 152148 -17489 152204 -17445
rect 152248 -17489 152304 -17445
rect 152348 -17489 152404 -17445
rect 152448 -17489 173611 -17445
rect 109734 -17545 173611 -17489
rect 109734 -17589 144904 -17545
rect 144948 -17589 145004 -17545
rect 145048 -17589 145104 -17545
rect 145148 -17589 145204 -17545
rect 145248 -17589 145304 -17545
rect 145348 -17589 145404 -17545
rect 145448 -17589 145504 -17545
rect 145548 -17589 145604 -17545
rect 145648 -17589 145704 -17545
rect 145748 -17589 145804 -17545
rect 145848 -17589 145904 -17545
rect 145948 -17589 146004 -17545
rect 146048 -17589 146104 -17545
rect 146148 -17589 146204 -17545
rect 146248 -17589 146304 -17545
rect 146348 -17589 146404 -17545
rect 146448 -17589 146904 -17545
rect 146948 -17589 147004 -17545
rect 147048 -17589 147104 -17545
rect 147148 -17589 147204 -17545
rect 147248 -17589 147304 -17545
rect 147348 -17589 147404 -17545
rect 147448 -17589 147504 -17545
rect 147548 -17589 147604 -17545
rect 147648 -17589 147704 -17545
rect 147748 -17589 147804 -17545
rect 147848 -17589 147904 -17545
rect 147948 -17589 148004 -17545
rect 148048 -17589 148104 -17545
rect 148148 -17589 148204 -17545
rect 148248 -17589 148304 -17545
rect 148348 -17589 148404 -17545
rect 148448 -17589 148904 -17545
rect 148948 -17589 149004 -17545
rect 149048 -17589 149104 -17545
rect 149148 -17589 149204 -17545
rect 149248 -17589 149304 -17545
rect 149348 -17589 149404 -17545
rect 149448 -17589 149504 -17545
rect 149548 -17589 149604 -17545
rect 149648 -17589 149704 -17545
rect 149748 -17589 149804 -17545
rect 149848 -17589 149904 -17545
rect 149948 -17589 150004 -17545
rect 150048 -17589 150104 -17545
rect 150148 -17589 150204 -17545
rect 150248 -17589 150304 -17545
rect 150348 -17589 150404 -17545
rect 150448 -17589 150904 -17545
rect 150948 -17589 151004 -17545
rect 151048 -17589 151104 -17545
rect 151148 -17589 151204 -17545
rect 151248 -17589 151304 -17545
rect 151348 -17589 151404 -17545
rect 151448 -17589 151504 -17545
rect 151548 -17589 151604 -17545
rect 151648 -17589 151704 -17545
rect 151748 -17589 151804 -17545
rect 151848 -17589 151904 -17545
rect 151948 -17589 152004 -17545
rect 152048 -17589 152104 -17545
rect 152148 -17589 152204 -17545
rect 152248 -17589 152304 -17545
rect 152348 -17589 152404 -17545
rect 152448 -17589 173611 -17545
rect 109734 -17645 173611 -17589
rect 109734 -17689 144904 -17645
rect 144948 -17689 145004 -17645
rect 145048 -17689 145104 -17645
rect 145148 -17689 145204 -17645
rect 145248 -17689 145304 -17645
rect 145348 -17689 145404 -17645
rect 145448 -17689 145504 -17645
rect 145548 -17689 145604 -17645
rect 145648 -17689 145704 -17645
rect 145748 -17689 145804 -17645
rect 145848 -17689 145904 -17645
rect 145948 -17689 146004 -17645
rect 146048 -17689 146104 -17645
rect 146148 -17689 146204 -17645
rect 146248 -17689 146304 -17645
rect 146348 -17689 146404 -17645
rect 146448 -17689 146904 -17645
rect 146948 -17689 147004 -17645
rect 147048 -17689 147104 -17645
rect 147148 -17689 147204 -17645
rect 147248 -17689 147304 -17645
rect 147348 -17689 147404 -17645
rect 147448 -17689 147504 -17645
rect 147548 -17689 147604 -17645
rect 147648 -17689 147704 -17645
rect 147748 -17689 147804 -17645
rect 147848 -17689 147904 -17645
rect 147948 -17689 148004 -17645
rect 148048 -17689 148104 -17645
rect 148148 -17689 148204 -17645
rect 148248 -17689 148304 -17645
rect 148348 -17689 148404 -17645
rect 148448 -17689 148904 -17645
rect 148948 -17689 149004 -17645
rect 149048 -17689 149104 -17645
rect 149148 -17689 149204 -17645
rect 149248 -17689 149304 -17645
rect 149348 -17689 149404 -17645
rect 149448 -17689 149504 -17645
rect 149548 -17689 149604 -17645
rect 149648 -17689 149704 -17645
rect 149748 -17689 149804 -17645
rect 149848 -17689 149904 -17645
rect 149948 -17689 150004 -17645
rect 150048 -17689 150104 -17645
rect 150148 -17689 150204 -17645
rect 150248 -17689 150304 -17645
rect 150348 -17689 150404 -17645
rect 150448 -17689 150904 -17645
rect 150948 -17689 151004 -17645
rect 151048 -17689 151104 -17645
rect 151148 -17689 151204 -17645
rect 151248 -17689 151304 -17645
rect 151348 -17689 151404 -17645
rect 151448 -17689 151504 -17645
rect 151548 -17689 151604 -17645
rect 151648 -17689 151704 -17645
rect 151748 -17689 151804 -17645
rect 151848 -17689 151904 -17645
rect 151948 -17689 152004 -17645
rect 152048 -17689 152104 -17645
rect 152148 -17689 152204 -17645
rect 152248 -17689 152304 -17645
rect 152348 -17689 152404 -17645
rect 152448 -17689 173611 -17645
rect 109734 -17745 173611 -17689
rect 109734 -17789 144904 -17745
rect 144948 -17789 145004 -17745
rect 145048 -17789 145104 -17745
rect 145148 -17789 145204 -17745
rect 145248 -17789 145304 -17745
rect 145348 -17789 145404 -17745
rect 145448 -17789 145504 -17745
rect 145548 -17789 145604 -17745
rect 145648 -17789 145704 -17745
rect 145748 -17789 145804 -17745
rect 145848 -17789 145904 -17745
rect 145948 -17789 146004 -17745
rect 146048 -17789 146104 -17745
rect 146148 -17789 146204 -17745
rect 146248 -17789 146304 -17745
rect 146348 -17789 146404 -17745
rect 146448 -17789 146904 -17745
rect 146948 -17789 147004 -17745
rect 147048 -17789 147104 -17745
rect 147148 -17789 147204 -17745
rect 147248 -17789 147304 -17745
rect 147348 -17789 147404 -17745
rect 147448 -17789 147504 -17745
rect 147548 -17789 147604 -17745
rect 147648 -17789 147704 -17745
rect 147748 -17789 147804 -17745
rect 147848 -17789 147904 -17745
rect 147948 -17789 148004 -17745
rect 148048 -17789 148104 -17745
rect 148148 -17789 148204 -17745
rect 148248 -17789 148304 -17745
rect 148348 -17789 148404 -17745
rect 148448 -17789 148904 -17745
rect 148948 -17789 149004 -17745
rect 149048 -17789 149104 -17745
rect 149148 -17789 149204 -17745
rect 149248 -17789 149304 -17745
rect 149348 -17789 149404 -17745
rect 149448 -17789 149504 -17745
rect 149548 -17789 149604 -17745
rect 149648 -17789 149704 -17745
rect 149748 -17789 149804 -17745
rect 149848 -17789 149904 -17745
rect 149948 -17789 150004 -17745
rect 150048 -17789 150104 -17745
rect 150148 -17789 150204 -17745
rect 150248 -17789 150304 -17745
rect 150348 -17789 150404 -17745
rect 150448 -17789 150904 -17745
rect 150948 -17789 151004 -17745
rect 151048 -17789 151104 -17745
rect 151148 -17789 151204 -17745
rect 151248 -17789 151304 -17745
rect 151348 -17789 151404 -17745
rect 151448 -17789 151504 -17745
rect 151548 -17789 151604 -17745
rect 151648 -17789 151704 -17745
rect 151748 -17789 151804 -17745
rect 151848 -17789 151904 -17745
rect 151948 -17789 152004 -17745
rect 152048 -17789 152104 -17745
rect 152148 -17789 152204 -17745
rect 152248 -17789 152304 -17745
rect 152348 -17789 152404 -17745
rect 152448 -17789 173611 -17745
rect 109734 -17830 173611 -17789
rect 174124 -17830 178142 -17214
rect 109734 -17845 178142 -17830
rect 109734 -17889 144904 -17845
rect 144948 -17889 145004 -17845
rect 145048 -17889 145104 -17845
rect 145148 -17889 145204 -17845
rect 145248 -17889 145304 -17845
rect 145348 -17889 145404 -17845
rect 145448 -17889 145504 -17845
rect 145548 -17889 145604 -17845
rect 145648 -17889 145704 -17845
rect 145748 -17889 145804 -17845
rect 145848 -17889 145904 -17845
rect 145948 -17889 146004 -17845
rect 146048 -17889 146104 -17845
rect 146148 -17889 146204 -17845
rect 146248 -17889 146304 -17845
rect 146348 -17889 146404 -17845
rect 146448 -17889 146904 -17845
rect 146948 -17889 147004 -17845
rect 147048 -17889 147104 -17845
rect 147148 -17889 147204 -17845
rect 147248 -17889 147304 -17845
rect 147348 -17889 147404 -17845
rect 147448 -17889 147504 -17845
rect 147548 -17889 147604 -17845
rect 147648 -17889 147704 -17845
rect 147748 -17889 147804 -17845
rect 147848 -17889 147904 -17845
rect 147948 -17889 148004 -17845
rect 148048 -17889 148104 -17845
rect 148148 -17889 148204 -17845
rect 148248 -17889 148304 -17845
rect 148348 -17889 148404 -17845
rect 148448 -17889 148904 -17845
rect 148948 -17889 149004 -17845
rect 149048 -17889 149104 -17845
rect 149148 -17889 149204 -17845
rect 149248 -17889 149304 -17845
rect 149348 -17889 149404 -17845
rect 149448 -17889 149504 -17845
rect 149548 -17889 149604 -17845
rect 149648 -17889 149704 -17845
rect 149748 -17889 149804 -17845
rect 149848 -17889 149904 -17845
rect 149948 -17889 150004 -17845
rect 150048 -17889 150104 -17845
rect 150148 -17889 150204 -17845
rect 150248 -17889 150304 -17845
rect 150348 -17889 150404 -17845
rect 150448 -17889 150904 -17845
rect 150948 -17889 151004 -17845
rect 151048 -17889 151104 -17845
rect 151148 -17889 151204 -17845
rect 151248 -17889 151304 -17845
rect 151348 -17889 151404 -17845
rect 151448 -17889 151504 -17845
rect 151548 -17889 151604 -17845
rect 151648 -17889 151704 -17845
rect 151748 -17889 151804 -17845
rect 151848 -17889 151904 -17845
rect 151948 -17889 152004 -17845
rect 152048 -17889 152104 -17845
rect 152148 -17889 152204 -17845
rect 152248 -17889 152304 -17845
rect 152348 -17889 152404 -17845
rect 152448 -17889 178142 -17845
rect 109734 -17945 178142 -17889
rect 109734 -17989 144904 -17945
rect 144948 -17989 145004 -17945
rect 145048 -17989 145104 -17945
rect 145148 -17989 145204 -17945
rect 145248 -17989 145304 -17945
rect 145348 -17989 145404 -17945
rect 145448 -17989 145504 -17945
rect 145548 -17989 145604 -17945
rect 145648 -17989 145704 -17945
rect 145748 -17989 145804 -17945
rect 145848 -17989 145904 -17945
rect 145948 -17989 146004 -17945
rect 146048 -17989 146104 -17945
rect 146148 -17989 146204 -17945
rect 146248 -17989 146304 -17945
rect 146348 -17989 146404 -17945
rect 146448 -17989 146904 -17945
rect 146948 -17989 147004 -17945
rect 147048 -17989 147104 -17945
rect 147148 -17989 147204 -17945
rect 147248 -17989 147304 -17945
rect 147348 -17989 147404 -17945
rect 147448 -17989 147504 -17945
rect 147548 -17989 147604 -17945
rect 147648 -17989 147704 -17945
rect 147748 -17989 147804 -17945
rect 147848 -17989 147904 -17945
rect 147948 -17989 148004 -17945
rect 148048 -17989 148104 -17945
rect 148148 -17989 148204 -17945
rect 148248 -17989 148304 -17945
rect 148348 -17989 148404 -17945
rect 148448 -17989 148904 -17945
rect 148948 -17989 149004 -17945
rect 149048 -17989 149104 -17945
rect 149148 -17989 149204 -17945
rect 149248 -17989 149304 -17945
rect 149348 -17989 149404 -17945
rect 149448 -17989 149504 -17945
rect 149548 -17989 149604 -17945
rect 149648 -17989 149704 -17945
rect 149748 -17989 149804 -17945
rect 149848 -17989 149904 -17945
rect 149948 -17989 150004 -17945
rect 150048 -17989 150104 -17945
rect 150148 -17989 150204 -17945
rect 150248 -17989 150304 -17945
rect 150348 -17989 150404 -17945
rect 150448 -17989 150904 -17945
rect 150948 -17989 151004 -17945
rect 151048 -17989 151104 -17945
rect 151148 -17989 151204 -17945
rect 151248 -17989 151304 -17945
rect 151348 -17989 151404 -17945
rect 151448 -17989 151504 -17945
rect 151548 -17989 151604 -17945
rect 151648 -17989 151704 -17945
rect 151748 -17989 151804 -17945
rect 151848 -17989 151904 -17945
rect 151948 -17989 152004 -17945
rect 152048 -17989 152104 -17945
rect 152148 -17989 152204 -17945
rect 152248 -17989 152304 -17945
rect 152348 -17989 152404 -17945
rect 152448 -17989 178142 -17945
rect 109734 -18045 178142 -17989
rect 109734 -18089 144904 -18045
rect 144948 -18089 145004 -18045
rect 145048 -18089 145104 -18045
rect 145148 -18089 145204 -18045
rect 145248 -18089 145304 -18045
rect 145348 -18089 145404 -18045
rect 145448 -18089 145504 -18045
rect 145548 -18089 145604 -18045
rect 145648 -18089 145704 -18045
rect 145748 -18089 145804 -18045
rect 145848 -18089 145904 -18045
rect 145948 -18089 146004 -18045
rect 146048 -18089 146104 -18045
rect 146148 -18089 146204 -18045
rect 146248 -18089 146304 -18045
rect 146348 -18089 146404 -18045
rect 146448 -18089 146904 -18045
rect 146948 -18089 147004 -18045
rect 147048 -18089 147104 -18045
rect 147148 -18089 147204 -18045
rect 147248 -18089 147304 -18045
rect 147348 -18089 147404 -18045
rect 147448 -18089 147504 -18045
rect 147548 -18089 147604 -18045
rect 147648 -18089 147704 -18045
rect 147748 -18089 147804 -18045
rect 147848 -18089 147904 -18045
rect 147948 -18089 148004 -18045
rect 148048 -18089 148104 -18045
rect 148148 -18089 148204 -18045
rect 148248 -18089 148304 -18045
rect 148348 -18089 148404 -18045
rect 148448 -18089 148904 -18045
rect 148948 -18089 149004 -18045
rect 149048 -18089 149104 -18045
rect 149148 -18089 149204 -18045
rect 149248 -18089 149304 -18045
rect 149348 -18089 149404 -18045
rect 149448 -18089 149504 -18045
rect 149548 -18089 149604 -18045
rect 149648 -18089 149704 -18045
rect 149748 -18089 149804 -18045
rect 149848 -18089 149904 -18045
rect 149948 -18089 150004 -18045
rect 150048 -18089 150104 -18045
rect 150148 -18089 150204 -18045
rect 150248 -18089 150304 -18045
rect 150348 -18089 150404 -18045
rect 150448 -18089 150904 -18045
rect 150948 -18089 151004 -18045
rect 151048 -18089 151104 -18045
rect 151148 -18089 151204 -18045
rect 151248 -18089 151304 -18045
rect 151348 -18089 151404 -18045
rect 151448 -18089 151504 -18045
rect 151548 -18089 151604 -18045
rect 151648 -18089 151704 -18045
rect 151748 -18089 151804 -18045
rect 151848 -18089 151904 -18045
rect 151948 -18089 152004 -18045
rect 152048 -18089 152104 -18045
rect 152148 -18089 152204 -18045
rect 152248 -18089 152304 -18045
rect 152348 -18089 152404 -18045
rect 152448 -18089 178142 -18045
rect 109734 -18145 178142 -18089
rect 109734 -18189 144904 -18145
rect 144948 -18189 145004 -18145
rect 145048 -18189 145104 -18145
rect 145148 -18189 145204 -18145
rect 145248 -18189 145304 -18145
rect 145348 -18189 145404 -18145
rect 145448 -18189 145504 -18145
rect 145548 -18189 145604 -18145
rect 145648 -18189 145704 -18145
rect 145748 -18189 145804 -18145
rect 145848 -18189 145904 -18145
rect 145948 -18189 146004 -18145
rect 146048 -18189 146104 -18145
rect 146148 -18189 146204 -18145
rect 146248 -18189 146304 -18145
rect 146348 -18189 146404 -18145
rect 146448 -18189 146904 -18145
rect 146948 -18189 147004 -18145
rect 147048 -18189 147104 -18145
rect 147148 -18189 147204 -18145
rect 147248 -18189 147304 -18145
rect 147348 -18189 147404 -18145
rect 147448 -18189 147504 -18145
rect 147548 -18189 147604 -18145
rect 147648 -18189 147704 -18145
rect 147748 -18189 147804 -18145
rect 147848 -18189 147904 -18145
rect 147948 -18189 148004 -18145
rect 148048 -18189 148104 -18145
rect 148148 -18189 148204 -18145
rect 148248 -18189 148304 -18145
rect 148348 -18189 148404 -18145
rect 148448 -18189 148904 -18145
rect 148948 -18189 149004 -18145
rect 149048 -18189 149104 -18145
rect 149148 -18189 149204 -18145
rect 149248 -18189 149304 -18145
rect 149348 -18189 149404 -18145
rect 149448 -18189 149504 -18145
rect 149548 -18189 149604 -18145
rect 149648 -18189 149704 -18145
rect 149748 -18189 149804 -18145
rect 149848 -18189 149904 -18145
rect 149948 -18189 150004 -18145
rect 150048 -18189 150104 -18145
rect 150148 -18189 150204 -18145
rect 150248 -18189 150304 -18145
rect 150348 -18189 150404 -18145
rect 150448 -18189 150904 -18145
rect 150948 -18189 151004 -18145
rect 151048 -18189 151104 -18145
rect 151148 -18189 151204 -18145
rect 151248 -18189 151304 -18145
rect 151348 -18189 151404 -18145
rect 151448 -18189 151504 -18145
rect 151548 -18189 151604 -18145
rect 151648 -18189 151704 -18145
rect 151748 -18189 151804 -18145
rect 151848 -18189 151904 -18145
rect 151948 -18189 152004 -18145
rect 152048 -18189 152104 -18145
rect 152148 -18189 152204 -18145
rect 152248 -18189 152304 -18145
rect 152348 -18189 152404 -18145
rect 152448 -18189 178142 -18145
rect 109734 -18245 178142 -18189
rect 109734 -18289 144904 -18245
rect 144948 -18289 145004 -18245
rect 145048 -18289 145104 -18245
rect 145148 -18289 145204 -18245
rect 145248 -18289 145304 -18245
rect 145348 -18289 145404 -18245
rect 145448 -18289 145504 -18245
rect 145548 -18289 145604 -18245
rect 145648 -18289 145704 -18245
rect 145748 -18289 145804 -18245
rect 145848 -18289 145904 -18245
rect 145948 -18289 146004 -18245
rect 146048 -18289 146104 -18245
rect 146148 -18289 146204 -18245
rect 146248 -18289 146304 -18245
rect 146348 -18289 146404 -18245
rect 146448 -18289 146904 -18245
rect 146948 -18289 147004 -18245
rect 147048 -18289 147104 -18245
rect 147148 -18289 147204 -18245
rect 147248 -18289 147304 -18245
rect 147348 -18289 147404 -18245
rect 147448 -18289 147504 -18245
rect 147548 -18289 147604 -18245
rect 147648 -18289 147704 -18245
rect 147748 -18289 147804 -18245
rect 147848 -18289 147904 -18245
rect 147948 -18289 148004 -18245
rect 148048 -18289 148104 -18245
rect 148148 -18289 148204 -18245
rect 148248 -18289 148304 -18245
rect 148348 -18289 148404 -18245
rect 148448 -18289 148904 -18245
rect 148948 -18289 149004 -18245
rect 149048 -18289 149104 -18245
rect 149148 -18289 149204 -18245
rect 149248 -18289 149304 -18245
rect 149348 -18289 149404 -18245
rect 149448 -18289 149504 -18245
rect 149548 -18289 149604 -18245
rect 149648 -18289 149704 -18245
rect 149748 -18289 149804 -18245
rect 149848 -18289 149904 -18245
rect 149948 -18289 150004 -18245
rect 150048 -18289 150104 -18245
rect 150148 -18289 150204 -18245
rect 150248 -18289 150304 -18245
rect 150348 -18289 150404 -18245
rect 150448 -18289 150904 -18245
rect 150948 -18289 151004 -18245
rect 151048 -18289 151104 -18245
rect 151148 -18289 151204 -18245
rect 151248 -18289 151304 -18245
rect 151348 -18289 151404 -18245
rect 151448 -18289 151504 -18245
rect 151548 -18289 151604 -18245
rect 151648 -18289 151704 -18245
rect 151748 -18289 151804 -18245
rect 151848 -18289 151904 -18245
rect 151948 -18289 152004 -18245
rect 152048 -18289 152104 -18245
rect 152148 -18289 152204 -18245
rect 152248 -18289 152304 -18245
rect 152348 -18289 152404 -18245
rect 152448 -18289 178142 -18245
rect 109734 -18345 178142 -18289
rect 109734 -18389 144904 -18345
rect 144948 -18389 145004 -18345
rect 145048 -18389 145104 -18345
rect 145148 -18389 145204 -18345
rect 145248 -18389 145304 -18345
rect 145348 -18389 145404 -18345
rect 145448 -18389 145504 -18345
rect 145548 -18389 145604 -18345
rect 145648 -18389 145704 -18345
rect 145748 -18389 145804 -18345
rect 145848 -18389 145904 -18345
rect 145948 -18389 146004 -18345
rect 146048 -18389 146104 -18345
rect 146148 -18389 146204 -18345
rect 146248 -18389 146304 -18345
rect 146348 -18389 146404 -18345
rect 146448 -18389 146904 -18345
rect 146948 -18389 147004 -18345
rect 147048 -18389 147104 -18345
rect 147148 -18389 147204 -18345
rect 147248 -18389 147304 -18345
rect 147348 -18389 147404 -18345
rect 147448 -18389 147504 -18345
rect 147548 -18389 147604 -18345
rect 147648 -18389 147704 -18345
rect 147748 -18389 147804 -18345
rect 147848 -18389 147904 -18345
rect 147948 -18389 148004 -18345
rect 148048 -18389 148104 -18345
rect 148148 -18389 148204 -18345
rect 148248 -18389 148304 -18345
rect 148348 -18389 148404 -18345
rect 148448 -18389 148904 -18345
rect 148948 -18389 149004 -18345
rect 149048 -18389 149104 -18345
rect 149148 -18389 149204 -18345
rect 149248 -18389 149304 -18345
rect 149348 -18389 149404 -18345
rect 149448 -18389 149504 -18345
rect 149548 -18389 149604 -18345
rect 149648 -18389 149704 -18345
rect 149748 -18389 149804 -18345
rect 149848 -18389 149904 -18345
rect 149948 -18389 150004 -18345
rect 150048 -18389 150104 -18345
rect 150148 -18389 150204 -18345
rect 150248 -18389 150304 -18345
rect 150348 -18389 150404 -18345
rect 150448 -18389 150904 -18345
rect 150948 -18389 151004 -18345
rect 151048 -18389 151104 -18345
rect 151148 -18389 151204 -18345
rect 151248 -18389 151304 -18345
rect 151348 -18389 151404 -18345
rect 151448 -18389 151504 -18345
rect 151548 -18389 151604 -18345
rect 151648 -18389 151704 -18345
rect 151748 -18389 151804 -18345
rect 151848 -18389 151904 -18345
rect 151948 -18389 152004 -18345
rect 152048 -18389 152104 -18345
rect 152148 -18389 152204 -18345
rect 152248 -18389 152304 -18345
rect 152348 -18389 152404 -18345
rect 152448 -18389 178142 -18345
rect 109734 -18445 178142 -18389
rect 109734 -18489 144904 -18445
rect 144948 -18489 145004 -18445
rect 145048 -18489 145104 -18445
rect 145148 -18489 145204 -18445
rect 145248 -18489 145304 -18445
rect 145348 -18489 145404 -18445
rect 145448 -18489 145504 -18445
rect 145548 -18489 145604 -18445
rect 145648 -18489 145704 -18445
rect 145748 -18489 145804 -18445
rect 145848 -18489 145904 -18445
rect 145948 -18489 146004 -18445
rect 146048 -18489 146104 -18445
rect 146148 -18489 146204 -18445
rect 146248 -18489 146304 -18445
rect 146348 -18489 146404 -18445
rect 146448 -18489 146904 -18445
rect 146948 -18489 147004 -18445
rect 147048 -18489 147104 -18445
rect 147148 -18489 147204 -18445
rect 147248 -18489 147304 -18445
rect 147348 -18489 147404 -18445
rect 147448 -18489 147504 -18445
rect 147548 -18489 147604 -18445
rect 147648 -18489 147704 -18445
rect 147748 -18489 147804 -18445
rect 147848 -18489 147904 -18445
rect 147948 -18489 148004 -18445
rect 148048 -18489 148104 -18445
rect 148148 -18489 148204 -18445
rect 148248 -18489 148304 -18445
rect 148348 -18489 148404 -18445
rect 148448 -18489 148904 -18445
rect 148948 -18489 149004 -18445
rect 149048 -18489 149104 -18445
rect 149148 -18489 149204 -18445
rect 149248 -18489 149304 -18445
rect 149348 -18489 149404 -18445
rect 149448 -18489 149504 -18445
rect 149548 -18489 149604 -18445
rect 149648 -18489 149704 -18445
rect 149748 -18489 149804 -18445
rect 149848 -18489 149904 -18445
rect 149948 -18489 150004 -18445
rect 150048 -18489 150104 -18445
rect 150148 -18489 150204 -18445
rect 150248 -18489 150304 -18445
rect 150348 -18489 150404 -18445
rect 150448 -18489 150904 -18445
rect 150948 -18489 151004 -18445
rect 151048 -18489 151104 -18445
rect 151148 -18489 151204 -18445
rect 151248 -18489 151304 -18445
rect 151348 -18489 151404 -18445
rect 151448 -18489 151504 -18445
rect 151548 -18489 151604 -18445
rect 151648 -18489 151704 -18445
rect 151748 -18489 151804 -18445
rect 151848 -18489 151904 -18445
rect 151948 -18489 152004 -18445
rect 152048 -18489 152104 -18445
rect 152148 -18489 152204 -18445
rect 152248 -18489 152304 -18445
rect 152348 -18489 152404 -18445
rect 152448 -18489 178142 -18445
rect 109734 -18545 178142 -18489
rect 109734 -18589 144904 -18545
rect 144948 -18589 145004 -18545
rect 145048 -18589 145104 -18545
rect 145148 -18589 145204 -18545
rect 145248 -18589 145304 -18545
rect 145348 -18589 145404 -18545
rect 145448 -18589 145504 -18545
rect 145548 -18589 145604 -18545
rect 145648 -18589 145704 -18545
rect 145748 -18589 145804 -18545
rect 145848 -18589 145904 -18545
rect 145948 -18589 146004 -18545
rect 146048 -18589 146104 -18545
rect 146148 -18589 146204 -18545
rect 146248 -18589 146304 -18545
rect 146348 -18589 146404 -18545
rect 146448 -18589 146904 -18545
rect 146948 -18589 147004 -18545
rect 147048 -18589 147104 -18545
rect 147148 -18589 147204 -18545
rect 147248 -18589 147304 -18545
rect 147348 -18589 147404 -18545
rect 147448 -18589 147504 -18545
rect 147548 -18589 147604 -18545
rect 147648 -18589 147704 -18545
rect 147748 -18589 147804 -18545
rect 147848 -18589 147904 -18545
rect 147948 -18589 148004 -18545
rect 148048 -18589 148104 -18545
rect 148148 -18589 148204 -18545
rect 148248 -18589 148304 -18545
rect 148348 -18589 148404 -18545
rect 148448 -18589 148904 -18545
rect 148948 -18589 149004 -18545
rect 149048 -18589 149104 -18545
rect 149148 -18589 149204 -18545
rect 149248 -18589 149304 -18545
rect 149348 -18589 149404 -18545
rect 149448 -18589 149504 -18545
rect 149548 -18589 149604 -18545
rect 149648 -18589 149704 -18545
rect 149748 -18589 149804 -18545
rect 149848 -18589 149904 -18545
rect 149948 -18589 150004 -18545
rect 150048 -18589 150104 -18545
rect 150148 -18589 150204 -18545
rect 150248 -18589 150304 -18545
rect 150348 -18589 150404 -18545
rect 150448 -18589 150904 -18545
rect 150948 -18589 151004 -18545
rect 151048 -18589 151104 -18545
rect 151148 -18589 151204 -18545
rect 151248 -18589 151304 -18545
rect 151348 -18589 151404 -18545
rect 151448 -18589 151504 -18545
rect 151548 -18589 151604 -18545
rect 151648 -18589 151704 -18545
rect 151748 -18589 151804 -18545
rect 151848 -18589 151904 -18545
rect 151948 -18589 152004 -18545
rect 152048 -18589 152104 -18545
rect 152148 -18589 152204 -18545
rect 152248 -18589 152304 -18545
rect 152348 -18589 152404 -18545
rect 152448 -18589 178142 -18545
rect 109734 -18645 178142 -18589
rect 109734 -18689 144904 -18645
rect 144948 -18689 145004 -18645
rect 145048 -18689 145104 -18645
rect 145148 -18689 145204 -18645
rect 145248 -18689 145304 -18645
rect 145348 -18689 145404 -18645
rect 145448 -18689 145504 -18645
rect 145548 -18689 145604 -18645
rect 145648 -18689 145704 -18645
rect 145748 -18689 145804 -18645
rect 145848 -18689 145904 -18645
rect 145948 -18689 146004 -18645
rect 146048 -18689 146104 -18645
rect 146148 -18689 146204 -18645
rect 146248 -18689 146304 -18645
rect 146348 -18689 146404 -18645
rect 146448 -18689 146904 -18645
rect 146948 -18689 147004 -18645
rect 147048 -18689 147104 -18645
rect 147148 -18689 147204 -18645
rect 147248 -18689 147304 -18645
rect 147348 -18689 147404 -18645
rect 147448 -18689 147504 -18645
rect 147548 -18689 147604 -18645
rect 147648 -18689 147704 -18645
rect 147748 -18689 147804 -18645
rect 147848 -18689 147904 -18645
rect 147948 -18689 148004 -18645
rect 148048 -18689 148104 -18645
rect 148148 -18689 148204 -18645
rect 148248 -18689 148304 -18645
rect 148348 -18689 148404 -18645
rect 148448 -18689 148904 -18645
rect 148948 -18689 149004 -18645
rect 149048 -18689 149104 -18645
rect 149148 -18689 149204 -18645
rect 149248 -18689 149304 -18645
rect 149348 -18689 149404 -18645
rect 149448 -18689 149504 -18645
rect 149548 -18689 149604 -18645
rect 149648 -18689 149704 -18645
rect 149748 -18689 149804 -18645
rect 149848 -18689 149904 -18645
rect 149948 -18689 150004 -18645
rect 150048 -18689 150104 -18645
rect 150148 -18689 150204 -18645
rect 150248 -18689 150304 -18645
rect 150348 -18689 150404 -18645
rect 150448 -18689 150904 -18645
rect 150948 -18689 151004 -18645
rect 151048 -18689 151104 -18645
rect 151148 -18689 151204 -18645
rect 151248 -18689 151304 -18645
rect 151348 -18689 151404 -18645
rect 151448 -18689 151504 -18645
rect 151548 -18689 151604 -18645
rect 151648 -18689 151704 -18645
rect 151748 -18689 151804 -18645
rect 151848 -18689 151904 -18645
rect 151948 -18689 152004 -18645
rect 152048 -18689 152104 -18645
rect 152148 -18689 152204 -18645
rect 152248 -18689 152304 -18645
rect 152348 -18689 152404 -18645
rect 152448 -18689 178142 -18645
rect 109734 -18745 178142 -18689
rect 109734 -18789 144904 -18745
rect 144948 -18789 145004 -18745
rect 145048 -18789 145104 -18745
rect 145148 -18789 145204 -18745
rect 145248 -18789 145304 -18745
rect 145348 -18789 145404 -18745
rect 145448 -18789 145504 -18745
rect 145548 -18789 145604 -18745
rect 145648 -18789 145704 -18745
rect 145748 -18789 145804 -18745
rect 145848 -18789 145904 -18745
rect 145948 -18789 146004 -18745
rect 146048 -18789 146104 -18745
rect 146148 -18789 146204 -18745
rect 146248 -18789 146304 -18745
rect 146348 -18789 146404 -18745
rect 146448 -18789 146904 -18745
rect 146948 -18789 147004 -18745
rect 147048 -18789 147104 -18745
rect 147148 -18789 147204 -18745
rect 147248 -18789 147304 -18745
rect 147348 -18789 147404 -18745
rect 147448 -18789 147504 -18745
rect 147548 -18789 147604 -18745
rect 147648 -18789 147704 -18745
rect 147748 -18789 147804 -18745
rect 147848 -18789 147904 -18745
rect 147948 -18789 148004 -18745
rect 148048 -18789 148104 -18745
rect 148148 -18789 148204 -18745
rect 148248 -18789 148304 -18745
rect 148348 -18789 148404 -18745
rect 148448 -18789 148904 -18745
rect 148948 -18789 149004 -18745
rect 149048 -18789 149104 -18745
rect 149148 -18789 149204 -18745
rect 149248 -18789 149304 -18745
rect 149348 -18789 149404 -18745
rect 149448 -18789 149504 -18745
rect 149548 -18789 149604 -18745
rect 149648 -18789 149704 -18745
rect 149748 -18789 149804 -18745
rect 149848 -18789 149904 -18745
rect 149948 -18789 150004 -18745
rect 150048 -18789 150104 -18745
rect 150148 -18789 150204 -18745
rect 150248 -18789 150304 -18745
rect 150348 -18789 150404 -18745
rect 150448 -18789 150904 -18745
rect 150948 -18789 151004 -18745
rect 151048 -18789 151104 -18745
rect 151148 -18789 151204 -18745
rect 151248 -18789 151304 -18745
rect 151348 -18789 151404 -18745
rect 151448 -18789 151504 -18745
rect 151548 -18789 151604 -18745
rect 151648 -18789 151704 -18745
rect 151748 -18789 151804 -18745
rect 151848 -18789 151904 -18745
rect 151948 -18789 152004 -18745
rect 152048 -18789 152104 -18745
rect 152148 -18789 152204 -18745
rect 152248 -18789 152304 -18745
rect 152348 -18789 152404 -18745
rect 152448 -18789 178142 -18745
rect 109734 -18845 178142 -18789
rect 109734 -18889 144904 -18845
rect 144948 -18889 145004 -18845
rect 145048 -18889 145104 -18845
rect 145148 -18889 145204 -18845
rect 145248 -18889 145304 -18845
rect 145348 -18889 145404 -18845
rect 145448 -18889 145504 -18845
rect 145548 -18889 145604 -18845
rect 145648 -18889 145704 -18845
rect 145748 -18889 145804 -18845
rect 145848 -18889 145904 -18845
rect 145948 -18889 146004 -18845
rect 146048 -18889 146104 -18845
rect 146148 -18889 146204 -18845
rect 146248 -18889 146304 -18845
rect 146348 -18889 146404 -18845
rect 146448 -18889 146904 -18845
rect 146948 -18889 147004 -18845
rect 147048 -18889 147104 -18845
rect 147148 -18889 147204 -18845
rect 147248 -18889 147304 -18845
rect 147348 -18889 147404 -18845
rect 147448 -18889 147504 -18845
rect 147548 -18889 147604 -18845
rect 147648 -18889 147704 -18845
rect 147748 -18889 147804 -18845
rect 147848 -18889 147904 -18845
rect 147948 -18889 148004 -18845
rect 148048 -18889 148104 -18845
rect 148148 -18889 148204 -18845
rect 148248 -18889 148304 -18845
rect 148348 -18889 148404 -18845
rect 148448 -18889 148904 -18845
rect 148948 -18889 149004 -18845
rect 149048 -18889 149104 -18845
rect 149148 -18889 149204 -18845
rect 149248 -18889 149304 -18845
rect 149348 -18889 149404 -18845
rect 149448 -18889 149504 -18845
rect 149548 -18889 149604 -18845
rect 149648 -18889 149704 -18845
rect 149748 -18889 149804 -18845
rect 149848 -18889 149904 -18845
rect 149948 -18889 150004 -18845
rect 150048 -18889 150104 -18845
rect 150148 -18889 150204 -18845
rect 150248 -18889 150304 -18845
rect 150348 -18889 150404 -18845
rect 150448 -18889 150904 -18845
rect 150948 -18889 151004 -18845
rect 151048 -18889 151104 -18845
rect 151148 -18889 151204 -18845
rect 151248 -18889 151304 -18845
rect 151348 -18889 151404 -18845
rect 151448 -18889 151504 -18845
rect 151548 -18889 151604 -18845
rect 151648 -18889 151704 -18845
rect 151748 -18889 151804 -18845
rect 151848 -18889 151904 -18845
rect 151948 -18889 152004 -18845
rect 152048 -18889 152104 -18845
rect 152148 -18889 152204 -18845
rect 152248 -18889 152304 -18845
rect 152348 -18889 152404 -18845
rect 152448 -18889 178142 -18845
rect 109734 -18945 178142 -18889
rect 109734 -18989 144904 -18945
rect 144948 -18989 145004 -18945
rect 145048 -18989 145104 -18945
rect 145148 -18989 145204 -18945
rect 145248 -18989 145304 -18945
rect 145348 -18989 145404 -18945
rect 145448 -18989 145504 -18945
rect 145548 -18989 145604 -18945
rect 145648 -18989 145704 -18945
rect 145748 -18989 145804 -18945
rect 145848 -18989 145904 -18945
rect 145948 -18989 146004 -18945
rect 146048 -18989 146104 -18945
rect 146148 -18989 146204 -18945
rect 146248 -18989 146304 -18945
rect 146348 -18989 146404 -18945
rect 146448 -18989 146904 -18945
rect 146948 -18989 147004 -18945
rect 147048 -18989 147104 -18945
rect 147148 -18989 147204 -18945
rect 147248 -18989 147304 -18945
rect 147348 -18989 147404 -18945
rect 147448 -18989 147504 -18945
rect 147548 -18989 147604 -18945
rect 147648 -18989 147704 -18945
rect 147748 -18989 147804 -18945
rect 147848 -18989 147904 -18945
rect 147948 -18989 148004 -18945
rect 148048 -18989 148104 -18945
rect 148148 -18989 148204 -18945
rect 148248 -18989 148304 -18945
rect 148348 -18989 148404 -18945
rect 148448 -18989 148904 -18945
rect 148948 -18989 149004 -18945
rect 149048 -18989 149104 -18945
rect 149148 -18989 149204 -18945
rect 149248 -18989 149304 -18945
rect 149348 -18989 149404 -18945
rect 149448 -18989 149504 -18945
rect 149548 -18989 149604 -18945
rect 149648 -18989 149704 -18945
rect 149748 -18989 149804 -18945
rect 149848 -18989 149904 -18945
rect 149948 -18989 150004 -18945
rect 150048 -18989 150104 -18945
rect 150148 -18989 150204 -18945
rect 150248 -18989 150304 -18945
rect 150348 -18989 150404 -18945
rect 150448 -18989 150904 -18945
rect 150948 -18989 151004 -18945
rect 151048 -18989 151104 -18945
rect 151148 -18989 151204 -18945
rect 151248 -18989 151304 -18945
rect 151348 -18989 151404 -18945
rect 151448 -18989 151504 -18945
rect 151548 -18989 151604 -18945
rect 151648 -18989 151704 -18945
rect 151748 -18989 151804 -18945
rect 151848 -18989 151904 -18945
rect 151948 -18989 152004 -18945
rect 152048 -18989 152104 -18945
rect 152148 -18989 152204 -18945
rect 152248 -18989 152304 -18945
rect 152348 -18989 152404 -18945
rect 152448 -18989 178142 -18945
rect 58258 -20180 58334 -19695
rect 58746 -20180 58822 -19695
rect 59234 -20180 59310 -19695
rect 59722 -20180 59798 -19695
rect 60210 -20180 60286 -19695
rect 60698 -20180 60774 -19695
rect 61186 -20180 61262 -19695
rect 61674 -20180 61750 -19695
rect 62162 -20180 62238 -19695
rect 62650 -20180 62726 -19695
rect 63138 -20180 63214 -19695
rect 63626 -20180 63702 -19695
rect 64114 -20180 64190 -19695
rect 64602 -20180 64678 -19695
rect 65090 -20180 65166 -19695
rect 65578 -20180 65654 -19695
rect 66066 -20180 66142 -19695
rect 66554 -20180 66630 -19695
rect 67042 -20180 67118 -19695
rect 67530 -20180 67606 -19695
rect 68018 -20180 68094 -19695
rect 68506 -20180 68582 -19695
rect 68994 -20180 69070 -19695
rect 69482 -20180 69558 -19695
rect 69970 -20180 70046 -19695
rect 70458 -20180 70534 -19695
rect 70946 -20180 71022 -19695
rect 71434 -20180 71510 -19695
rect 71922 -20180 71998 -19695
rect 72410 -20180 72486 -19695
rect 72898 -20180 72974 -19695
rect 73386 -20180 73462 -19695
rect 73874 -20180 73950 -19695
rect 74362 -20180 74438 -19695
rect 74850 -20180 74926 -19695
rect 75338 -20180 75414 -19695
rect 75826 -20180 75902 -19695
rect 76314 -20180 76390 -19695
rect 76802 -20180 76878 -19695
rect 77290 -20180 77366 -19695
rect 77778 -20180 77854 -19695
rect 78266 -20180 78342 -19695
rect 78754 -20180 78830 -19695
rect 79242 -20180 79318 -19695
rect 79730 -20180 79806 -19695
rect 80218 -20180 80294 -19695
rect 80706 -20180 80782 -19695
rect 81194 -20180 81270 -19695
rect 81682 -20180 81758 -19695
rect 82170 -20180 82246 -19695
rect 85258 -20180 85334 -19695
rect 85746 -20180 85822 -19695
rect 86234 -20180 86310 -19695
rect 86722 -20180 86798 -19695
rect 87210 -20180 87286 -19695
rect 87698 -20180 87774 -19695
rect 88186 -20180 88262 -19695
rect 88674 -20180 88750 -19695
rect 89162 -20180 89238 -19695
rect 89650 -20180 89726 -19695
rect 90138 -20180 90214 -19695
rect 90626 -20180 90702 -19695
rect 91114 -20180 91190 -19695
rect 91602 -20180 91678 -19695
rect 92090 -20180 92166 -19695
rect 92578 -20180 92654 -19695
rect 93066 -20180 93142 -19695
rect 93554 -20180 93630 -19695
rect 94042 -20180 94118 -19695
rect 94530 -20180 94606 -19695
rect 95018 -20180 95094 -19695
rect 95506 -20180 95582 -19695
rect 95994 -20180 96070 -19695
rect 96482 -20180 96558 -19695
rect 96970 -20180 97046 -19695
rect 97458 -20180 97534 -19695
rect 97946 -20180 98022 -19695
rect 98434 -20180 98510 -19695
rect 98922 -20180 98998 -19695
rect 99410 -20180 99486 -19695
rect 99898 -20180 99974 -19695
rect 100386 -20180 100462 -19695
rect 100874 -20180 100950 -19695
rect 101362 -20180 101438 -19695
rect 101850 -20180 101926 -19695
rect 102338 -20180 102414 -19695
rect 102826 -20180 102902 -19695
rect 103314 -20180 103390 -19695
rect 103802 -20180 103878 -19695
rect 104290 -20180 104366 -19695
rect 104778 -20180 104854 -19695
rect 105266 -20180 105342 -19695
rect 105754 -20180 105830 -19695
rect 106242 -20180 106318 -19695
rect 106730 -20180 106806 -19695
rect 107218 -20180 107294 -19695
rect 107706 -20180 107782 -19695
rect 108194 -20180 108270 -19695
rect 108682 -20180 108758 -19695
rect 109170 -20180 109246 -19695
rect 109734 -20180 178142 -18989
rect 58258 -20875 178142 -20180
rect -109116 -24026 177360 -23015
rect -109116 -24070 80849 -24026
rect 80893 -24070 80949 -24026
rect 80993 -24070 81049 -24026
rect 81093 -24070 81149 -24026
rect 81193 -24070 81249 -24026
rect 81293 -24070 81349 -24026
rect 81393 -24070 81449 -24026
rect 81493 -24070 81549 -24026
rect 81593 -24070 81649 -24026
rect 81693 -24070 81749 -24026
rect 81793 -24070 81849 -24026
rect 81893 -24070 81949 -24026
rect 81993 -24070 82049 -24026
rect 82093 -24070 82149 -24026
rect 82193 -24070 82249 -24026
rect 82293 -24070 82349 -24026
rect 82393 -24070 82849 -24026
rect 82893 -24070 82949 -24026
rect 82993 -24070 83049 -24026
rect 83093 -24070 83149 -24026
rect 83193 -24070 83249 -24026
rect 83293 -24070 83349 -24026
rect 83393 -24070 83449 -24026
rect 83493 -24070 83549 -24026
rect 83593 -24070 83649 -24026
rect 83693 -24070 83749 -24026
rect 83793 -24070 83849 -24026
rect 83893 -24070 83949 -24026
rect 83993 -24070 84049 -24026
rect 84093 -24070 84149 -24026
rect 84193 -24070 84249 -24026
rect 84293 -24070 84349 -24026
rect 84393 -24070 84849 -24026
rect 84893 -24070 84949 -24026
rect 84993 -24070 85049 -24026
rect 85093 -24070 85149 -24026
rect 85193 -24070 85249 -24026
rect 85293 -24070 85349 -24026
rect 85393 -24070 85449 -24026
rect 85493 -24070 85549 -24026
rect 85593 -24070 85649 -24026
rect 85693 -24070 85749 -24026
rect 85793 -24070 85849 -24026
rect 85893 -24070 85949 -24026
rect 85993 -24070 86049 -24026
rect 86093 -24070 86149 -24026
rect 86193 -24070 86249 -24026
rect 86293 -24070 86349 -24026
rect 86393 -24070 86849 -24026
rect 86893 -24070 86949 -24026
rect 86993 -24070 87049 -24026
rect 87093 -24070 87149 -24026
rect 87193 -24070 87249 -24026
rect 87293 -24070 87349 -24026
rect 87393 -24070 87449 -24026
rect 87493 -24070 87549 -24026
rect 87593 -24070 87649 -24026
rect 87693 -24070 87749 -24026
rect 87793 -24070 87849 -24026
rect 87893 -24070 87949 -24026
rect 87993 -24070 88049 -24026
rect 88093 -24070 88149 -24026
rect 88193 -24070 88249 -24026
rect 88293 -24070 88349 -24026
rect 88393 -24070 177360 -24026
rect -109116 -24126 177360 -24070
rect -109116 -24170 80849 -24126
rect 80893 -24170 80949 -24126
rect 80993 -24170 81049 -24126
rect 81093 -24170 81149 -24126
rect 81193 -24170 81249 -24126
rect 81293 -24170 81349 -24126
rect 81393 -24170 81449 -24126
rect 81493 -24170 81549 -24126
rect 81593 -24170 81649 -24126
rect 81693 -24170 81749 -24126
rect 81793 -24170 81849 -24126
rect 81893 -24170 81949 -24126
rect 81993 -24170 82049 -24126
rect 82093 -24170 82149 -24126
rect 82193 -24170 82249 -24126
rect 82293 -24170 82349 -24126
rect 82393 -24170 82849 -24126
rect 82893 -24170 82949 -24126
rect 82993 -24170 83049 -24126
rect 83093 -24170 83149 -24126
rect 83193 -24170 83249 -24126
rect 83293 -24170 83349 -24126
rect 83393 -24170 83449 -24126
rect 83493 -24170 83549 -24126
rect 83593 -24170 83649 -24126
rect 83693 -24170 83749 -24126
rect 83793 -24170 83849 -24126
rect 83893 -24170 83949 -24126
rect 83993 -24170 84049 -24126
rect 84093 -24170 84149 -24126
rect 84193 -24170 84249 -24126
rect 84293 -24170 84349 -24126
rect 84393 -24170 84849 -24126
rect 84893 -24170 84949 -24126
rect 84993 -24170 85049 -24126
rect 85093 -24170 85149 -24126
rect 85193 -24170 85249 -24126
rect 85293 -24170 85349 -24126
rect 85393 -24170 85449 -24126
rect 85493 -24170 85549 -24126
rect 85593 -24170 85649 -24126
rect 85693 -24170 85749 -24126
rect 85793 -24170 85849 -24126
rect 85893 -24170 85949 -24126
rect 85993 -24170 86049 -24126
rect 86093 -24170 86149 -24126
rect 86193 -24170 86249 -24126
rect 86293 -24170 86349 -24126
rect 86393 -24170 86849 -24126
rect 86893 -24170 86949 -24126
rect 86993 -24170 87049 -24126
rect 87093 -24170 87149 -24126
rect 87193 -24170 87249 -24126
rect 87293 -24170 87349 -24126
rect 87393 -24170 87449 -24126
rect 87493 -24170 87549 -24126
rect 87593 -24170 87649 -24126
rect 87693 -24170 87749 -24126
rect 87793 -24170 87849 -24126
rect 87893 -24170 87949 -24126
rect 87993 -24170 88049 -24126
rect 88093 -24170 88149 -24126
rect 88193 -24170 88249 -24126
rect 88293 -24170 88349 -24126
rect 88393 -24170 177360 -24126
rect -109116 -24195 177360 -24170
rect -109116 -24226 109104 -24195
rect -109116 -24270 80849 -24226
rect 80893 -24270 80949 -24226
rect 80993 -24270 81049 -24226
rect 81093 -24270 81149 -24226
rect 81193 -24270 81249 -24226
rect 81293 -24270 81349 -24226
rect 81393 -24270 81449 -24226
rect 81493 -24270 81549 -24226
rect 81593 -24270 81649 -24226
rect 81693 -24270 81749 -24226
rect 81793 -24270 81849 -24226
rect 81893 -24270 81949 -24226
rect 81993 -24270 82049 -24226
rect 82093 -24270 82149 -24226
rect 82193 -24270 82249 -24226
rect 82293 -24270 82349 -24226
rect 82393 -24270 82849 -24226
rect 82893 -24270 82949 -24226
rect 82993 -24270 83049 -24226
rect 83093 -24270 83149 -24226
rect 83193 -24270 83249 -24226
rect 83293 -24270 83349 -24226
rect 83393 -24270 83449 -24226
rect 83493 -24270 83549 -24226
rect 83593 -24270 83649 -24226
rect 83693 -24270 83749 -24226
rect 83793 -24270 83849 -24226
rect 83893 -24270 83949 -24226
rect 83993 -24270 84049 -24226
rect 84093 -24270 84149 -24226
rect 84193 -24270 84249 -24226
rect 84293 -24270 84349 -24226
rect 84393 -24270 84849 -24226
rect 84893 -24270 84949 -24226
rect 84993 -24270 85049 -24226
rect 85093 -24270 85149 -24226
rect 85193 -24270 85249 -24226
rect 85293 -24270 85349 -24226
rect 85393 -24270 85449 -24226
rect 85493 -24270 85549 -24226
rect 85593 -24270 85649 -24226
rect 85693 -24270 85749 -24226
rect 85793 -24270 85849 -24226
rect 85893 -24270 85949 -24226
rect 85993 -24270 86049 -24226
rect 86093 -24270 86149 -24226
rect 86193 -24270 86249 -24226
rect 86293 -24270 86349 -24226
rect 86393 -24270 86849 -24226
rect 86893 -24270 86949 -24226
rect 86993 -24270 87049 -24226
rect 87093 -24270 87149 -24226
rect 87193 -24270 87249 -24226
rect 87293 -24270 87349 -24226
rect 87393 -24270 87449 -24226
rect 87493 -24270 87549 -24226
rect 87593 -24270 87649 -24226
rect 87693 -24270 87749 -24226
rect 87793 -24270 87849 -24226
rect 87893 -24270 87949 -24226
rect 87993 -24270 88049 -24226
rect 88093 -24270 88149 -24226
rect 88193 -24270 88249 -24226
rect 88293 -24270 88349 -24226
rect 88393 -24239 109104 -24226
rect 109148 -24239 109204 -24195
rect 109248 -24239 109304 -24195
rect 109348 -24239 109404 -24195
rect 109448 -24239 109504 -24195
rect 109548 -24239 109604 -24195
rect 109648 -24239 109704 -24195
rect 109748 -24239 109804 -24195
rect 109848 -24239 109904 -24195
rect 109948 -24239 110004 -24195
rect 110048 -24239 110104 -24195
rect 110148 -24239 110204 -24195
rect 110248 -24239 110304 -24195
rect 110348 -24239 110404 -24195
rect 110448 -24239 110504 -24195
rect 110548 -24239 110604 -24195
rect 110648 -24239 111104 -24195
rect 111148 -24239 111204 -24195
rect 111248 -24239 111304 -24195
rect 111348 -24239 111404 -24195
rect 111448 -24239 111504 -24195
rect 111548 -24239 111604 -24195
rect 111648 -24239 111704 -24195
rect 111748 -24239 111804 -24195
rect 111848 -24239 111904 -24195
rect 111948 -24239 112004 -24195
rect 112048 -24239 112104 -24195
rect 112148 -24239 112204 -24195
rect 112248 -24239 112304 -24195
rect 112348 -24239 112404 -24195
rect 112448 -24239 112504 -24195
rect 112548 -24239 112604 -24195
rect 112648 -24239 113104 -24195
rect 113148 -24239 113204 -24195
rect 113248 -24239 113304 -24195
rect 113348 -24239 113404 -24195
rect 113448 -24239 113504 -24195
rect 113548 -24239 113604 -24195
rect 113648 -24239 113704 -24195
rect 113748 -24239 113804 -24195
rect 113848 -24239 113904 -24195
rect 113948 -24239 114004 -24195
rect 114048 -24239 114104 -24195
rect 114148 -24239 114204 -24195
rect 114248 -24239 114304 -24195
rect 114348 -24239 114404 -24195
rect 114448 -24239 114504 -24195
rect 114548 -24239 114604 -24195
rect 114648 -24239 115104 -24195
rect 115148 -24239 115204 -24195
rect 115248 -24239 115304 -24195
rect 115348 -24239 115404 -24195
rect 115448 -24239 115504 -24195
rect 115548 -24239 115604 -24195
rect 115648 -24239 115704 -24195
rect 115748 -24239 115804 -24195
rect 115848 -24239 115904 -24195
rect 115948 -24239 116004 -24195
rect 116048 -24239 116104 -24195
rect 116148 -24239 116204 -24195
rect 116248 -24239 116304 -24195
rect 116348 -24239 116404 -24195
rect 116448 -24239 116504 -24195
rect 116548 -24239 116604 -24195
rect 116648 -24239 177360 -24195
rect 88393 -24270 177360 -24239
rect -109116 -24295 177360 -24270
rect -109116 -24326 109104 -24295
rect -109116 -24366 80849 -24326
rect -109116 -24410 -82799 -24366
rect -82755 -24410 -82699 -24366
rect -82655 -24410 -82599 -24366
rect -82555 -24410 -82499 -24366
rect -82455 -24410 -82399 -24366
rect -82355 -24410 -82299 -24366
rect -82255 -24410 -82199 -24366
rect -82155 -24410 -82099 -24366
rect -82055 -24410 -81999 -24366
rect -81955 -24410 -81899 -24366
rect -81855 -24410 -81799 -24366
rect -81755 -24410 -81699 -24366
rect -81655 -24410 -81599 -24366
rect -81555 -24410 -81499 -24366
rect -81455 -24410 -81399 -24366
rect -81355 -24410 -81299 -24366
rect -81255 -24410 -80799 -24366
rect -80755 -24410 -80699 -24366
rect -80655 -24410 -80599 -24366
rect -80555 -24410 -80499 -24366
rect -80455 -24410 -80399 -24366
rect -80355 -24410 -80299 -24366
rect -80255 -24410 -80199 -24366
rect -80155 -24410 -80099 -24366
rect -80055 -24410 -79999 -24366
rect -79955 -24410 -79899 -24366
rect -79855 -24410 -79799 -24366
rect -79755 -24410 -79699 -24366
rect -79655 -24410 -79599 -24366
rect -79555 -24410 -79499 -24366
rect -79455 -24410 -79399 -24366
rect -79355 -24410 -79299 -24366
rect -79255 -24410 -78799 -24366
rect -78755 -24410 -78699 -24366
rect -78655 -24410 -78599 -24366
rect -78555 -24410 -78499 -24366
rect -78455 -24410 -78399 -24366
rect -78355 -24410 -78299 -24366
rect -78255 -24410 -78199 -24366
rect -78155 -24410 -78099 -24366
rect -78055 -24410 -77999 -24366
rect -77955 -24410 -77899 -24366
rect -77855 -24410 -77799 -24366
rect -77755 -24410 -77699 -24366
rect -77655 -24410 -77599 -24366
rect -77555 -24410 -77499 -24366
rect -77455 -24410 -77399 -24366
rect -77355 -24410 -77299 -24366
rect -77255 -24410 -76799 -24366
rect -76755 -24410 -76699 -24366
rect -76655 -24410 -76599 -24366
rect -76555 -24410 -76499 -24366
rect -76455 -24410 -76399 -24366
rect -76355 -24410 -76299 -24366
rect -76255 -24410 -76199 -24366
rect -76155 -24410 -76099 -24366
rect -76055 -24410 -75999 -24366
rect -75955 -24410 -75899 -24366
rect -75855 -24410 -75799 -24366
rect -75755 -24410 -75699 -24366
rect -75655 -24410 -75599 -24366
rect -75555 -24410 -75499 -24366
rect -75455 -24410 -75399 -24366
rect -75355 -24410 -75299 -24366
rect -75255 -24370 80849 -24366
rect 80893 -24370 80949 -24326
rect 80993 -24370 81049 -24326
rect 81093 -24370 81149 -24326
rect 81193 -24370 81249 -24326
rect 81293 -24370 81349 -24326
rect 81393 -24370 81449 -24326
rect 81493 -24370 81549 -24326
rect 81593 -24370 81649 -24326
rect 81693 -24370 81749 -24326
rect 81793 -24370 81849 -24326
rect 81893 -24370 81949 -24326
rect 81993 -24370 82049 -24326
rect 82093 -24370 82149 -24326
rect 82193 -24370 82249 -24326
rect 82293 -24370 82349 -24326
rect 82393 -24370 82849 -24326
rect 82893 -24370 82949 -24326
rect 82993 -24370 83049 -24326
rect 83093 -24370 83149 -24326
rect 83193 -24370 83249 -24326
rect 83293 -24370 83349 -24326
rect 83393 -24370 83449 -24326
rect 83493 -24370 83549 -24326
rect 83593 -24370 83649 -24326
rect 83693 -24370 83749 -24326
rect 83793 -24370 83849 -24326
rect 83893 -24370 83949 -24326
rect 83993 -24370 84049 -24326
rect 84093 -24370 84149 -24326
rect 84193 -24370 84249 -24326
rect 84293 -24370 84349 -24326
rect 84393 -24370 84849 -24326
rect 84893 -24370 84949 -24326
rect 84993 -24370 85049 -24326
rect 85093 -24370 85149 -24326
rect 85193 -24370 85249 -24326
rect 85293 -24370 85349 -24326
rect 85393 -24370 85449 -24326
rect 85493 -24370 85549 -24326
rect 85593 -24370 85649 -24326
rect 85693 -24370 85749 -24326
rect 85793 -24370 85849 -24326
rect 85893 -24370 85949 -24326
rect 85993 -24370 86049 -24326
rect 86093 -24370 86149 -24326
rect 86193 -24370 86249 -24326
rect 86293 -24370 86349 -24326
rect 86393 -24370 86849 -24326
rect 86893 -24370 86949 -24326
rect 86993 -24370 87049 -24326
rect 87093 -24370 87149 -24326
rect 87193 -24370 87249 -24326
rect 87293 -24370 87349 -24326
rect 87393 -24370 87449 -24326
rect 87493 -24370 87549 -24326
rect 87593 -24370 87649 -24326
rect 87693 -24370 87749 -24326
rect 87793 -24370 87849 -24326
rect 87893 -24370 87949 -24326
rect 87993 -24370 88049 -24326
rect 88093 -24370 88149 -24326
rect 88193 -24370 88249 -24326
rect 88293 -24370 88349 -24326
rect 88393 -24339 109104 -24326
rect 109148 -24339 109204 -24295
rect 109248 -24339 109304 -24295
rect 109348 -24339 109404 -24295
rect 109448 -24339 109504 -24295
rect 109548 -24339 109604 -24295
rect 109648 -24339 109704 -24295
rect 109748 -24339 109804 -24295
rect 109848 -24339 109904 -24295
rect 109948 -24339 110004 -24295
rect 110048 -24339 110104 -24295
rect 110148 -24339 110204 -24295
rect 110248 -24339 110304 -24295
rect 110348 -24339 110404 -24295
rect 110448 -24339 110504 -24295
rect 110548 -24339 110604 -24295
rect 110648 -24339 111104 -24295
rect 111148 -24339 111204 -24295
rect 111248 -24339 111304 -24295
rect 111348 -24339 111404 -24295
rect 111448 -24339 111504 -24295
rect 111548 -24339 111604 -24295
rect 111648 -24339 111704 -24295
rect 111748 -24339 111804 -24295
rect 111848 -24339 111904 -24295
rect 111948 -24339 112004 -24295
rect 112048 -24339 112104 -24295
rect 112148 -24339 112204 -24295
rect 112248 -24339 112304 -24295
rect 112348 -24339 112404 -24295
rect 112448 -24339 112504 -24295
rect 112548 -24339 112604 -24295
rect 112648 -24339 113104 -24295
rect 113148 -24339 113204 -24295
rect 113248 -24339 113304 -24295
rect 113348 -24339 113404 -24295
rect 113448 -24339 113504 -24295
rect 113548 -24339 113604 -24295
rect 113648 -24339 113704 -24295
rect 113748 -24339 113804 -24295
rect 113848 -24339 113904 -24295
rect 113948 -24339 114004 -24295
rect 114048 -24339 114104 -24295
rect 114148 -24339 114204 -24295
rect 114248 -24339 114304 -24295
rect 114348 -24339 114404 -24295
rect 114448 -24339 114504 -24295
rect 114548 -24339 114604 -24295
rect 114648 -24339 115104 -24295
rect 115148 -24339 115204 -24295
rect 115248 -24339 115304 -24295
rect 115348 -24339 115404 -24295
rect 115448 -24339 115504 -24295
rect 115548 -24339 115604 -24295
rect 115648 -24339 115704 -24295
rect 115748 -24339 115804 -24295
rect 115848 -24339 115904 -24295
rect 115948 -24339 116004 -24295
rect 116048 -24339 116104 -24295
rect 116148 -24339 116204 -24295
rect 116248 -24339 116304 -24295
rect 116348 -24339 116404 -24295
rect 116448 -24339 116504 -24295
rect 116548 -24339 116604 -24295
rect 116648 -24339 177360 -24295
rect 88393 -24370 177360 -24339
rect -75255 -24395 177360 -24370
rect -75255 -24410 109104 -24395
rect -109116 -24426 109104 -24410
rect -109116 -24466 80849 -24426
rect -109116 -24510 -82799 -24466
rect -82755 -24510 -82699 -24466
rect -82655 -24510 -82599 -24466
rect -82555 -24510 -82499 -24466
rect -82455 -24510 -82399 -24466
rect -82355 -24510 -82299 -24466
rect -82255 -24510 -82199 -24466
rect -82155 -24510 -82099 -24466
rect -82055 -24510 -81999 -24466
rect -81955 -24510 -81899 -24466
rect -81855 -24510 -81799 -24466
rect -81755 -24510 -81699 -24466
rect -81655 -24510 -81599 -24466
rect -81555 -24510 -81499 -24466
rect -81455 -24510 -81399 -24466
rect -81355 -24510 -81299 -24466
rect -81255 -24510 -80799 -24466
rect -80755 -24510 -80699 -24466
rect -80655 -24510 -80599 -24466
rect -80555 -24510 -80499 -24466
rect -80455 -24510 -80399 -24466
rect -80355 -24510 -80299 -24466
rect -80255 -24510 -80199 -24466
rect -80155 -24510 -80099 -24466
rect -80055 -24510 -79999 -24466
rect -79955 -24510 -79899 -24466
rect -79855 -24510 -79799 -24466
rect -79755 -24510 -79699 -24466
rect -79655 -24510 -79599 -24466
rect -79555 -24510 -79499 -24466
rect -79455 -24510 -79399 -24466
rect -79355 -24510 -79299 -24466
rect -79255 -24510 -78799 -24466
rect -78755 -24510 -78699 -24466
rect -78655 -24510 -78599 -24466
rect -78555 -24510 -78499 -24466
rect -78455 -24510 -78399 -24466
rect -78355 -24510 -78299 -24466
rect -78255 -24510 -78199 -24466
rect -78155 -24510 -78099 -24466
rect -78055 -24510 -77999 -24466
rect -77955 -24510 -77899 -24466
rect -77855 -24510 -77799 -24466
rect -77755 -24510 -77699 -24466
rect -77655 -24510 -77599 -24466
rect -77555 -24510 -77499 -24466
rect -77455 -24510 -77399 -24466
rect -77355 -24510 -77299 -24466
rect -77255 -24510 -76799 -24466
rect -76755 -24510 -76699 -24466
rect -76655 -24510 -76599 -24466
rect -76555 -24510 -76499 -24466
rect -76455 -24510 -76399 -24466
rect -76355 -24510 -76299 -24466
rect -76255 -24510 -76199 -24466
rect -76155 -24510 -76099 -24466
rect -76055 -24510 -75999 -24466
rect -75955 -24510 -75899 -24466
rect -75855 -24510 -75799 -24466
rect -75755 -24510 -75699 -24466
rect -75655 -24510 -75599 -24466
rect -75555 -24510 -75499 -24466
rect -75455 -24510 -75399 -24466
rect -75355 -24510 -75299 -24466
rect -75255 -24470 80849 -24466
rect 80893 -24470 80949 -24426
rect 80993 -24470 81049 -24426
rect 81093 -24470 81149 -24426
rect 81193 -24470 81249 -24426
rect 81293 -24470 81349 -24426
rect 81393 -24470 81449 -24426
rect 81493 -24470 81549 -24426
rect 81593 -24470 81649 -24426
rect 81693 -24470 81749 -24426
rect 81793 -24470 81849 -24426
rect 81893 -24470 81949 -24426
rect 81993 -24470 82049 -24426
rect 82093 -24470 82149 -24426
rect 82193 -24470 82249 -24426
rect 82293 -24470 82349 -24426
rect 82393 -24470 82849 -24426
rect 82893 -24470 82949 -24426
rect 82993 -24470 83049 -24426
rect 83093 -24470 83149 -24426
rect 83193 -24470 83249 -24426
rect 83293 -24470 83349 -24426
rect 83393 -24470 83449 -24426
rect 83493 -24470 83549 -24426
rect 83593 -24470 83649 -24426
rect 83693 -24470 83749 -24426
rect 83793 -24470 83849 -24426
rect 83893 -24470 83949 -24426
rect 83993 -24470 84049 -24426
rect 84093 -24470 84149 -24426
rect 84193 -24470 84249 -24426
rect 84293 -24470 84349 -24426
rect 84393 -24470 84849 -24426
rect 84893 -24470 84949 -24426
rect 84993 -24470 85049 -24426
rect 85093 -24470 85149 -24426
rect 85193 -24470 85249 -24426
rect 85293 -24470 85349 -24426
rect 85393 -24470 85449 -24426
rect 85493 -24470 85549 -24426
rect 85593 -24470 85649 -24426
rect 85693 -24470 85749 -24426
rect 85793 -24470 85849 -24426
rect 85893 -24470 85949 -24426
rect 85993 -24470 86049 -24426
rect 86093 -24470 86149 -24426
rect 86193 -24470 86249 -24426
rect 86293 -24470 86349 -24426
rect 86393 -24470 86849 -24426
rect 86893 -24470 86949 -24426
rect 86993 -24470 87049 -24426
rect 87093 -24470 87149 -24426
rect 87193 -24470 87249 -24426
rect 87293 -24470 87349 -24426
rect 87393 -24470 87449 -24426
rect 87493 -24470 87549 -24426
rect 87593 -24470 87649 -24426
rect 87693 -24470 87749 -24426
rect 87793 -24470 87849 -24426
rect 87893 -24470 87949 -24426
rect 87993 -24470 88049 -24426
rect 88093 -24470 88149 -24426
rect 88193 -24470 88249 -24426
rect 88293 -24470 88349 -24426
rect 88393 -24439 109104 -24426
rect 109148 -24439 109204 -24395
rect 109248 -24439 109304 -24395
rect 109348 -24439 109404 -24395
rect 109448 -24439 109504 -24395
rect 109548 -24439 109604 -24395
rect 109648 -24439 109704 -24395
rect 109748 -24439 109804 -24395
rect 109848 -24439 109904 -24395
rect 109948 -24439 110004 -24395
rect 110048 -24439 110104 -24395
rect 110148 -24439 110204 -24395
rect 110248 -24439 110304 -24395
rect 110348 -24439 110404 -24395
rect 110448 -24439 110504 -24395
rect 110548 -24439 110604 -24395
rect 110648 -24439 111104 -24395
rect 111148 -24439 111204 -24395
rect 111248 -24439 111304 -24395
rect 111348 -24439 111404 -24395
rect 111448 -24439 111504 -24395
rect 111548 -24439 111604 -24395
rect 111648 -24439 111704 -24395
rect 111748 -24439 111804 -24395
rect 111848 -24439 111904 -24395
rect 111948 -24439 112004 -24395
rect 112048 -24439 112104 -24395
rect 112148 -24439 112204 -24395
rect 112248 -24439 112304 -24395
rect 112348 -24439 112404 -24395
rect 112448 -24439 112504 -24395
rect 112548 -24439 112604 -24395
rect 112648 -24439 113104 -24395
rect 113148 -24439 113204 -24395
rect 113248 -24439 113304 -24395
rect 113348 -24439 113404 -24395
rect 113448 -24439 113504 -24395
rect 113548 -24439 113604 -24395
rect 113648 -24439 113704 -24395
rect 113748 -24439 113804 -24395
rect 113848 -24439 113904 -24395
rect 113948 -24439 114004 -24395
rect 114048 -24439 114104 -24395
rect 114148 -24439 114204 -24395
rect 114248 -24439 114304 -24395
rect 114348 -24439 114404 -24395
rect 114448 -24439 114504 -24395
rect 114548 -24439 114604 -24395
rect 114648 -24439 115104 -24395
rect 115148 -24439 115204 -24395
rect 115248 -24439 115304 -24395
rect 115348 -24439 115404 -24395
rect 115448 -24439 115504 -24395
rect 115548 -24439 115604 -24395
rect 115648 -24439 115704 -24395
rect 115748 -24439 115804 -24395
rect 115848 -24439 115904 -24395
rect 115948 -24439 116004 -24395
rect 116048 -24439 116104 -24395
rect 116148 -24439 116204 -24395
rect 116248 -24439 116304 -24395
rect 116348 -24439 116404 -24395
rect 116448 -24439 116504 -24395
rect 116548 -24439 116604 -24395
rect 116648 -24439 177360 -24395
rect 88393 -24470 177360 -24439
rect -75255 -24495 177360 -24470
rect -75255 -24510 109104 -24495
rect -109116 -24526 109104 -24510
rect -109116 -24566 80849 -24526
rect -109116 -24610 -82799 -24566
rect -82755 -24610 -82699 -24566
rect -82655 -24610 -82599 -24566
rect -82555 -24610 -82499 -24566
rect -82455 -24610 -82399 -24566
rect -82355 -24610 -82299 -24566
rect -82255 -24610 -82199 -24566
rect -82155 -24610 -82099 -24566
rect -82055 -24610 -81999 -24566
rect -81955 -24610 -81899 -24566
rect -81855 -24610 -81799 -24566
rect -81755 -24610 -81699 -24566
rect -81655 -24610 -81599 -24566
rect -81555 -24610 -81499 -24566
rect -81455 -24610 -81399 -24566
rect -81355 -24610 -81299 -24566
rect -81255 -24610 -80799 -24566
rect -80755 -24610 -80699 -24566
rect -80655 -24610 -80599 -24566
rect -80555 -24610 -80499 -24566
rect -80455 -24610 -80399 -24566
rect -80355 -24610 -80299 -24566
rect -80255 -24610 -80199 -24566
rect -80155 -24610 -80099 -24566
rect -80055 -24610 -79999 -24566
rect -79955 -24610 -79899 -24566
rect -79855 -24610 -79799 -24566
rect -79755 -24610 -79699 -24566
rect -79655 -24610 -79599 -24566
rect -79555 -24610 -79499 -24566
rect -79455 -24610 -79399 -24566
rect -79355 -24610 -79299 -24566
rect -79255 -24610 -78799 -24566
rect -78755 -24610 -78699 -24566
rect -78655 -24610 -78599 -24566
rect -78555 -24610 -78499 -24566
rect -78455 -24610 -78399 -24566
rect -78355 -24610 -78299 -24566
rect -78255 -24610 -78199 -24566
rect -78155 -24610 -78099 -24566
rect -78055 -24610 -77999 -24566
rect -77955 -24610 -77899 -24566
rect -77855 -24610 -77799 -24566
rect -77755 -24610 -77699 -24566
rect -77655 -24610 -77599 -24566
rect -77555 -24610 -77499 -24566
rect -77455 -24610 -77399 -24566
rect -77355 -24610 -77299 -24566
rect -77255 -24610 -76799 -24566
rect -76755 -24610 -76699 -24566
rect -76655 -24610 -76599 -24566
rect -76555 -24610 -76499 -24566
rect -76455 -24610 -76399 -24566
rect -76355 -24610 -76299 -24566
rect -76255 -24610 -76199 -24566
rect -76155 -24610 -76099 -24566
rect -76055 -24610 -75999 -24566
rect -75955 -24610 -75899 -24566
rect -75855 -24610 -75799 -24566
rect -75755 -24610 -75699 -24566
rect -75655 -24610 -75599 -24566
rect -75555 -24610 -75499 -24566
rect -75455 -24610 -75399 -24566
rect -75355 -24610 -75299 -24566
rect -75255 -24570 80849 -24566
rect 80893 -24570 80949 -24526
rect 80993 -24570 81049 -24526
rect 81093 -24570 81149 -24526
rect 81193 -24570 81249 -24526
rect 81293 -24570 81349 -24526
rect 81393 -24570 81449 -24526
rect 81493 -24570 81549 -24526
rect 81593 -24570 81649 -24526
rect 81693 -24570 81749 -24526
rect 81793 -24570 81849 -24526
rect 81893 -24570 81949 -24526
rect 81993 -24570 82049 -24526
rect 82093 -24570 82149 -24526
rect 82193 -24570 82249 -24526
rect 82293 -24570 82349 -24526
rect 82393 -24570 82849 -24526
rect 82893 -24570 82949 -24526
rect 82993 -24570 83049 -24526
rect 83093 -24570 83149 -24526
rect 83193 -24570 83249 -24526
rect 83293 -24570 83349 -24526
rect 83393 -24570 83449 -24526
rect 83493 -24570 83549 -24526
rect 83593 -24570 83649 -24526
rect 83693 -24570 83749 -24526
rect 83793 -24570 83849 -24526
rect 83893 -24570 83949 -24526
rect 83993 -24570 84049 -24526
rect 84093 -24570 84149 -24526
rect 84193 -24570 84249 -24526
rect 84293 -24570 84349 -24526
rect 84393 -24570 84849 -24526
rect 84893 -24570 84949 -24526
rect 84993 -24570 85049 -24526
rect 85093 -24570 85149 -24526
rect 85193 -24570 85249 -24526
rect 85293 -24570 85349 -24526
rect 85393 -24570 85449 -24526
rect 85493 -24570 85549 -24526
rect 85593 -24570 85649 -24526
rect 85693 -24570 85749 -24526
rect 85793 -24570 85849 -24526
rect 85893 -24570 85949 -24526
rect 85993 -24570 86049 -24526
rect 86093 -24570 86149 -24526
rect 86193 -24570 86249 -24526
rect 86293 -24570 86349 -24526
rect 86393 -24570 86849 -24526
rect 86893 -24570 86949 -24526
rect 86993 -24570 87049 -24526
rect 87093 -24570 87149 -24526
rect 87193 -24570 87249 -24526
rect 87293 -24570 87349 -24526
rect 87393 -24570 87449 -24526
rect 87493 -24570 87549 -24526
rect 87593 -24570 87649 -24526
rect 87693 -24570 87749 -24526
rect 87793 -24570 87849 -24526
rect 87893 -24570 87949 -24526
rect 87993 -24570 88049 -24526
rect 88093 -24570 88149 -24526
rect 88193 -24570 88249 -24526
rect 88293 -24570 88349 -24526
rect 88393 -24539 109104 -24526
rect 109148 -24539 109204 -24495
rect 109248 -24539 109304 -24495
rect 109348 -24539 109404 -24495
rect 109448 -24539 109504 -24495
rect 109548 -24539 109604 -24495
rect 109648 -24539 109704 -24495
rect 109748 -24539 109804 -24495
rect 109848 -24539 109904 -24495
rect 109948 -24539 110004 -24495
rect 110048 -24539 110104 -24495
rect 110148 -24539 110204 -24495
rect 110248 -24539 110304 -24495
rect 110348 -24539 110404 -24495
rect 110448 -24539 110504 -24495
rect 110548 -24539 110604 -24495
rect 110648 -24539 111104 -24495
rect 111148 -24539 111204 -24495
rect 111248 -24539 111304 -24495
rect 111348 -24539 111404 -24495
rect 111448 -24539 111504 -24495
rect 111548 -24539 111604 -24495
rect 111648 -24539 111704 -24495
rect 111748 -24539 111804 -24495
rect 111848 -24539 111904 -24495
rect 111948 -24539 112004 -24495
rect 112048 -24539 112104 -24495
rect 112148 -24539 112204 -24495
rect 112248 -24539 112304 -24495
rect 112348 -24539 112404 -24495
rect 112448 -24539 112504 -24495
rect 112548 -24539 112604 -24495
rect 112648 -24539 113104 -24495
rect 113148 -24539 113204 -24495
rect 113248 -24539 113304 -24495
rect 113348 -24539 113404 -24495
rect 113448 -24539 113504 -24495
rect 113548 -24539 113604 -24495
rect 113648 -24539 113704 -24495
rect 113748 -24539 113804 -24495
rect 113848 -24539 113904 -24495
rect 113948 -24539 114004 -24495
rect 114048 -24539 114104 -24495
rect 114148 -24539 114204 -24495
rect 114248 -24539 114304 -24495
rect 114348 -24539 114404 -24495
rect 114448 -24539 114504 -24495
rect 114548 -24539 114604 -24495
rect 114648 -24539 115104 -24495
rect 115148 -24539 115204 -24495
rect 115248 -24539 115304 -24495
rect 115348 -24539 115404 -24495
rect 115448 -24539 115504 -24495
rect 115548 -24539 115604 -24495
rect 115648 -24539 115704 -24495
rect 115748 -24539 115804 -24495
rect 115848 -24539 115904 -24495
rect 115948 -24539 116004 -24495
rect 116048 -24539 116104 -24495
rect 116148 -24539 116204 -24495
rect 116248 -24539 116304 -24495
rect 116348 -24539 116404 -24495
rect 116448 -24539 116504 -24495
rect 116548 -24539 116604 -24495
rect 116648 -24539 177360 -24495
rect 88393 -24570 177360 -24539
rect -75255 -24595 177360 -24570
rect -75255 -24610 109104 -24595
rect -109116 -24626 109104 -24610
rect -109116 -24666 80849 -24626
rect -109116 -24710 -82799 -24666
rect -82755 -24710 -82699 -24666
rect -82655 -24710 -82599 -24666
rect -82555 -24710 -82499 -24666
rect -82455 -24710 -82399 -24666
rect -82355 -24710 -82299 -24666
rect -82255 -24710 -82199 -24666
rect -82155 -24710 -82099 -24666
rect -82055 -24710 -81999 -24666
rect -81955 -24710 -81899 -24666
rect -81855 -24710 -81799 -24666
rect -81755 -24710 -81699 -24666
rect -81655 -24710 -81599 -24666
rect -81555 -24710 -81499 -24666
rect -81455 -24710 -81399 -24666
rect -81355 -24710 -81299 -24666
rect -81255 -24710 -80799 -24666
rect -80755 -24710 -80699 -24666
rect -80655 -24710 -80599 -24666
rect -80555 -24710 -80499 -24666
rect -80455 -24710 -80399 -24666
rect -80355 -24710 -80299 -24666
rect -80255 -24710 -80199 -24666
rect -80155 -24710 -80099 -24666
rect -80055 -24710 -79999 -24666
rect -79955 -24710 -79899 -24666
rect -79855 -24710 -79799 -24666
rect -79755 -24710 -79699 -24666
rect -79655 -24710 -79599 -24666
rect -79555 -24710 -79499 -24666
rect -79455 -24710 -79399 -24666
rect -79355 -24710 -79299 -24666
rect -79255 -24710 -78799 -24666
rect -78755 -24710 -78699 -24666
rect -78655 -24710 -78599 -24666
rect -78555 -24710 -78499 -24666
rect -78455 -24710 -78399 -24666
rect -78355 -24710 -78299 -24666
rect -78255 -24710 -78199 -24666
rect -78155 -24710 -78099 -24666
rect -78055 -24710 -77999 -24666
rect -77955 -24710 -77899 -24666
rect -77855 -24710 -77799 -24666
rect -77755 -24710 -77699 -24666
rect -77655 -24710 -77599 -24666
rect -77555 -24710 -77499 -24666
rect -77455 -24710 -77399 -24666
rect -77355 -24710 -77299 -24666
rect -77255 -24710 -76799 -24666
rect -76755 -24710 -76699 -24666
rect -76655 -24710 -76599 -24666
rect -76555 -24710 -76499 -24666
rect -76455 -24710 -76399 -24666
rect -76355 -24710 -76299 -24666
rect -76255 -24710 -76199 -24666
rect -76155 -24710 -76099 -24666
rect -76055 -24710 -75999 -24666
rect -75955 -24710 -75899 -24666
rect -75855 -24710 -75799 -24666
rect -75755 -24710 -75699 -24666
rect -75655 -24710 -75599 -24666
rect -75555 -24710 -75499 -24666
rect -75455 -24710 -75399 -24666
rect -75355 -24710 -75299 -24666
rect -75255 -24670 80849 -24666
rect 80893 -24670 80949 -24626
rect 80993 -24670 81049 -24626
rect 81093 -24670 81149 -24626
rect 81193 -24670 81249 -24626
rect 81293 -24670 81349 -24626
rect 81393 -24670 81449 -24626
rect 81493 -24670 81549 -24626
rect 81593 -24670 81649 -24626
rect 81693 -24670 81749 -24626
rect 81793 -24670 81849 -24626
rect 81893 -24670 81949 -24626
rect 81993 -24670 82049 -24626
rect 82093 -24670 82149 -24626
rect 82193 -24670 82249 -24626
rect 82293 -24670 82349 -24626
rect 82393 -24670 82849 -24626
rect 82893 -24670 82949 -24626
rect 82993 -24670 83049 -24626
rect 83093 -24670 83149 -24626
rect 83193 -24670 83249 -24626
rect 83293 -24670 83349 -24626
rect 83393 -24670 83449 -24626
rect 83493 -24670 83549 -24626
rect 83593 -24670 83649 -24626
rect 83693 -24670 83749 -24626
rect 83793 -24670 83849 -24626
rect 83893 -24670 83949 -24626
rect 83993 -24670 84049 -24626
rect 84093 -24670 84149 -24626
rect 84193 -24670 84249 -24626
rect 84293 -24670 84349 -24626
rect 84393 -24670 84849 -24626
rect 84893 -24670 84949 -24626
rect 84993 -24670 85049 -24626
rect 85093 -24670 85149 -24626
rect 85193 -24670 85249 -24626
rect 85293 -24670 85349 -24626
rect 85393 -24670 85449 -24626
rect 85493 -24670 85549 -24626
rect 85593 -24670 85649 -24626
rect 85693 -24670 85749 -24626
rect 85793 -24670 85849 -24626
rect 85893 -24670 85949 -24626
rect 85993 -24670 86049 -24626
rect 86093 -24670 86149 -24626
rect 86193 -24670 86249 -24626
rect 86293 -24670 86349 -24626
rect 86393 -24670 86849 -24626
rect 86893 -24670 86949 -24626
rect 86993 -24670 87049 -24626
rect 87093 -24670 87149 -24626
rect 87193 -24670 87249 -24626
rect 87293 -24670 87349 -24626
rect 87393 -24670 87449 -24626
rect 87493 -24670 87549 -24626
rect 87593 -24670 87649 -24626
rect 87693 -24670 87749 -24626
rect 87793 -24670 87849 -24626
rect 87893 -24670 87949 -24626
rect 87993 -24670 88049 -24626
rect 88093 -24670 88149 -24626
rect 88193 -24670 88249 -24626
rect 88293 -24670 88349 -24626
rect 88393 -24639 109104 -24626
rect 109148 -24639 109204 -24595
rect 109248 -24639 109304 -24595
rect 109348 -24639 109404 -24595
rect 109448 -24639 109504 -24595
rect 109548 -24639 109604 -24595
rect 109648 -24639 109704 -24595
rect 109748 -24639 109804 -24595
rect 109848 -24639 109904 -24595
rect 109948 -24639 110004 -24595
rect 110048 -24639 110104 -24595
rect 110148 -24639 110204 -24595
rect 110248 -24639 110304 -24595
rect 110348 -24639 110404 -24595
rect 110448 -24639 110504 -24595
rect 110548 -24639 110604 -24595
rect 110648 -24639 111104 -24595
rect 111148 -24639 111204 -24595
rect 111248 -24639 111304 -24595
rect 111348 -24639 111404 -24595
rect 111448 -24639 111504 -24595
rect 111548 -24639 111604 -24595
rect 111648 -24639 111704 -24595
rect 111748 -24639 111804 -24595
rect 111848 -24639 111904 -24595
rect 111948 -24639 112004 -24595
rect 112048 -24639 112104 -24595
rect 112148 -24639 112204 -24595
rect 112248 -24639 112304 -24595
rect 112348 -24639 112404 -24595
rect 112448 -24639 112504 -24595
rect 112548 -24639 112604 -24595
rect 112648 -24639 113104 -24595
rect 113148 -24639 113204 -24595
rect 113248 -24639 113304 -24595
rect 113348 -24639 113404 -24595
rect 113448 -24639 113504 -24595
rect 113548 -24639 113604 -24595
rect 113648 -24639 113704 -24595
rect 113748 -24639 113804 -24595
rect 113848 -24639 113904 -24595
rect 113948 -24639 114004 -24595
rect 114048 -24639 114104 -24595
rect 114148 -24639 114204 -24595
rect 114248 -24639 114304 -24595
rect 114348 -24639 114404 -24595
rect 114448 -24639 114504 -24595
rect 114548 -24639 114604 -24595
rect 114648 -24639 115104 -24595
rect 115148 -24639 115204 -24595
rect 115248 -24639 115304 -24595
rect 115348 -24639 115404 -24595
rect 115448 -24639 115504 -24595
rect 115548 -24639 115604 -24595
rect 115648 -24639 115704 -24595
rect 115748 -24639 115804 -24595
rect 115848 -24639 115904 -24595
rect 115948 -24639 116004 -24595
rect 116048 -24639 116104 -24595
rect 116148 -24639 116204 -24595
rect 116248 -24639 116304 -24595
rect 116348 -24639 116404 -24595
rect 116448 -24639 116504 -24595
rect 116548 -24639 116604 -24595
rect 116648 -24639 177360 -24595
rect 88393 -24670 177360 -24639
rect -75255 -24695 177360 -24670
rect -75255 -24710 109104 -24695
rect -109116 -24726 109104 -24710
rect -109116 -24766 80849 -24726
rect -109116 -24810 -82799 -24766
rect -82755 -24810 -82699 -24766
rect -82655 -24810 -82599 -24766
rect -82555 -24810 -82499 -24766
rect -82455 -24810 -82399 -24766
rect -82355 -24810 -82299 -24766
rect -82255 -24810 -82199 -24766
rect -82155 -24810 -82099 -24766
rect -82055 -24810 -81999 -24766
rect -81955 -24810 -81899 -24766
rect -81855 -24810 -81799 -24766
rect -81755 -24810 -81699 -24766
rect -81655 -24810 -81599 -24766
rect -81555 -24810 -81499 -24766
rect -81455 -24810 -81399 -24766
rect -81355 -24810 -81299 -24766
rect -81255 -24810 -80799 -24766
rect -80755 -24810 -80699 -24766
rect -80655 -24810 -80599 -24766
rect -80555 -24810 -80499 -24766
rect -80455 -24810 -80399 -24766
rect -80355 -24810 -80299 -24766
rect -80255 -24810 -80199 -24766
rect -80155 -24810 -80099 -24766
rect -80055 -24810 -79999 -24766
rect -79955 -24810 -79899 -24766
rect -79855 -24810 -79799 -24766
rect -79755 -24810 -79699 -24766
rect -79655 -24810 -79599 -24766
rect -79555 -24810 -79499 -24766
rect -79455 -24810 -79399 -24766
rect -79355 -24810 -79299 -24766
rect -79255 -24810 -78799 -24766
rect -78755 -24810 -78699 -24766
rect -78655 -24810 -78599 -24766
rect -78555 -24810 -78499 -24766
rect -78455 -24810 -78399 -24766
rect -78355 -24810 -78299 -24766
rect -78255 -24810 -78199 -24766
rect -78155 -24810 -78099 -24766
rect -78055 -24810 -77999 -24766
rect -77955 -24810 -77899 -24766
rect -77855 -24810 -77799 -24766
rect -77755 -24810 -77699 -24766
rect -77655 -24810 -77599 -24766
rect -77555 -24810 -77499 -24766
rect -77455 -24810 -77399 -24766
rect -77355 -24810 -77299 -24766
rect -77255 -24810 -76799 -24766
rect -76755 -24810 -76699 -24766
rect -76655 -24810 -76599 -24766
rect -76555 -24810 -76499 -24766
rect -76455 -24810 -76399 -24766
rect -76355 -24810 -76299 -24766
rect -76255 -24810 -76199 -24766
rect -76155 -24810 -76099 -24766
rect -76055 -24810 -75999 -24766
rect -75955 -24810 -75899 -24766
rect -75855 -24810 -75799 -24766
rect -75755 -24810 -75699 -24766
rect -75655 -24810 -75599 -24766
rect -75555 -24810 -75499 -24766
rect -75455 -24810 -75399 -24766
rect -75355 -24810 -75299 -24766
rect -75255 -24770 80849 -24766
rect 80893 -24770 80949 -24726
rect 80993 -24770 81049 -24726
rect 81093 -24770 81149 -24726
rect 81193 -24770 81249 -24726
rect 81293 -24770 81349 -24726
rect 81393 -24770 81449 -24726
rect 81493 -24770 81549 -24726
rect 81593 -24770 81649 -24726
rect 81693 -24770 81749 -24726
rect 81793 -24770 81849 -24726
rect 81893 -24770 81949 -24726
rect 81993 -24770 82049 -24726
rect 82093 -24770 82149 -24726
rect 82193 -24770 82249 -24726
rect 82293 -24770 82349 -24726
rect 82393 -24770 82849 -24726
rect 82893 -24770 82949 -24726
rect 82993 -24770 83049 -24726
rect 83093 -24770 83149 -24726
rect 83193 -24770 83249 -24726
rect 83293 -24770 83349 -24726
rect 83393 -24770 83449 -24726
rect 83493 -24770 83549 -24726
rect 83593 -24770 83649 -24726
rect 83693 -24770 83749 -24726
rect 83793 -24770 83849 -24726
rect 83893 -24770 83949 -24726
rect 83993 -24770 84049 -24726
rect 84093 -24770 84149 -24726
rect 84193 -24770 84249 -24726
rect 84293 -24770 84349 -24726
rect 84393 -24770 84849 -24726
rect 84893 -24770 84949 -24726
rect 84993 -24770 85049 -24726
rect 85093 -24770 85149 -24726
rect 85193 -24770 85249 -24726
rect 85293 -24770 85349 -24726
rect 85393 -24770 85449 -24726
rect 85493 -24770 85549 -24726
rect 85593 -24770 85649 -24726
rect 85693 -24770 85749 -24726
rect 85793 -24770 85849 -24726
rect 85893 -24770 85949 -24726
rect 85993 -24770 86049 -24726
rect 86093 -24770 86149 -24726
rect 86193 -24770 86249 -24726
rect 86293 -24770 86349 -24726
rect 86393 -24770 86849 -24726
rect 86893 -24770 86949 -24726
rect 86993 -24770 87049 -24726
rect 87093 -24770 87149 -24726
rect 87193 -24770 87249 -24726
rect 87293 -24770 87349 -24726
rect 87393 -24770 87449 -24726
rect 87493 -24770 87549 -24726
rect 87593 -24770 87649 -24726
rect 87693 -24770 87749 -24726
rect 87793 -24770 87849 -24726
rect 87893 -24770 87949 -24726
rect 87993 -24770 88049 -24726
rect 88093 -24770 88149 -24726
rect 88193 -24770 88249 -24726
rect 88293 -24770 88349 -24726
rect 88393 -24739 109104 -24726
rect 109148 -24739 109204 -24695
rect 109248 -24739 109304 -24695
rect 109348 -24739 109404 -24695
rect 109448 -24739 109504 -24695
rect 109548 -24739 109604 -24695
rect 109648 -24739 109704 -24695
rect 109748 -24739 109804 -24695
rect 109848 -24739 109904 -24695
rect 109948 -24739 110004 -24695
rect 110048 -24739 110104 -24695
rect 110148 -24739 110204 -24695
rect 110248 -24739 110304 -24695
rect 110348 -24739 110404 -24695
rect 110448 -24739 110504 -24695
rect 110548 -24739 110604 -24695
rect 110648 -24739 111104 -24695
rect 111148 -24739 111204 -24695
rect 111248 -24739 111304 -24695
rect 111348 -24739 111404 -24695
rect 111448 -24739 111504 -24695
rect 111548 -24739 111604 -24695
rect 111648 -24739 111704 -24695
rect 111748 -24739 111804 -24695
rect 111848 -24739 111904 -24695
rect 111948 -24739 112004 -24695
rect 112048 -24739 112104 -24695
rect 112148 -24739 112204 -24695
rect 112248 -24739 112304 -24695
rect 112348 -24739 112404 -24695
rect 112448 -24739 112504 -24695
rect 112548 -24739 112604 -24695
rect 112648 -24739 113104 -24695
rect 113148 -24739 113204 -24695
rect 113248 -24739 113304 -24695
rect 113348 -24739 113404 -24695
rect 113448 -24739 113504 -24695
rect 113548 -24739 113604 -24695
rect 113648 -24739 113704 -24695
rect 113748 -24739 113804 -24695
rect 113848 -24739 113904 -24695
rect 113948 -24739 114004 -24695
rect 114048 -24739 114104 -24695
rect 114148 -24739 114204 -24695
rect 114248 -24739 114304 -24695
rect 114348 -24739 114404 -24695
rect 114448 -24739 114504 -24695
rect 114548 -24739 114604 -24695
rect 114648 -24739 115104 -24695
rect 115148 -24739 115204 -24695
rect 115248 -24739 115304 -24695
rect 115348 -24739 115404 -24695
rect 115448 -24739 115504 -24695
rect 115548 -24739 115604 -24695
rect 115648 -24739 115704 -24695
rect 115748 -24739 115804 -24695
rect 115848 -24739 115904 -24695
rect 115948 -24739 116004 -24695
rect 116048 -24739 116104 -24695
rect 116148 -24739 116204 -24695
rect 116248 -24739 116304 -24695
rect 116348 -24739 116404 -24695
rect 116448 -24739 116504 -24695
rect 116548 -24739 116604 -24695
rect 116648 -24739 177360 -24695
rect 88393 -24770 177360 -24739
rect -75255 -24795 177360 -24770
rect -75255 -24810 109104 -24795
rect -109116 -24826 109104 -24810
rect -109116 -24866 80849 -24826
rect -109116 -24910 -82799 -24866
rect -82755 -24910 -82699 -24866
rect -82655 -24910 -82599 -24866
rect -82555 -24910 -82499 -24866
rect -82455 -24910 -82399 -24866
rect -82355 -24910 -82299 -24866
rect -82255 -24910 -82199 -24866
rect -82155 -24910 -82099 -24866
rect -82055 -24910 -81999 -24866
rect -81955 -24910 -81899 -24866
rect -81855 -24910 -81799 -24866
rect -81755 -24910 -81699 -24866
rect -81655 -24910 -81599 -24866
rect -81555 -24910 -81499 -24866
rect -81455 -24910 -81399 -24866
rect -81355 -24910 -81299 -24866
rect -81255 -24910 -80799 -24866
rect -80755 -24910 -80699 -24866
rect -80655 -24910 -80599 -24866
rect -80555 -24910 -80499 -24866
rect -80455 -24910 -80399 -24866
rect -80355 -24910 -80299 -24866
rect -80255 -24910 -80199 -24866
rect -80155 -24910 -80099 -24866
rect -80055 -24910 -79999 -24866
rect -79955 -24910 -79899 -24866
rect -79855 -24910 -79799 -24866
rect -79755 -24910 -79699 -24866
rect -79655 -24910 -79599 -24866
rect -79555 -24910 -79499 -24866
rect -79455 -24910 -79399 -24866
rect -79355 -24910 -79299 -24866
rect -79255 -24910 -78799 -24866
rect -78755 -24910 -78699 -24866
rect -78655 -24910 -78599 -24866
rect -78555 -24910 -78499 -24866
rect -78455 -24910 -78399 -24866
rect -78355 -24910 -78299 -24866
rect -78255 -24910 -78199 -24866
rect -78155 -24910 -78099 -24866
rect -78055 -24910 -77999 -24866
rect -77955 -24910 -77899 -24866
rect -77855 -24910 -77799 -24866
rect -77755 -24910 -77699 -24866
rect -77655 -24910 -77599 -24866
rect -77555 -24910 -77499 -24866
rect -77455 -24910 -77399 -24866
rect -77355 -24910 -77299 -24866
rect -77255 -24910 -76799 -24866
rect -76755 -24910 -76699 -24866
rect -76655 -24910 -76599 -24866
rect -76555 -24910 -76499 -24866
rect -76455 -24910 -76399 -24866
rect -76355 -24910 -76299 -24866
rect -76255 -24910 -76199 -24866
rect -76155 -24910 -76099 -24866
rect -76055 -24910 -75999 -24866
rect -75955 -24910 -75899 -24866
rect -75855 -24910 -75799 -24866
rect -75755 -24910 -75699 -24866
rect -75655 -24910 -75599 -24866
rect -75555 -24910 -75499 -24866
rect -75455 -24910 -75399 -24866
rect -75355 -24910 -75299 -24866
rect -75255 -24870 80849 -24866
rect 80893 -24870 80949 -24826
rect 80993 -24870 81049 -24826
rect 81093 -24870 81149 -24826
rect 81193 -24870 81249 -24826
rect 81293 -24870 81349 -24826
rect 81393 -24870 81449 -24826
rect 81493 -24870 81549 -24826
rect 81593 -24870 81649 -24826
rect 81693 -24870 81749 -24826
rect 81793 -24870 81849 -24826
rect 81893 -24870 81949 -24826
rect 81993 -24870 82049 -24826
rect 82093 -24870 82149 -24826
rect 82193 -24870 82249 -24826
rect 82293 -24870 82349 -24826
rect 82393 -24870 82849 -24826
rect 82893 -24870 82949 -24826
rect 82993 -24870 83049 -24826
rect 83093 -24870 83149 -24826
rect 83193 -24870 83249 -24826
rect 83293 -24870 83349 -24826
rect 83393 -24870 83449 -24826
rect 83493 -24870 83549 -24826
rect 83593 -24870 83649 -24826
rect 83693 -24870 83749 -24826
rect 83793 -24870 83849 -24826
rect 83893 -24870 83949 -24826
rect 83993 -24870 84049 -24826
rect 84093 -24870 84149 -24826
rect 84193 -24870 84249 -24826
rect 84293 -24870 84349 -24826
rect 84393 -24870 84849 -24826
rect 84893 -24870 84949 -24826
rect 84993 -24870 85049 -24826
rect 85093 -24870 85149 -24826
rect 85193 -24870 85249 -24826
rect 85293 -24870 85349 -24826
rect 85393 -24870 85449 -24826
rect 85493 -24870 85549 -24826
rect 85593 -24870 85649 -24826
rect 85693 -24870 85749 -24826
rect 85793 -24870 85849 -24826
rect 85893 -24870 85949 -24826
rect 85993 -24870 86049 -24826
rect 86093 -24870 86149 -24826
rect 86193 -24870 86249 -24826
rect 86293 -24870 86349 -24826
rect 86393 -24870 86849 -24826
rect 86893 -24870 86949 -24826
rect 86993 -24870 87049 -24826
rect 87093 -24870 87149 -24826
rect 87193 -24870 87249 -24826
rect 87293 -24870 87349 -24826
rect 87393 -24870 87449 -24826
rect 87493 -24870 87549 -24826
rect 87593 -24870 87649 -24826
rect 87693 -24870 87749 -24826
rect 87793 -24870 87849 -24826
rect 87893 -24870 87949 -24826
rect 87993 -24870 88049 -24826
rect 88093 -24870 88149 -24826
rect 88193 -24870 88249 -24826
rect 88293 -24870 88349 -24826
rect 88393 -24839 109104 -24826
rect 109148 -24839 109204 -24795
rect 109248 -24839 109304 -24795
rect 109348 -24839 109404 -24795
rect 109448 -24839 109504 -24795
rect 109548 -24839 109604 -24795
rect 109648 -24839 109704 -24795
rect 109748 -24839 109804 -24795
rect 109848 -24839 109904 -24795
rect 109948 -24839 110004 -24795
rect 110048 -24839 110104 -24795
rect 110148 -24839 110204 -24795
rect 110248 -24839 110304 -24795
rect 110348 -24839 110404 -24795
rect 110448 -24839 110504 -24795
rect 110548 -24839 110604 -24795
rect 110648 -24839 111104 -24795
rect 111148 -24839 111204 -24795
rect 111248 -24839 111304 -24795
rect 111348 -24839 111404 -24795
rect 111448 -24839 111504 -24795
rect 111548 -24839 111604 -24795
rect 111648 -24839 111704 -24795
rect 111748 -24839 111804 -24795
rect 111848 -24839 111904 -24795
rect 111948 -24839 112004 -24795
rect 112048 -24839 112104 -24795
rect 112148 -24839 112204 -24795
rect 112248 -24839 112304 -24795
rect 112348 -24839 112404 -24795
rect 112448 -24839 112504 -24795
rect 112548 -24839 112604 -24795
rect 112648 -24839 113104 -24795
rect 113148 -24839 113204 -24795
rect 113248 -24839 113304 -24795
rect 113348 -24839 113404 -24795
rect 113448 -24839 113504 -24795
rect 113548 -24839 113604 -24795
rect 113648 -24839 113704 -24795
rect 113748 -24839 113804 -24795
rect 113848 -24839 113904 -24795
rect 113948 -24839 114004 -24795
rect 114048 -24839 114104 -24795
rect 114148 -24839 114204 -24795
rect 114248 -24839 114304 -24795
rect 114348 -24839 114404 -24795
rect 114448 -24839 114504 -24795
rect 114548 -24839 114604 -24795
rect 114648 -24839 115104 -24795
rect 115148 -24839 115204 -24795
rect 115248 -24839 115304 -24795
rect 115348 -24839 115404 -24795
rect 115448 -24839 115504 -24795
rect 115548 -24839 115604 -24795
rect 115648 -24839 115704 -24795
rect 115748 -24839 115804 -24795
rect 115848 -24839 115904 -24795
rect 115948 -24839 116004 -24795
rect 116048 -24839 116104 -24795
rect 116148 -24839 116204 -24795
rect 116248 -24839 116304 -24795
rect 116348 -24839 116404 -24795
rect 116448 -24839 116504 -24795
rect 116548 -24839 116604 -24795
rect 116648 -24839 177360 -24795
rect 88393 -24870 177360 -24839
rect -75255 -24895 177360 -24870
rect -75255 -24910 109104 -24895
rect -109116 -24926 109104 -24910
rect -109116 -24966 80849 -24926
rect -109116 -25010 -82799 -24966
rect -82755 -25010 -82699 -24966
rect -82655 -25010 -82599 -24966
rect -82555 -25010 -82499 -24966
rect -82455 -25010 -82399 -24966
rect -82355 -25010 -82299 -24966
rect -82255 -25010 -82199 -24966
rect -82155 -25010 -82099 -24966
rect -82055 -25010 -81999 -24966
rect -81955 -25010 -81899 -24966
rect -81855 -25010 -81799 -24966
rect -81755 -25010 -81699 -24966
rect -81655 -25010 -81599 -24966
rect -81555 -25010 -81499 -24966
rect -81455 -25010 -81399 -24966
rect -81355 -25010 -81299 -24966
rect -81255 -25010 -80799 -24966
rect -80755 -25010 -80699 -24966
rect -80655 -25010 -80599 -24966
rect -80555 -25010 -80499 -24966
rect -80455 -25010 -80399 -24966
rect -80355 -25010 -80299 -24966
rect -80255 -25010 -80199 -24966
rect -80155 -25010 -80099 -24966
rect -80055 -25010 -79999 -24966
rect -79955 -25010 -79899 -24966
rect -79855 -25010 -79799 -24966
rect -79755 -25010 -79699 -24966
rect -79655 -25010 -79599 -24966
rect -79555 -25010 -79499 -24966
rect -79455 -25010 -79399 -24966
rect -79355 -25010 -79299 -24966
rect -79255 -25010 -78799 -24966
rect -78755 -25010 -78699 -24966
rect -78655 -25010 -78599 -24966
rect -78555 -25010 -78499 -24966
rect -78455 -25010 -78399 -24966
rect -78355 -25010 -78299 -24966
rect -78255 -25010 -78199 -24966
rect -78155 -25010 -78099 -24966
rect -78055 -25010 -77999 -24966
rect -77955 -25010 -77899 -24966
rect -77855 -25010 -77799 -24966
rect -77755 -25010 -77699 -24966
rect -77655 -25010 -77599 -24966
rect -77555 -25010 -77499 -24966
rect -77455 -25010 -77399 -24966
rect -77355 -25010 -77299 -24966
rect -77255 -25010 -76799 -24966
rect -76755 -25010 -76699 -24966
rect -76655 -25010 -76599 -24966
rect -76555 -25010 -76499 -24966
rect -76455 -25010 -76399 -24966
rect -76355 -25010 -76299 -24966
rect -76255 -25010 -76199 -24966
rect -76155 -25010 -76099 -24966
rect -76055 -25010 -75999 -24966
rect -75955 -25010 -75899 -24966
rect -75855 -25010 -75799 -24966
rect -75755 -25010 -75699 -24966
rect -75655 -25010 -75599 -24966
rect -75555 -25010 -75499 -24966
rect -75455 -25010 -75399 -24966
rect -75355 -25010 -75299 -24966
rect -75255 -24970 80849 -24966
rect 80893 -24970 80949 -24926
rect 80993 -24970 81049 -24926
rect 81093 -24970 81149 -24926
rect 81193 -24970 81249 -24926
rect 81293 -24970 81349 -24926
rect 81393 -24970 81449 -24926
rect 81493 -24970 81549 -24926
rect 81593 -24970 81649 -24926
rect 81693 -24970 81749 -24926
rect 81793 -24970 81849 -24926
rect 81893 -24970 81949 -24926
rect 81993 -24970 82049 -24926
rect 82093 -24970 82149 -24926
rect 82193 -24970 82249 -24926
rect 82293 -24970 82349 -24926
rect 82393 -24970 82849 -24926
rect 82893 -24970 82949 -24926
rect 82993 -24970 83049 -24926
rect 83093 -24970 83149 -24926
rect 83193 -24970 83249 -24926
rect 83293 -24970 83349 -24926
rect 83393 -24970 83449 -24926
rect 83493 -24970 83549 -24926
rect 83593 -24970 83649 -24926
rect 83693 -24970 83749 -24926
rect 83793 -24970 83849 -24926
rect 83893 -24970 83949 -24926
rect 83993 -24970 84049 -24926
rect 84093 -24970 84149 -24926
rect 84193 -24970 84249 -24926
rect 84293 -24970 84349 -24926
rect 84393 -24970 84849 -24926
rect 84893 -24970 84949 -24926
rect 84993 -24970 85049 -24926
rect 85093 -24970 85149 -24926
rect 85193 -24970 85249 -24926
rect 85293 -24970 85349 -24926
rect 85393 -24970 85449 -24926
rect 85493 -24970 85549 -24926
rect 85593 -24970 85649 -24926
rect 85693 -24970 85749 -24926
rect 85793 -24970 85849 -24926
rect 85893 -24970 85949 -24926
rect 85993 -24970 86049 -24926
rect 86093 -24970 86149 -24926
rect 86193 -24970 86249 -24926
rect 86293 -24970 86349 -24926
rect 86393 -24970 86849 -24926
rect 86893 -24970 86949 -24926
rect 86993 -24970 87049 -24926
rect 87093 -24970 87149 -24926
rect 87193 -24970 87249 -24926
rect 87293 -24970 87349 -24926
rect 87393 -24970 87449 -24926
rect 87493 -24970 87549 -24926
rect 87593 -24970 87649 -24926
rect 87693 -24970 87749 -24926
rect 87793 -24970 87849 -24926
rect 87893 -24970 87949 -24926
rect 87993 -24970 88049 -24926
rect 88093 -24970 88149 -24926
rect 88193 -24970 88249 -24926
rect 88293 -24970 88349 -24926
rect 88393 -24939 109104 -24926
rect 109148 -24939 109204 -24895
rect 109248 -24939 109304 -24895
rect 109348 -24939 109404 -24895
rect 109448 -24939 109504 -24895
rect 109548 -24939 109604 -24895
rect 109648 -24939 109704 -24895
rect 109748 -24939 109804 -24895
rect 109848 -24939 109904 -24895
rect 109948 -24939 110004 -24895
rect 110048 -24939 110104 -24895
rect 110148 -24939 110204 -24895
rect 110248 -24939 110304 -24895
rect 110348 -24939 110404 -24895
rect 110448 -24939 110504 -24895
rect 110548 -24939 110604 -24895
rect 110648 -24939 111104 -24895
rect 111148 -24939 111204 -24895
rect 111248 -24939 111304 -24895
rect 111348 -24939 111404 -24895
rect 111448 -24939 111504 -24895
rect 111548 -24939 111604 -24895
rect 111648 -24939 111704 -24895
rect 111748 -24939 111804 -24895
rect 111848 -24939 111904 -24895
rect 111948 -24939 112004 -24895
rect 112048 -24939 112104 -24895
rect 112148 -24939 112204 -24895
rect 112248 -24939 112304 -24895
rect 112348 -24939 112404 -24895
rect 112448 -24939 112504 -24895
rect 112548 -24939 112604 -24895
rect 112648 -24939 113104 -24895
rect 113148 -24939 113204 -24895
rect 113248 -24939 113304 -24895
rect 113348 -24939 113404 -24895
rect 113448 -24939 113504 -24895
rect 113548 -24939 113604 -24895
rect 113648 -24939 113704 -24895
rect 113748 -24939 113804 -24895
rect 113848 -24939 113904 -24895
rect 113948 -24939 114004 -24895
rect 114048 -24939 114104 -24895
rect 114148 -24939 114204 -24895
rect 114248 -24939 114304 -24895
rect 114348 -24939 114404 -24895
rect 114448 -24939 114504 -24895
rect 114548 -24939 114604 -24895
rect 114648 -24939 115104 -24895
rect 115148 -24939 115204 -24895
rect 115248 -24939 115304 -24895
rect 115348 -24939 115404 -24895
rect 115448 -24939 115504 -24895
rect 115548 -24939 115604 -24895
rect 115648 -24939 115704 -24895
rect 115748 -24939 115804 -24895
rect 115848 -24939 115904 -24895
rect 115948 -24939 116004 -24895
rect 116048 -24939 116104 -24895
rect 116148 -24939 116204 -24895
rect 116248 -24939 116304 -24895
rect 116348 -24939 116404 -24895
rect 116448 -24939 116504 -24895
rect 116548 -24939 116604 -24895
rect 116648 -24939 177360 -24895
rect 88393 -24970 177360 -24939
rect -75255 -24995 177360 -24970
rect -75255 -25010 109104 -24995
rect -109116 -25026 109104 -25010
rect -109116 -25066 80849 -25026
rect -109116 -25110 -82799 -25066
rect -82755 -25110 -82699 -25066
rect -82655 -25110 -82599 -25066
rect -82555 -25110 -82499 -25066
rect -82455 -25110 -82399 -25066
rect -82355 -25110 -82299 -25066
rect -82255 -25110 -82199 -25066
rect -82155 -25110 -82099 -25066
rect -82055 -25110 -81999 -25066
rect -81955 -25110 -81899 -25066
rect -81855 -25110 -81799 -25066
rect -81755 -25110 -81699 -25066
rect -81655 -25110 -81599 -25066
rect -81555 -25110 -81499 -25066
rect -81455 -25110 -81399 -25066
rect -81355 -25110 -81299 -25066
rect -81255 -25110 -80799 -25066
rect -80755 -25110 -80699 -25066
rect -80655 -25110 -80599 -25066
rect -80555 -25110 -80499 -25066
rect -80455 -25110 -80399 -25066
rect -80355 -25110 -80299 -25066
rect -80255 -25110 -80199 -25066
rect -80155 -25110 -80099 -25066
rect -80055 -25110 -79999 -25066
rect -79955 -25110 -79899 -25066
rect -79855 -25110 -79799 -25066
rect -79755 -25110 -79699 -25066
rect -79655 -25110 -79599 -25066
rect -79555 -25110 -79499 -25066
rect -79455 -25110 -79399 -25066
rect -79355 -25110 -79299 -25066
rect -79255 -25110 -78799 -25066
rect -78755 -25110 -78699 -25066
rect -78655 -25110 -78599 -25066
rect -78555 -25110 -78499 -25066
rect -78455 -25110 -78399 -25066
rect -78355 -25110 -78299 -25066
rect -78255 -25110 -78199 -25066
rect -78155 -25110 -78099 -25066
rect -78055 -25110 -77999 -25066
rect -77955 -25110 -77899 -25066
rect -77855 -25110 -77799 -25066
rect -77755 -25110 -77699 -25066
rect -77655 -25110 -77599 -25066
rect -77555 -25110 -77499 -25066
rect -77455 -25110 -77399 -25066
rect -77355 -25110 -77299 -25066
rect -77255 -25110 -76799 -25066
rect -76755 -25110 -76699 -25066
rect -76655 -25110 -76599 -25066
rect -76555 -25110 -76499 -25066
rect -76455 -25110 -76399 -25066
rect -76355 -25110 -76299 -25066
rect -76255 -25110 -76199 -25066
rect -76155 -25110 -76099 -25066
rect -76055 -25110 -75999 -25066
rect -75955 -25110 -75899 -25066
rect -75855 -25110 -75799 -25066
rect -75755 -25110 -75699 -25066
rect -75655 -25110 -75599 -25066
rect -75555 -25110 -75499 -25066
rect -75455 -25110 -75399 -25066
rect -75355 -25110 -75299 -25066
rect -75255 -25070 80849 -25066
rect 80893 -25070 80949 -25026
rect 80993 -25070 81049 -25026
rect 81093 -25070 81149 -25026
rect 81193 -25070 81249 -25026
rect 81293 -25070 81349 -25026
rect 81393 -25070 81449 -25026
rect 81493 -25070 81549 -25026
rect 81593 -25070 81649 -25026
rect 81693 -25070 81749 -25026
rect 81793 -25070 81849 -25026
rect 81893 -25070 81949 -25026
rect 81993 -25070 82049 -25026
rect 82093 -25070 82149 -25026
rect 82193 -25070 82249 -25026
rect 82293 -25070 82349 -25026
rect 82393 -25070 82849 -25026
rect 82893 -25070 82949 -25026
rect 82993 -25070 83049 -25026
rect 83093 -25070 83149 -25026
rect 83193 -25070 83249 -25026
rect 83293 -25070 83349 -25026
rect 83393 -25070 83449 -25026
rect 83493 -25070 83549 -25026
rect 83593 -25070 83649 -25026
rect 83693 -25070 83749 -25026
rect 83793 -25070 83849 -25026
rect 83893 -25070 83949 -25026
rect 83993 -25070 84049 -25026
rect 84093 -25070 84149 -25026
rect 84193 -25070 84249 -25026
rect 84293 -25070 84349 -25026
rect 84393 -25070 84849 -25026
rect 84893 -25070 84949 -25026
rect 84993 -25070 85049 -25026
rect 85093 -25070 85149 -25026
rect 85193 -25070 85249 -25026
rect 85293 -25070 85349 -25026
rect 85393 -25070 85449 -25026
rect 85493 -25070 85549 -25026
rect 85593 -25070 85649 -25026
rect 85693 -25070 85749 -25026
rect 85793 -25070 85849 -25026
rect 85893 -25070 85949 -25026
rect 85993 -25070 86049 -25026
rect 86093 -25070 86149 -25026
rect 86193 -25070 86249 -25026
rect 86293 -25070 86349 -25026
rect 86393 -25070 86849 -25026
rect 86893 -25070 86949 -25026
rect 86993 -25070 87049 -25026
rect 87093 -25070 87149 -25026
rect 87193 -25070 87249 -25026
rect 87293 -25070 87349 -25026
rect 87393 -25070 87449 -25026
rect 87493 -25070 87549 -25026
rect 87593 -25070 87649 -25026
rect 87693 -25070 87749 -25026
rect 87793 -25070 87849 -25026
rect 87893 -25070 87949 -25026
rect 87993 -25070 88049 -25026
rect 88093 -25070 88149 -25026
rect 88193 -25070 88249 -25026
rect 88293 -25070 88349 -25026
rect 88393 -25039 109104 -25026
rect 109148 -25039 109204 -24995
rect 109248 -25039 109304 -24995
rect 109348 -25039 109404 -24995
rect 109448 -25039 109504 -24995
rect 109548 -25039 109604 -24995
rect 109648 -25039 109704 -24995
rect 109748 -25039 109804 -24995
rect 109848 -25039 109904 -24995
rect 109948 -25039 110004 -24995
rect 110048 -25039 110104 -24995
rect 110148 -25039 110204 -24995
rect 110248 -25039 110304 -24995
rect 110348 -25039 110404 -24995
rect 110448 -25039 110504 -24995
rect 110548 -25039 110604 -24995
rect 110648 -25039 111104 -24995
rect 111148 -25039 111204 -24995
rect 111248 -25039 111304 -24995
rect 111348 -25039 111404 -24995
rect 111448 -25039 111504 -24995
rect 111548 -25039 111604 -24995
rect 111648 -25039 111704 -24995
rect 111748 -25039 111804 -24995
rect 111848 -25039 111904 -24995
rect 111948 -25039 112004 -24995
rect 112048 -25039 112104 -24995
rect 112148 -25039 112204 -24995
rect 112248 -25039 112304 -24995
rect 112348 -25039 112404 -24995
rect 112448 -25039 112504 -24995
rect 112548 -25039 112604 -24995
rect 112648 -25039 113104 -24995
rect 113148 -25039 113204 -24995
rect 113248 -25039 113304 -24995
rect 113348 -25039 113404 -24995
rect 113448 -25039 113504 -24995
rect 113548 -25039 113604 -24995
rect 113648 -25039 113704 -24995
rect 113748 -25039 113804 -24995
rect 113848 -25039 113904 -24995
rect 113948 -25039 114004 -24995
rect 114048 -25039 114104 -24995
rect 114148 -25039 114204 -24995
rect 114248 -25039 114304 -24995
rect 114348 -25039 114404 -24995
rect 114448 -25039 114504 -24995
rect 114548 -25039 114604 -24995
rect 114648 -25039 115104 -24995
rect 115148 -25039 115204 -24995
rect 115248 -25039 115304 -24995
rect 115348 -25039 115404 -24995
rect 115448 -25039 115504 -24995
rect 115548 -25039 115604 -24995
rect 115648 -25039 115704 -24995
rect 115748 -25039 115804 -24995
rect 115848 -25039 115904 -24995
rect 115948 -25039 116004 -24995
rect 116048 -25039 116104 -24995
rect 116148 -25039 116204 -24995
rect 116248 -25039 116304 -24995
rect 116348 -25039 116404 -24995
rect 116448 -25039 116504 -24995
rect 116548 -25039 116604 -24995
rect 116648 -25039 177360 -24995
rect 88393 -25070 177360 -25039
rect -75255 -25095 177360 -25070
rect -75255 -25110 109104 -25095
rect -109116 -25126 109104 -25110
rect -109116 -25166 80849 -25126
rect -109116 -25210 -82799 -25166
rect -82755 -25210 -82699 -25166
rect -82655 -25210 -82599 -25166
rect -82555 -25210 -82499 -25166
rect -82455 -25210 -82399 -25166
rect -82355 -25210 -82299 -25166
rect -82255 -25210 -82199 -25166
rect -82155 -25210 -82099 -25166
rect -82055 -25210 -81999 -25166
rect -81955 -25210 -81899 -25166
rect -81855 -25210 -81799 -25166
rect -81755 -25210 -81699 -25166
rect -81655 -25210 -81599 -25166
rect -81555 -25210 -81499 -25166
rect -81455 -25210 -81399 -25166
rect -81355 -25210 -81299 -25166
rect -81255 -25210 -80799 -25166
rect -80755 -25210 -80699 -25166
rect -80655 -25210 -80599 -25166
rect -80555 -25210 -80499 -25166
rect -80455 -25210 -80399 -25166
rect -80355 -25210 -80299 -25166
rect -80255 -25210 -80199 -25166
rect -80155 -25210 -80099 -25166
rect -80055 -25210 -79999 -25166
rect -79955 -25210 -79899 -25166
rect -79855 -25210 -79799 -25166
rect -79755 -25210 -79699 -25166
rect -79655 -25210 -79599 -25166
rect -79555 -25210 -79499 -25166
rect -79455 -25210 -79399 -25166
rect -79355 -25210 -79299 -25166
rect -79255 -25210 -78799 -25166
rect -78755 -25210 -78699 -25166
rect -78655 -25210 -78599 -25166
rect -78555 -25210 -78499 -25166
rect -78455 -25210 -78399 -25166
rect -78355 -25210 -78299 -25166
rect -78255 -25210 -78199 -25166
rect -78155 -25210 -78099 -25166
rect -78055 -25210 -77999 -25166
rect -77955 -25210 -77899 -25166
rect -77855 -25210 -77799 -25166
rect -77755 -25210 -77699 -25166
rect -77655 -25210 -77599 -25166
rect -77555 -25210 -77499 -25166
rect -77455 -25210 -77399 -25166
rect -77355 -25210 -77299 -25166
rect -77255 -25210 -76799 -25166
rect -76755 -25210 -76699 -25166
rect -76655 -25210 -76599 -25166
rect -76555 -25210 -76499 -25166
rect -76455 -25210 -76399 -25166
rect -76355 -25210 -76299 -25166
rect -76255 -25210 -76199 -25166
rect -76155 -25210 -76099 -25166
rect -76055 -25210 -75999 -25166
rect -75955 -25210 -75899 -25166
rect -75855 -25210 -75799 -25166
rect -75755 -25210 -75699 -25166
rect -75655 -25210 -75599 -25166
rect -75555 -25210 -75499 -25166
rect -75455 -25210 -75399 -25166
rect -75355 -25210 -75299 -25166
rect -75255 -25170 80849 -25166
rect 80893 -25170 80949 -25126
rect 80993 -25170 81049 -25126
rect 81093 -25170 81149 -25126
rect 81193 -25170 81249 -25126
rect 81293 -25170 81349 -25126
rect 81393 -25170 81449 -25126
rect 81493 -25170 81549 -25126
rect 81593 -25170 81649 -25126
rect 81693 -25170 81749 -25126
rect 81793 -25170 81849 -25126
rect 81893 -25170 81949 -25126
rect 81993 -25170 82049 -25126
rect 82093 -25170 82149 -25126
rect 82193 -25170 82249 -25126
rect 82293 -25170 82349 -25126
rect 82393 -25170 82849 -25126
rect 82893 -25170 82949 -25126
rect 82993 -25170 83049 -25126
rect 83093 -25170 83149 -25126
rect 83193 -25170 83249 -25126
rect 83293 -25170 83349 -25126
rect 83393 -25170 83449 -25126
rect 83493 -25170 83549 -25126
rect 83593 -25170 83649 -25126
rect 83693 -25170 83749 -25126
rect 83793 -25170 83849 -25126
rect 83893 -25170 83949 -25126
rect 83993 -25170 84049 -25126
rect 84093 -25170 84149 -25126
rect 84193 -25170 84249 -25126
rect 84293 -25170 84349 -25126
rect 84393 -25170 84849 -25126
rect 84893 -25170 84949 -25126
rect 84993 -25170 85049 -25126
rect 85093 -25170 85149 -25126
rect 85193 -25170 85249 -25126
rect 85293 -25170 85349 -25126
rect 85393 -25170 85449 -25126
rect 85493 -25170 85549 -25126
rect 85593 -25170 85649 -25126
rect 85693 -25170 85749 -25126
rect 85793 -25170 85849 -25126
rect 85893 -25170 85949 -25126
rect 85993 -25170 86049 -25126
rect 86093 -25170 86149 -25126
rect 86193 -25170 86249 -25126
rect 86293 -25170 86349 -25126
rect 86393 -25170 86849 -25126
rect 86893 -25170 86949 -25126
rect 86993 -25170 87049 -25126
rect 87093 -25170 87149 -25126
rect 87193 -25170 87249 -25126
rect 87293 -25170 87349 -25126
rect 87393 -25170 87449 -25126
rect 87493 -25170 87549 -25126
rect 87593 -25170 87649 -25126
rect 87693 -25170 87749 -25126
rect 87793 -25170 87849 -25126
rect 87893 -25170 87949 -25126
rect 87993 -25170 88049 -25126
rect 88093 -25170 88149 -25126
rect 88193 -25170 88249 -25126
rect 88293 -25170 88349 -25126
rect 88393 -25139 109104 -25126
rect 109148 -25139 109204 -25095
rect 109248 -25139 109304 -25095
rect 109348 -25139 109404 -25095
rect 109448 -25139 109504 -25095
rect 109548 -25139 109604 -25095
rect 109648 -25139 109704 -25095
rect 109748 -25139 109804 -25095
rect 109848 -25139 109904 -25095
rect 109948 -25139 110004 -25095
rect 110048 -25139 110104 -25095
rect 110148 -25139 110204 -25095
rect 110248 -25139 110304 -25095
rect 110348 -25139 110404 -25095
rect 110448 -25139 110504 -25095
rect 110548 -25139 110604 -25095
rect 110648 -25139 111104 -25095
rect 111148 -25139 111204 -25095
rect 111248 -25139 111304 -25095
rect 111348 -25139 111404 -25095
rect 111448 -25139 111504 -25095
rect 111548 -25139 111604 -25095
rect 111648 -25139 111704 -25095
rect 111748 -25139 111804 -25095
rect 111848 -25139 111904 -25095
rect 111948 -25139 112004 -25095
rect 112048 -25139 112104 -25095
rect 112148 -25139 112204 -25095
rect 112248 -25139 112304 -25095
rect 112348 -25139 112404 -25095
rect 112448 -25139 112504 -25095
rect 112548 -25139 112604 -25095
rect 112648 -25139 113104 -25095
rect 113148 -25139 113204 -25095
rect 113248 -25139 113304 -25095
rect 113348 -25139 113404 -25095
rect 113448 -25139 113504 -25095
rect 113548 -25139 113604 -25095
rect 113648 -25139 113704 -25095
rect 113748 -25139 113804 -25095
rect 113848 -25139 113904 -25095
rect 113948 -25139 114004 -25095
rect 114048 -25139 114104 -25095
rect 114148 -25139 114204 -25095
rect 114248 -25139 114304 -25095
rect 114348 -25139 114404 -25095
rect 114448 -25139 114504 -25095
rect 114548 -25139 114604 -25095
rect 114648 -25139 115104 -25095
rect 115148 -25139 115204 -25095
rect 115248 -25139 115304 -25095
rect 115348 -25139 115404 -25095
rect 115448 -25139 115504 -25095
rect 115548 -25139 115604 -25095
rect 115648 -25139 115704 -25095
rect 115748 -25139 115804 -25095
rect 115848 -25139 115904 -25095
rect 115948 -25139 116004 -25095
rect 116048 -25139 116104 -25095
rect 116148 -25139 116204 -25095
rect 116248 -25139 116304 -25095
rect 116348 -25139 116404 -25095
rect 116448 -25139 116504 -25095
rect 116548 -25139 116604 -25095
rect 116648 -25139 177360 -25095
rect 88393 -25170 177360 -25139
rect -75255 -25195 177360 -25170
rect -75255 -25210 109104 -25195
rect -109116 -25226 109104 -25210
rect -109116 -25266 80849 -25226
rect -109116 -25310 -82799 -25266
rect -82755 -25310 -82699 -25266
rect -82655 -25310 -82599 -25266
rect -82555 -25310 -82499 -25266
rect -82455 -25310 -82399 -25266
rect -82355 -25310 -82299 -25266
rect -82255 -25310 -82199 -25266
rect -82155 -25310 -82099 -25266
rect -82055 -25310 -81999 -25266
rect -81955 -25310 -81899 -25266
rect -81855 -25310 -81799 -25266
rect -81755 -25310 -81699 -25266
rect -81655 -25310 -81599 -25266
rect -81555 -25310 -81499 -25266
rect -81455 -25310 -81399 -25266
rect -81355 -25310 -81299 -25266
rect -81255 -25310 -80799 -25266
rect -80755 -25310 -80699 -25266
rect -80655 -25310 -80599 -25266
rect -80555 -25310 -80499 -25266
rect -80455 -25310 -80399 -25266
rect -80355 -25310 -80299 -25266
rect -80255 -25310 -80199 -25266
rect -80155 -25310 -80099 -25266
rect -80055 -25310 -79999 -25266
rect -79955 -25310 -79899 -25266
rect -79855 -25310 -79799 -25266
rect -79755 -25310 -79699 -25266
rect -79655 -25310 -79599 -25266
rect -79555 -25310 -79499 -25266
rect -79455 -25310 -79399 -25266
rect -79355 -25310 -79299 -25266
rect -79255 -25310 -78799 -25266
rect -78755 -25310 -78699 -25266
rect -78655 -25310 -78599 -25266
rect -78555 -25310 -78499 -25266
rect -78455 -25310 -78399 -25266
rect -78355 -25310 -78299 -25266
rect -78255 -25310 -78199 -25266
rect -78155 -25310 -78099 -25266
rect -78055 -25310 -77999 -25266
rect -77955 -25310 -77899 -25266
rect -77855 -25310 -77799 -25266
rect -77755 -25310 -77699 -25266
rect -77655 -25310 -77599 -25266
rect -77555 -25310 -77499 -25266
rect -77455 -25310 -77399 -25266
rect -77355 -25310 -77299 -25266
rect -77255 -25310 -76799 -25266
rect -76755 -25310 -76699 -25266
rect -76655 -25310 -76599 -25266
rect -76555 -25310 -76499 -25266
rect -76455 -25310 -76399 -25266
rect -76355 -25310 -76299 -25266
rect -76255 -25310 -76199 -25266
rect -76155 -25310 -76099 -25266
rect -76055 -25310 -75999 -25266
rect -75955 -25310 -75899 -25266
rect -75855 -25310 -75799 -25266
rect -75755 -25310 -75699 -25266
rect -75655 -25310 -75599 -25266
rect -75555 -25310 -75499 -25266
rect -75455 -25310 -75399 -25266
rect -75355 -25310 -75299 -25266
rect -75255 -25270 80849 -25266
rect 80893 -25270 80949 -25226
rect 80993 -25270 81049 -25226
rect 81093 -25270 81149 -25226
rect 81193 -25270 81249 -25226
rect 81293 -25270 81349 -25226
rect 81393 -25270 81449 -25226
rect 81493 -25270 81549 -25226
rect 81593 -25270 81649 -25226
rect 81693 -25270 81749 -25226
rect 81793 -25270 81849 -25226
rect 81893 -25270 81949 -25226
rect 81993 -25270 82049 -25226
rect 82093 -25270 82149 -25226
rect 82193 -25270 82249 -25226
rect 82293 -25270 82349 -25226
rect 82393 -25270 82849 -25226
rect 82893 -25270 82949 -25226
rect 82993 -25270 83049 -25226
rect 83093 -25270 83149 -25226
rect 83193 -25270 83249 -25226
rect 83293 -25270 83349 -25226
rect 83393 -25270 83449 -25226
rect 83493 -25270 83549 -25226
rect 83593 -25270 83649 -25226
rect 83693 -25270 83749 -25226
rect 83793 -25270 83849 -25226
rect 83893 -25270 83949 -25226
rect 83993 -25270 84049 -25226
rect 84093 -25270 84149 -25226
rect 84193 -25270 84249 -25226
rect 84293 -25270 84349 -25226
rect 84393 -25270 84849 -25226
rect 84893 -25270 84949 -25226
rect 84993 -25270 85049 -25226
rect 85093 -25270 85149 -25226
rect 85193 -25270 85249 -25226
rect 85293 -25270 85349 -25226
rect 85393 -25270 85449 -25226
rect 85493 -25270 85549 -25226
rect 85593 -25270 85649 -25226
rect 85693 -25270 85749 -25226
rect 85793 -25270 85849 -25226
rect 85893 -25270 85949 -25226
rect 85993 -25270 86049 -25226
rect 86093 -25270 86149 -25226
rect 86193 -25270 86249 -25226
rect 86293 -25270 86349 -25226
rect 86393 -25270 86849 -25226
rect 86893 -25270 86949 -25226
rect 86993 -25270 87049 -25226
rect 87093 -25270 87149 -25226
rect 87193 -25270 87249 -25226
rect 87293 -25270 87349 -25226
rect 87393 -25270 87449 -25226
rect 87493 -25270 87549 -25226
rect 87593 -25270 87649 -25226
rect 87693 -25270 87749 -25226
rect 87793 -25270 87849 -25226
rect 87893 -25270 87949 -25226
rect 87993 -25270 88049 -25226
rect 88093 -25270 88149 -25226
rect 88193 -25270 88249 -25226
rect 88293 -25270 88349 -25226
rect 88393 -25239 109104 -25226
rect 109148 -25239 109204 -25195
rect 109248 -25239 109304 -25195
rect 109348 -25239 109404 -25195
rect 109448 -25239 109504 -25195
rect 109548 -25239 109604 -25195
rect 109648 -25239 109704 -25195
rect 109748 -25239 109804 -25195
rect 109848 -25239 109904 -25195
rect 109948 -25239 110004 -25195
rect 110048 -25239 110104 -25195
rect 110148 -25239 110204 -25195
rect 110248 -25239 110304 -25195
rect 110348 -25239 110404 -25195
rect 110448 -25239 110504 -25195
rect 110548 -25239 110604 -25195
rect 110648 -25239 111104 -25195
rect 111148 -25239 111204 -25195
rect 111248 -25239 111304 -25195
rect 111348 -25239 111404 -25195
rect 111448 -25239 111504 -25195
rect 111548 -25239 111604 -25195
rect 111648 -25239 111704 -25195
rect 111748 -25239 111804 -25195
rect 111848 -25239 111904 -25195
rect 111948 -25239 112004 -25195
rect 112048 -25239 112104 -25195
rect 112148 -25239 112204 -25195
rect 112248 -25239 112304 -25195
rect 112348 -25239 112404 -25195
rect 112448 -25239 112504 -25195
rect 112548 -25239 112604 -25195
rect 112648 -25239 113104 -25195
rect 113148 -25239 113204 -25195
rect 113248 -25239 113304 -25195
rect 113348 -25239 113404 -25195
rect 113448 -25239 113504 -25195
rect 113548 -25239 113604 -25195
rect 113648 -25239 113704 -25195
rect 113748 -25239 113804 -25195
rect 113848 -25239 113904 -25195
rect 113948 -25239 114004 -25195
rect 114048 -25239 114104 -25195
rect 114148 -25239 114204 -25195
rect 114248 -25239 114304 -25195
rect 114348 -25239 114404 -25195
rect 114448 -25239 114504 -25195
rect 114548 -25239 114604 -25195
rect 114648 -25239 115104 -25195
rect 115148 -25239 115204 -25195
rect 115248 -25239 115304 -25195
rect 115348 -25239 115404 -25195
rect 115448 -25239 115504 -25195
rect 115548 -25239 115604 -25195
rect 115648 -25239 115704 -25195
rect 115748 -25239 115804 -25195
rect 115848 -25239 115904 -25195
rect 115948 -25239 116004 -25195
rect 116048 -25239 116104 -25195
rect 116148 -25239 116204 -25195
rect 116248 -25239 116304 -25195
rect 116348 -25239 116404 -25195
rect 116448 -25239 116504 -25195
rect 116548 -25239 116604 -25195
rect 116648 -25239 177360 -25195
rect 88393 -25270 177360 -25239
rect -75255 -25295 177360 -25270
rect -75255 -25310 109104 -25295
rect -109116 -25326 109104 -25310
rect -109116 -25366 80849 -25326
rect -109116 -25410 -82799 -25366
rect -82755 -25410 -82699 -25366
rect -82655 -25410 -82599 -25366
rect -82555 -25410 -82499 -25366
rect -82455 -25410 -82399 -25366
rect -82355 -25410 -82299 -25366
rect -82255 -25410 -82199 -25366
rect -82155 -25410 -82099 -25366
rect -82055 -25410 -81999 -25366
rect -81955 -25410 -81899 -25366
rect -81855 -25410 -81799 -25366
rect -81755 -25410 -81699 -25366
rect -81655 -25410 -81599 -25366
rect -81555 -25410 -81499 -25366
rect -81455 -25410 -81399 -25366
rect -81355 -25410 -81299 -25366
rect -81255 -25410 -80799 -25366
rect -80755 -25410 -80699 -25366
rect -80655 -25410 -80599 -25366
rect -80555 -25410 -80499 -25366
rect -80455 -25410 -80399 -25366
rect -80355 -25410 -80299 -25366
rect -80255 -25410 -80199 -25366
rect -80155 -25410 -80099 -25366
rect -80055 -25410 -79999 -25366
rect -79955 -25410 -79899 -25366
rect -79855 -25410 -79799 -25366
rect -79755 -25410 -79699 -25366
rect -79655 -25410 -79599 -25366
rect -79555 -25410 -79499 -25366
rect -79455 -25410 -79399 -25366
rect -79355 -25410 -79299 -25366
rect -79255 -25410 -78799 -25366
rect -78755 -25410 -78699 -25366
rect -78655 -25410 -78599 -25366
rect -78555 -25410 -78499 -25366
rect -78455 -25410 -78399 -25366
rect -78355 -25410 -78299 -25366
rect -78255 -25410 -78199 -25366
rect -78155 -25410 -78099 -25366
rect -78055 -25410 -77999 -25366
rect -77955 -25410 -77899 -25366
rect -77855 -25410 -77799 -25366
rect -77755 -25410 -77699 -25366
rect -77655 -25410 -77599 -25366
rect -77555 -25410 -77499 -25366
rect -77455 -25410 -77399 -25366
rect -77355 -25410 -77299 -25366
rect -77255 -25410 -76799 -25366
rect -76755 -25410 -76699 -25366
rect -76655 -25410 -76599 -25366
rect -76555 -25410 -76499 -25366
rect -76455 -25410 -76399 -25366
rect -76355 -25410 -76299 -25366
rect -76255 -25410 -76199 -25366
rect -76155 -25410 -76099 -25366
rect -76055 -25410 -75999 -25366
rect -75955 -25410 -75899 -25366
rect -75855 -25410 -75799 -25366
rect -75755 -25410 -75699 -25366
rect -75655 -25410 -75599 -25366
rect -75555 -25410 -75499 -25366
rect -75455 -25410 -75399 -25366
rect -75355 -25410 -75299 -25366
rect -75255 -25370 80849 -25366
rect 80893 -25370 80949 -25326
rect 80993 -25370 81049 -25326
rect 81093 -25370 81149 -25326
rect 81193 -25370 81249 -25326
rect 81293 -25370 81349 -25326
rect 81393 -25370 81449 -25326
rect 81493 -25370 81549 -25326
rect 81593 -25370 81649 -25326
rect 81693 -25370 81749 -25326
rect 81793 -25370 81849 -25326
rect 81893 -25370 81949 -25326
rect 81993 -25370 82049 -25326
rect 82093 -25370 82149 -25326
rect 82193 -25370 82249 -25326
rect 82293 -25370 82349 -25326
rect 82393 -25370 82849 -25326
rect 82893 -25370 82949 -25326
rect 82993 -25370 83049 -25326
rect 83093 -25370 83149 -25326
rect 83193 -25370 83249 -25326
rect 83293 -25370 83349 -25326
rect 83393 -25370 83449 -25326
rect 83493 -25370 83549 -25326
rect 83593 -25370 83649 -25326
rect 83693 -25370 83749 -25326
rect 83793 -25370 83849 -25326
rect 83893 -25370 83949 -25326
rect 83993 -25370 84049 -25326
rect 84093 -25370 84149 -25326
rect 84193 -25370 84249 -25326
rect 84293 -25370 84349 -25326
rect 84393 -25370 84849 -25326
rect 84893 -25370 84949 -25326
rect 84993 -25370 85049 -25326
rect 85093 -25370 85149 -25326
rect 85193 -25370 85249 -25326
rect 85293 -25370 85349 -25326
rect 85393 -25370 85449 -25326
rect 85493 -25370 85549 -25326
rect 85593 -25370 85649 -25326
rect 85693 -25370 85749 -25326
rect 85793 -25370 85849 -25326
rect 85893 -25370 85949 -25326
rect 85993 -25370 86049 -25326
rect 86093 -25370 86149 -25326
rect 86193 -25370 86249 -25326
rect 86293 -25370 86349 -25326
rect 86393 -25370 86849 -25326
rect 86893 -25370 86949 -25326
rect 86993 -25370 87049 -25326
rect 87093 -25370 87149 -25326
rect 87193 -25370 87249 -25326
rect 87293 -25370 87349 -25326
rect 87393 -25370 87449 -25326
rect 87493 -25370 87549 -25326
rect 87593 -25370 87649 -25326
rect 87693 -25370 87749 -25326
rect 87793 -25370 87849 -25326
rect 87893 -25370 87949 -25326
rect 87993 -25370 88049 -25326
rect 88093 -25370 88149 -25326
rect 88193 -25370 88249 -25326
rect 88293 -25370 88349 -25326
rect 88393 -25339 109104 -25326
rect 109148 -25339 109204 -25295
rect 109248 -25339 109304 -25295
rect 109348 -25339 109404 -25295
rect 109448 -25339 109504 -25295
rect 109548 -25339 109604 -25295
rect 109648 -25339 109704 -25295
rect 109748 -25339 109804 -25295
rect 109848 -25339 109904 -25295
rect 109948 -25339 110004 -25295
rect 110048 -25339 110104 -25295
rect 110148 -25339 110204 -25295
rect 110248 -25339 110304 -25295
rect 110348 -25339 110404 -25295
rect 110448 -25339 110504 -25295
rect 110548 -25339 110604 -25295
rect 110648 -25339 111104 -25295
rect 111148 -25339 111204 -25295
rect 111248 -25339 111304 -25295
rect 111348 -25339 111404 -25295
rect 111448 -25339 111504 -25295
rect 111548 -25339 111604 -25295
rect 111648 -25339 111704 -25295
rect 111748 -25339 111804 -25295
rect 111848 -25339 111904 -25295
rect 111948 -25339 112004 -25295
rect 112048 -25339 112104 -25295
rect 112148 -25339 112204 -25295
rect 112248 -25339 112304 -25295
rect 112348 -25339 112404 -25295
rect 112448 -25339 112504 -25295
rect 112548 -25339 112604 -25295
rect 112648 -25339 113104 -25295
rect 113148 -25339 113204 -25295
rect 113248 -25339 113304 -25295
rect 113348 -25339 113404 -25295
rect 113448 -25339 113504 -25295
rect 113548 -25339 113604 -25295
rect 113648 -25339 113704 -25295
rect 113748 -25339 113804 -25295
rect 113848 -25339 113904 -25295
rect 113948 -25339 114004 -25295
rect 114048 -25339 114104 -25295
rect 114148 -25339 114204 -25295
rect 114248 -25339 114304 -25295
rect 114348 -25339 114404 -25295
rect 114448 -25339 114504 -25295
rect 114548 -25339 114604 -25295
rect 114648 -25339 115104 -25295
rect 115148 -25339 115204 -25295
rect 115248 -25339 115304 -25295
rect 115348 -25339 115404 -25295
rect 115448 -25339 115504 -25295
rect 115548 -25339 115604 -25295
rect 115648 -25339 115704 -25295
rect 115748 -25339 115804 -25295
rect 115848 -25339 115904 -25295
rect 115948 -25339 116004 -25295
rect 116048 -25339 116104 -25295
rect 116148 -25339 116204 -25295
rect 116248 -25339 116304 -25295
rect 116348 -25339 116404 -25295
rect 116448 -25339 116504 -25295
rect 116548 -25339 116604 -25295
rect 116648 -25339 177360 -25295
rect 88393 -25370 177360 -25339
rect -75255 -25395 177360 -25370
rect -75255 -25410 109104 -25395
rect -109116 -25426 109104 -25410
rect -109116 -25466 80849 -25426
rect -109116 -25510 -82799 -25466
rect -82755 -25510 -82699 -25466
rect -82655 -25510 -82599 -25466
rect -82555 -25510 -82499 -25466
rect -82455 -25510 -82399 -25466
rect -82355 -25510 -82299 -25466
rect -82255 -25510 -82199 -25466
rect -82155 -25510 -82099 -25466
rect -82055 -25510 -81999 -25466
rect -81955 -25510 -81899 -25466
rect -81855 -25510 -81799 -25466
rect -81755 -25510 -81699 -25466
rect -81655 -25510 -81599 -25466
rect -81555 -25510 -81499 -25466
rect -81455 -25510 -81399 -25466
rect -81355 -25510 -81299 -25466
rect -81255 -25510 -80799 -25466
rect -80755 -25510 -80699 -25466
rect -80655 -25510 -80599 -25466
rect -80555 -25510 -80499 -25466
rect -80455 -25510 -80399 -25466
rect -80355 -25510 -80299 -25466
rect -80255 -25510 -80199 -25466
rect -80155 -25510 -80099 -25466
rect -80055 -25510 -79999 -25466
rect -79955 -25510 -79899 -25466
rect -79855 -25510 -79799 -25466
rect -79755 -25510 -79699 -25466
rect -79655 -25510 -79599 -25466
rect -79555 -25510 -79499 -25466
rect -79455 -25510 -79399 -25466
rect -79355 -25510 -79299 -25466
rect -79255 -25510 -78799 -25466
rect -78755 -25510 -78699 -25466
rect -78655 -25510 -78599 -25466
rect -78555 -25510 -78499 -25466
rect -78455 -25510 -78399 -25466
rect -78355 -25510 -78299 -25466
rect -78255 -25510 -78199 -25466
rect -78155 -25510 -78099 -25466
rect -78055 -25510 -77999 -25466
rect -77955 -25510 -77899 -25466
rect -77855 -25510 -77799 -25466
rect -77755 -25510 -77699 -25466
rect -77655 -25510 -77599 -25466
rect -77555 -25510 -77499 -25466
rect -77455 -25510 -77399 -25466
rect -77355 -25510 -77299 -25466
rect -77255 -25510 -76799 -25466
rect -76755 -25510 -76699 -25466
rect -76655 -25510 -76599 -25466
rect -76555 -25510 -76499 -25466
rect -76455 -25510 -76399 -25466
rect -76355 -25510 -76299 -25466
rect -76255 -25510 -76199 -25466
rect -76155 -25510 -76099 -25466
rect -76055 -25510 -75999 -25466
rect -75955 -25510 -75899 -25466
rect -75855 -25510 -75799 -25466
rect -75755 -25510 -75699 -25466
rect -75655 -25510 -75599 -25466
rect -75555 -25510 -75499 -25466
rect -75455 -25510 -75399 -25466
rect -75355 -25510 -75299 -25466
rect -75255 -25470 80849 -25466
rect 80893 -25470 80949 -25426
rect 80993 -25470 81049 -25426
rect 81093 -25470 81149 -25426
rect 81193 -25470 81249 -25426
rect 81293 -25470 81349 -25426
rect 81393 -25470 81449 -25426
rect 81493 -25470 81549 -25426
rect 81593 -25470 81649 -25426
rect 81693 -25470 81749 -25426
rect 81793 -25470 81849 -25426
rect 81893 -25470 81949 -25426
rect 81993 -25470 82049 -25426
rect 82093 -25470 82149 -25426
rect 82193 -25470 82249 -25426
rect 82293 -25470 82349 -25426
rect 82393 -25470 82849 -25426
rect 82893 -25470 82949 -25426
rect 82993 -25470 83049 -25426
rect 83093 -25470 83149 -25426
rect 83193 -25470 83249 -25426
rect 83293 -25470 83349 -25426
rect 83393 -25470 83449 -25426
rect 83493 -25470 83549 -25426
rect 83593 -25470 83649 -25426
rect 83693 -25470 83749 -25426
rect 83793 -25470 83849 -25426
rect 83893 -25470 83949 -25426
rect 83993 -25470 84049 -25426
rect 84093 -25470 84149 -25426
rect 84193 -25470 84249 -25426
rect 84293 -25470 84349 -25426
rect 84393 -25470 84849 -25426
rect 84893 -25470 84949 -25426
rect 84993 -25470 85049 -25426
rect 85093 -25470 85149 -25426
rect 85193 -25470 85249 -25426
rect 85293 -25470 85349 -25426
rect 85393 -25470 85449 -25426
rect 85493 -25470 85549 -25426
rect 85593 -25470 85649 -25426
rect 85693 -25470 85749 -25426
rect 85793 -25470 85849 -25426
rect 85893 -25470 85949 -25426
rect 85993 -25470 86049 -25426
rect 86093 -25470 86149 -25426
rect 86193 -25470 86249 -25426
rect 86293 -25470 86349 -25426
rect 86393 -25470 86849 -25426
rect 86893 -25470 86949 -25426
rect 86993 -25470 87049 -25426
rect 87093 -25470 87149 -25426
rect 87193 -25470 87249 -25426
rect 87293 -25470 87349 -25426
rect 87393 -25470 87449 -25426
rect 87493 -25470 87549 -25426
rect 87593 -25470 87649 -25426
rect 87693 -25470 87749 -25426
rect 87793 -25470 87849 -25426
rect 87893 -25470 87949 -25426
rect 87993 -25470 88049 -25426
rect 88093 -25470 88149 -25426
rect 88193 -25470 88249 -25426
rect 88293 -25470 88349 -25426
rect 88393 -25439 109104 -25426
rect 109148 -25439 109204 -25395
rect 109248 -25439 109304 -25395
rect 109348 -25439 109404 -25395
rect 109448 -25439 109504 -25395
rect 109548 -25439 109604 -25395
rect 109648 -25439 109704 -25395
rect 109748 -25439 109804 -25395
rect 109848 -25439 109904 -25395
rect 109948 -25439 110004 -25395
rect 110048 -25439 110104 -25395
rect 110148 -25439 110204 -25395
rect 110248 -25439 110304 -25395
rect 110348 -25439 110404 -25395
rect 110448 -25439 110504 -25395
rect 110548 -25439 110604 -25395
rect 110648 -25439 111104 -25395
rect 111148 -25439 111204 -25395
rect 111248 -25439 111304 -25395
rect 111348 -25439 111404 -25395
rect 111448 -25439 111504 -25395
rect 111548 -25439 111604 -25395
rect 111648 -25439 111704 -25395
rect 111748 -25439 111804 -25395
rect 111848 -25439 111904 -25395
rect 111948 -25439 112004 -25395
rect 112048 -25439 112104 -25395
rect 112148 -25439 112204 -25395
rect 112248 -25439 112304 -25395
rect 112348 -25439 112404 -25395
rect 112448 -25439 112504 -25395
rect 112548 -25439 112604 -25395
rect 112648 -25439 113104 -25395
rect 113148 -25439 113204 -25395
rect 113248 -25439 113304 -25395
rect 113348 -25439 113404 -25395
rect 113448 -25439 113504 -25395
rect 113548 -25439 113604 -25395
rect 113648 -25439 113704 -25395
rect 113748 -25439 113804 -25395
rect 113848 -25439 113904 -25395
rect 113948 -25439 114004 -25395
rect 114048 -25439 114104 -25395
rect 114148 -25439 114204 -25395
rect 114248 -25439 114304 -25395
rect 114348 -25439 114404 -25395
rect 114448 -25439 114504 -25395
rect 114548 -25439 114604 -25395
rect 114648 -25439 115104 -25395
rect 115148 -25439 115204 -25395
rect 115248 -25439 115304 -25395
rect 115348 -25439 115404 -25395
rect 115448 -25439 115504 -25395
rect 115548 -25439 115604 -25395
rect 115648 -25439 115704 -25395
rect 115748 -25439 115804 -25395
rect 115848 -25439 115904 -25395
rect 115948 -25439 116004 -25395
rect 116048 -25439 116104 -25395
rect 116148 -25439 116204 -25395
rect 116248 -25439 116304 -25395
rect 116348 -25439 116404 -25395
rect 116448 -25439 116504 -25395
rect 116548 -25439 116604 -25395
rect 116648 -25439 177360 -25395
rect 88393 -25470 177360 -25439
rect -75255 -25495 177360 -25470
rect -75255 -25510 109104 -25495
rect -109116 -25526 109104 -25510
rect -109116 -25566 80849 -25526
rect -109116 -25610 -82799 -25566
rect -82755 -25610 -82699 -25566
rect -82655 -25610 -82599 -25566
rect -82555 -25610 -82499 -25566
rect -82455 -25610 -82399 -25566
rect -82355 -25610 -82299 -25566
rect -82255 -25610 -82199 -25566
rect -82155 -25610 -82099 -25566
rect -82055 -25610 -81999 -25566
rect -81955 -25610 -81899 -25566
rect -81855 -25610 -81799 -25566
rect -81755 -25610 -81699 -25566
rect -81655 -25610 -81599 -25566
rect -81555 -25610 -81499 -25566
rect -81455 -25610 -81399 -25566
rect -81355 -25610 -81299 -25566
rect -81255 -25610 -80799 -25566
rect -80755 -25610 -80699 -25566
rect -80655 -25610 -80599 -25566
rect -80555 -25610 -80499 -25566
rect -80455 -25610 -80399 -25566
rect -80355 -25610 -80299 -25566
rect -80255 -25610 -80199 -25566
rect -80155 -25610 -80099 -25566
rect -80055 -25610 -79999 -25566
rect -79955 -25610 -79899 -25566
rect -79855 -25610 -79799 -25566
rect -79755 -25610 -79699 -25566
rect -79655 -25610 -79599 -25566
rect -79555 -25610 -79499 -25566
rect -79455 -25610 -79399 -25566
rect -79355 -25610 -79299 -25566
rect -79255 -25610 -78799 -25566
rect -78755 -25610 -78699 -25566
rect -78655 -25610 -78599 -25566
rect -78555 -25610 -78499 -25566
rect -78455 -25610 -78399 -25566
rect -78355 -25610 -78299 -25566
rect -78255 -25610 -78199 -25566
rect -78155 -25610 -78099 -25566
rect -78055 -25610 -77999 -25566
rect -77955 -25610 -77899 -25566
rect -77855 -25610 -77799 -25566
rect -77755 -25610 -77699 -25566
rect -77655 -25610 -77599 -25566
rect -77555 -25610 -77499 -25566
rect -77455 -25610 -77399 -25566
rect -77355 -25610 -77299 -25566
rect -77255 -25610 -76799 -25566
rect -76755 -25610 -76699 -25566
rect -76655 -25610 -76599 -25566
rect -76555 -25610 -76499 -25566
rect -76455 -25610 -76399 -25566
rect -76355 -25610 -76299 -25566
rect -76255 -25610 -76199 -25566
rect -76155 -25610 -76099 -25566
rect -76055 -25610 -75999 -25566
rect -75955 -25610 -75899 -25566
rect -75855 -25610 -75799 -25566
rect -75755 -25610 -75699 -25566
rect -75655 -25610 -75599 -25566
rect -75555 -25610 -75499 -25566
rect -75455 -25610 -75399 -25566
rect -75355 -25610 -75299 -25566
rect -75255 -25570 80849 -25566
rect 80893 -25570 80949 -25526
rect 80993 -25570 81049 -25526
rect 81093 -25570 81149 -25526
rect 81193 -25570 81249 -25526
rect 81293 -25570 81349 -25526
rect 81393 -25570 81449 -25526
rect 81493 -25570 81549 -25526
rect 81593 -25570 81649 -25526
rect 81693 -25570 81749 -25526
rect 81793 -25570 81849 -25526
rect 81893 -25570 81949 -25526
rect 81993 -25570 82049 -25526
rect 82093 -25570 82149 -25526
rect 82193 -25570 82249 -25526
rect 82293 -25570 82349 -25526
rect 82393 -25570 82849 -25526
rect 82893 -25570 82949 -25526
rect 82993 -25570 83049 -25526
rect 83093 -25570 83149 -25526
rect 83193 -25570 83249 -25526
rect 83293 -25570 83349 -25526
rect 83393 -25570 83449 -25526
rect 83493 -25570 83549 -25526
rect 83593 -25570 83649 -25526
rect 83693 -25570 83749 -25526
rect 83793 -25570 83849 -25526
rect 83893 -25570 83949 -25526
rect 83993 -25570 84049 -25526
rect 84093 -25570 84149 -25526
rect 84193 -25570 84249 -25526
rect 84293 -25570 84349 -25526
rect 84393 -25570 84849 -25526
rect 84893 -25570 84949 -25526
rect 84993 -25570 85049 -25526
rect 85093 -25570 85149 -25526
rect 85193 -25570 85249 -25526
rect 85293 -25570 85349 -25526
rect 85393 -25570 85449 -25526
rect 85493 -25570 85549 -25526
rect 85593 -25570 85649 -25526
rect 85693 -25570 85749 -25526
rect 85793 -25570 85849 -25526
rect 85893 -25570 85949 -25526
rect 85993 -25570 86049 -25526
rect 86093 -25570 86149 -25526
rect 86193 -25570 86249 -25526
rect 86293 -25570 86349 -25526
rect 86393 -25570 86849 -25526
rect 86893 -25570 86949 -25526
rect 86993 -25570 87049 -25526
rect 87093 -25570 87149 -25526
rect 87193 -25570 87249 -25526
rect 87293 -25570 87349 -25526
rect 87393 -25570 87449 -25526
rect 87493 -25570 87549 -25526
rect 87593 -25570 87649 -25526
rect 87693 -25570 87749 -25526
rect 87793 -25570 87849 -25526
rect 87893 -25570 87949 -25526
rect 87993 -25570 88049 -25526
rect 88093 -25570 88149 -25526
rect 88193 -25570 88249 -25526
rect 88293 -25570 88349 -25526
rect 88393 -25539 109104 -25526
rect 109148 -25539 109204 -25495
rect 109248 -25539 109304 -25495
rect 109348 -25539 109404 -25495
rect 109448 -25539 109504 -25495
rect 109548 -25539 109604 -25495
rect 109648 -25539 109704 -25495
rect 109748 -25539 109804 -25495
rect 109848 -25539 109904 -25495
rect 109948 -25539 110004 -25495
rect 110048 -25539 110104 -25495
rect 110148 -25539 110204 -25495
rect 110248 -25539 110304 -25495
rect 110348 -25539 110404 -25495
rect 110448 -25539 110504 -25495
rect 110548 -25539 110604 -25495
rect 110648 -25539 111104 -25495
rect 111148 -25539 111204 -25495
rect 111248 -25539 111304 -25495
rect 111348 -25539 111404 -25495
rect 111448 -25539 111504 -25495
rect 111548 -25539 111604 -25495
rect 111648 -25539 111704 -25495
rect 111748 -25539 111804 -25495
rect 111848 -25539 111904 -25495
rect 111948 -25539 112004 -25495
rect 112048 -25539 112104 -25495
rect 112148 -25539 112204 -25495
rect 112248 -25539 112304 -25495
rect 112348 -25539 112404 -25495
rect 112448 -25539 112504 -25495
rect 112548 -25539 112604 -25495
rect 112648 -25539 113104 -25495
rect 113148 -25539 113204 -25495
rect 113248 -25539 113304 -25495
rect 113348 -25539 113404 -25495
rect 113448 -25539 113504 -25495
rect 113548 -25539 113604 -25495
rect 113648 -25539 113704 -25495
rect 113748 -25539 113804 -25495
rect 113848 -25539 113904 -25495
rect 113948 -25539 114004 -25495
rect 114048 -25539 114104 -25495
rect 114148 -25539 114204 -25495
rect 114248 -25539 114304 -25495
rect 114348 -25539 114404 -25495
rect 114448 -25539 114504 -25495
rect 114548 -25539 114604 -25495
rect 114648 -25539 115104 -25495
rect 115148 -25539 115204 -25495
rect 115248 -25539 115304 -25495
rect 115348 -25539 115404 -25495
rect 115448 -25539 115504 -25495
rect 115548 -25539 115604 -25495
rect 115648 -25539 115704 -25495
rect 115748 -25539 115804 -25495
rect 115848 -25539 115904 -25495
rect 115948 -25539 116004 -25495
rect 116048 -25539 116104 -25495
rect 116148 -25539 116204 -25495
rect 116248 -25539 116304 -25495
rect 116348 -25539 116404 -25495
rect 116448 -25539 116504 -25495
rect 116548 -25539 116604 -25495
rect 116648 -25539 177360 -25495
rect 88393 -25570 177360 -25539
rect -75255 -25595 177360 -25570
rect -75255 -25610 109104 -25595
rect -109116 -25639 109104 -25610
rect 109148 -25639 109204 -25595
rect 109248 -25639 109304 -25595
rect 109348 -25639 109404 -25595
rect 109448 -25639 109504 -25595
rect 109548 -25639 109604 -25595
rect 109648 -25639 109704 -25595
rect 109748 -25639 109804 -25595
rect 109848 -25639 109904 -25595
rect 109948 -25639 110004 -25595
rect 110048 -25639 110104 -25595
rect 110148 -25639 110204 -25595
rect 110248 -25639 110304 -25595
rect 110348 -25639 110404 -25595
rect 110448 -25639 110504 -25595
rect 110548 -25639 110604 -25595
rect 110648 -25639 111104 -25595
rect 111148 -25639 111204 -25595
rect 111248 -25639 111304 -25595
rect 111348 -25639 111404 -25595
rect 111448 -25639 111504 -25595
rect 111548 -25639 111604 -25595
rect 111648 -25639 111704 -25595
rect 111748 -25639 111804 -25595
rect 111848 -25639 111904 -25595
rect 111948 -25639 112004 -25595
rect 112048 -25639 112104 -25595
rect 112148 -25639 112204 -25595
rect 112248 -25639 112304 -25595
rect 112348 -25639 112404 -25595
rect 112448 -25639 112504 -25595
rect 112548 -25639 112604 -25595
rect 112648 -25639 113104 -25595
rect 113148 -25639 113204 -25595
rect 113248 -25639 113304 -25595
rect 113348 -25639 113404 -25595
rect 113448 -25639 113504 -25595
rect 113548 -25639 113604 -25595
rect 113648 -25639 113704 -25595
rect 113748 -25639 113804 -25595
rect 113848 -25639 113904 -25595
rect 113948 -25639 114004 -25595
rect 114048 -25639 114104 -25595
rect 114148 -25639 114204 -25595
rect 114248 -25639 114304 -25595
rect 114348 -25639 114404 -25595
rect 114448 -25639 114504 -25595
rect 114548 -25639 114604 -25595
rect 114648 -25639 115104 -25595
rect 115148 -25639 115204 -25595
rect 115248 -25639 115304 -25595
rect 115348 -25639 115404 -25595
rect 115448 -25639 115504 -25595
rect 115548 -25639 115604 -25595
rect 115648 -25639 115704 -25595
rect 115748 -25639 115804 -25595
rect 115848 -25639 115904 -25595
rect 115948 -25639 116004 -25595
rect 116048 -25639 116104 -25595
rect 116148 -25639 116204 -25595
rect 116248 -25639 116304 -25595
rect 116348 -25639 116404 -25595
rect 116448 -25639 116504 -25595
rect 116548 -25639 116604 -25595
rect 116648 -25639 177360 -25595
rect -109116 -25666 177360 -25639
rect -109116 -25710 -82799 -25666
rect -82755 -25710 -82699 -25666
rect -82655 -25710 -82599 -25666
rect -82555 -25710 -82499 -25666
rect -82455 -25710 -82399 -25666
rect -82355 -25710 -82299 -25666
rect -82255 -25710 -82199 -25666
rect -82155 -25710 -82099 -25666
rect -82055 -25710 -81999 -25666
rect -81955 -25710 -81899 -25666
rect -81855 -25710 -81799 -25666
rect -81755 -25710 -81699 -25666
rect -81655 -25710 -81599 -25666
rect -81555 -25710 -81499 -25666
rect -81455 -25710 -81399 -25666
rect -81355 -25710 -81299 -25666
rect -81255 -25710 -80799 -25666
rect -80755 -25710 -80699 -25666
rect -80655 -25710 -80599 -25666
rect -80555 -25710 -80499 -25666
rect -80455 -25710 -80399 -25666
rect -80355 -25710 -80299 -25666
rect -80255 -25710 -80199 -25666
rect -80155 -25710 -80099 -25666
rect -80055 -25710 -79999 -25666
rect -79955 -25710 -79899 -25666
rect -79855 -25710 -79799 -25666
rect -79755 -25710 -79699 -25666
rect -79655 -25710 -79599 -25666
rect -79555 -25710 -79499 -25666
rect -79455 -25710 -79399 -25666
rect -79355 -25710 -79299 -25666
rect -79255 -25710 -78799 -25666
rect -78755 -25710 -78699 -25666
rect -78655 -25710 -78599 -25666
rect -78555 -25710 -78499 -25666
rect -78455 -25710 -78399 -25666
rect -78355 -25710 -78299 -25666
rect -78255 -25710 -78199 -25666
rect -78155 -25710 -78099 -25666
rect -78055 -25710 -77999 -25666
rect -77955 -25710 -77899 -25666
rect -77855 -25710 -77799 -25666
rect -77755 -25710 -77699 -25666
rect -77655 -25710 -77599 -25666
rect -77555 -25710 -77499 -25666
rect -77455 -25710 -77399 -25666
rect -77355 -25710 -77299 -25666
rect -77255 -25710 -76799 -25666
rect -76755 -25710 -76699 -25666
rect -76655 -25710 -76599 -25666
rect -76555 -25710 -76499 -25666
rect -76455 -25710 -76399 -25666
rect -76355 -25710 -76299 -25666
rect -76255 -25710 -76199 -25666
rect -76155 -25710 -76099 -25666
rect -76055 -25710 -75999 -25666
rect -75955 -25710 -75899 -25666
rect -75855 -25710 -75799 -25666
rect -75755 -25710 -75699 -25666
rect -75655 -25710 -75599 -25666
rect -75555 -25710 -75499 -25666
rect -75455 -25710 -75399 -25666
rect -75355 -25710 -75299 -25666
rect -75255 -25695 177360 -25666
rect -75255 -25710 109104 -25695
rect -109116 -25739 109104 -25710
rect 109148 -25739 109204 -25695
rect 109248 -25739 109304 -25695
rect 109348 -25739 109404 -25695
rect 109448 -25739 109504 -25695
rect 109548 -25739 109604 -25695
rect 109648 -25739 109704 -25695
rect 109748 -25739 109804 -25695
rect 109848 -25739 109904 -25695
rect 109948 -25739 110004 -25695
rect 110048 -25739 110104 -25695
rect 110148 -25739 110204 -25695
rect 110248 -25739 110304 -25695
rect 110348 -25739 110404 -25695
rect 110448 -25739 110504 -25695
rect 110548 -25739 110604 -25695
rect 110648 -25739 111104 -25695
rect 111148 -25739 111204 -25695
rect 111248 -25739 111304 -25695
rect 111348 -25739 111404 -25695
rect 111448 -25739 111504 -25695
rect 111548 -25739 111604 -25695
rect 111648 -25739 111704 -25695
rect 111748 -25739 111804 -25695
rect 111848 -25739 111904 -25695
rect 111948 -25739 112004 -25695
rect 112048 -25739 112104 -25695
rect 112148 -25739 112204 -25695
rect 112248 -25739 112304 -25695
rect 112348 -25739 112404 -25695
rect 112448 -25739 112504 -25695
rect 112548 -25739 112604 -25695
rect 112648 -25739 113104 -25695
rect 113148 -25739 113204 -25695
rect 113248 -25739 113304 -25695
rect 113348 -25739 113404 -25695
rect 113448 -25739 113504 -25695
rect 113548 -25739 113604 -25695
rect 113648 -25739 113704 -25695
rect 113748 -25739 113804 -25695
rect 113848 -25739 113904 -25695
rect 113948 -25739 114004 -25695
rect 114048 -25739 114104 -25695
rect 114148 -25739 114204 -25695
rect 114248 -25739 114304 -25695
rect 114348 -25739 114404 -25695
rect 114448 -25739 114504 -25695
rect 114548 -25739 114604 -25695
rect 114648 -25739 115104 -25695
rect 115148 -25739 115204 -25695
rect 115248 -25739 115304 -25695
rect 115348 -25739 115404 -25695
rect 115448 -25739 115504 -25695
rect 115548 -25739 115604 -25695
rect 115648 -25739 115704 -25695
rect 115748 -25739 115804 -25695
rect 115848 -25739 115904 -25695
rect 115948 -25739 116004 -25695
rect 116048 -25739 116104 -25695
rect 116148 -25739 116204 -25695
rect 116248 -25739 116304 -25695
rect 116348 -25739 116404 -25695
rect 116448 -25739 116504 -25695
rect 116548 -25739 116604 -25695
rect 116648 -25739 177360 -25695
rect -109116 -25766 177360 -25739
rect -109116 -25810 -82799 -25766
rect -82755 -25810 -82699 -25766
rect -82655 -25810 -82599 -25766
rect -82555 -25810 -82499 -25766
rect -82455 -25810 -82399 -25766
rect -82355 -25810 -82299 -25766
rect -82255 -25810 -82199 -25766
rect -82155 -25810 -82099 -25766
rect -82055 -25810 -81999 -25766
rect -81955 -25810 -81899 -25766
rect -81855 -25810 -81799 -25766
rect -81755 -25810 -81699 -25766
rect -81655 -25810 -81599 -25766
rect -81555 -25810 -81499 -25766
rect -81455 -25810 -81399 -25766
rect -81355 -25810 -81299 -25766
rect -81255 -25810 -80799 -25766
rect -80755 -25810 -80699 -25766
rect -80655 -25810 -80599 -25766
rect -80555 -25810 -80499 -25766
rect -80455 -25810 -80399 -25766
rect -80355 -25810 -80299 -25766
rect -80255 -25810 -80199 -25766
rect -80155 -25810 -80099 -25766
rect -80055 -25810 -79999 -25766
rect -79955 -25810 -79899 -25766
rect -79855 -25810 -79799 -25766
rect -79755 -25810 -79699 -25766
rect -79655 -25810 -79599 -25766
rect -79555 -25810 -79499 -25766
rect -79455 -25810 -79399 -25766
rect -79355 -25810 -79299 -25766
rect -79255 -25810 -78799 -25766
rect -78755 -25810 -78699 -25766
rect -78655 -25810 -78599 -25766
rect -78555 -25810 -78499 -25766
rect -78455 -25810 -78399 -25766
rect -78355 -25810 -78299 -25766
rect -78255 -25810 -78199 -25766
rect -78155 -25810 -78099 -25766
rect -78055 -25810 -77999 -25766
rect -77955 -25810 -77899 -25766
rect -77855 -25810 -77799 -25766
rect -77755 -25810 -77699 -25766
rect -77655 -25810 -77599 -25766
rect -77555 -25810 -77499 -25766
rect -77455 -25810 -77399 -25766
rect -77355 -25810 -77299 -25766
rect -77255 -25810 -76799 -25766
rect -76755 -25810 -76699 -25766
rect -76655 -25810 -76599 -25766
rect -76555 -25810 -76499 -25766
rect -76455 -25810 -76399 -25766
rect -76355 -25810 -76299 -25766
rect -76255 -25810 -76199 -25766
rect -76155 -25810 -76099 -25766
rect -76055 -25810 -75999 -25766
rect -75955 -25810 -75899 -25766
rect -75855 -25810 -75799 -25766
rect -75755 -25810 -75699 -25766
rect -75655 -25810 -75599 -25766
rect -75555 -25810 -75499 -25766
rect -75455 -25810 -75399 -25766
rect -75355 -25810 -75299 -25766
rect -75255 -25810 177360 -25766
rect -109116 -25866 177360 -25810
rect -109116 -25910 -82799 -25866
rect -82755 -25910 -82699 -25866
rect -82655 -25910 -82599 -25866
rect -82555 -25910 -82499 -25866
rect -82455 -25910 -82399 -25866
rect -82355 -25910 -82299 -25866
rect -82255 -25910 -82199 -25866
rect -82155 -25910 -82099 -25866
rect -82055 -25910 -81999 -25866
rect -81955 -25910 -81899 -25866
rect -81855 -25910 -81799 -25866
rect -81755 -25910 -81699 -25866
rect -81655 -25910 -81599 -25866
rect -81555 -25910 -81499 -25866
rect -81455 -25910 -81399 -25866
rect -81355 -25910 -81299 -25866
rect -81255 -25910 -80799 -25866
rect -80755 -25910 -80699 -25866
rect -80655 -25910 -80599 -25866
rect -80555 -25910 -80499 -25866
rect -80455 -25910 -80399 -25866
rect -80355 -25910 -80299 -25866
rect -80255 -25910 -80199 -25866
rect -80155 -25910 -80099 -25866
rect -80055 -25910 -79999 -25866
rect -79955 -25910 -79899 -25866
rect -79855 -25910 -79799 -25866
rect -79755 -25910 -79699 -25866
rect -79655 -25910 -79599 -25866
rect -79555 -25910 -79499 -25866
rect -79455 -25910 -79399 -25866
rect -79355 -25910 -79299 -25866
rect -79255 -25910 -78799 -25866
rect -78755 -25910 -78699 -25866
rect -78655 -25910 -78599 -25866
rect -78555 -25910 -78499 -25866
rect -78455 -25910 -78399 -25866
rect -78355 -25910 -78299 -25866
rect -78255 -25910 -78199 -25866
rect -78155 -25910 -78099 -25866
rect -78055 -25910 -77999 -25866
rect -77955 -25910 -77899 -25866
rect -77855 -25910 -77799 -25866
rect -77755 -25910 -77699 -25866
rect -77655 -25910 -77599 -25866
rect -77555 -25910 -77499 -25866
rect -77455 -25910 -77399 -25866
rect -77355 -25910 -77299 -25866
rect -77255 -25910 -76799 -25866
rect -76755 -25910 -76699 -25866
rect -76655 -25910 -76599 -25866
rect -76555 -25910 -76499 -25866
rect -76455 -25910 -76399 -25866
rect -76355 -25910 -76299 -25866
rect -76255 -25910 -76199 -25866
rect -76155 -25910 -76099 -25866
rect -76055 -25910 -75999 -25866
rect -75955 -25910 -75899 -25866
rect -75855 -25910 -75799 -25866
rect -75755 -25910 -75699 -25866
rect -75655 -25910 -75599 -25866
rect -75555 -25910 -75499 -25866
rect -75455 -25910 -75399 -25866
rect -75355 -25910 -75299 -25866
rect -75255 -25910 177360 -25866
rect -109116 -27203 177360 -25910
rect -109116 -28117 -109040 -27203
rect -108508 -28117 -108432 -27203
rect -107900 -28117 -107824 -27203
rect -107292 -28117 -107216 -27203
rect -106684 -28117 -106608 -27203
rect -106076 -28117 -106000 -27203
rect -105468 -28117 -105392 -27203
rect -104860 -28117 -104784 -27203
rect -104252 -28117 -104176 -27203
rect -103644 -28117 -103568 -27203
rect -103036 -28117 -102960 -27203
rect -102428 -28117 -102352 -27203
rect -101820 -28117 -101744 -27203
rect -101212 -28117 -101136 -27203
rect -100604 -28117 -100528 -27203
rect -99996 -28117 -99920 -27203
rect -99388 -28117 -99312 -27203
rect -98780 -28117 -98704 -27203
rect -98172 -28117 -98096 -27203
rect -97564 -28117 -97488 -27203
rect -96956 -28117 -96880 -27203
rect -96348 -28117 -96272 -27203
rect -95740 -28117 -95664 -27203
rect -95132 -28117 -95056 -27203
rect -94524 -28117 -94448 -27203
rect -93916 -28117 -93840 -27203
rect -93308 -28117 -93232 -27203
rect -92700 -28117 -92624 -27203
rect -92092 -28117 -92016 -27203
rect -91484 -28117 -91408 -27203
rect -90876 -28117 -90800 -27203
rect -90268 -28117 -90192 -27203
rect -89660 -28117 -89584 -27203
rect -89052 -28117 -88976 -27203
rect -88444 -28117 -88368 -27203
rect -87836 -28117 -87760 -27203
rect -87228 -28117 -87152 -27203
rect -86620 -28117 -86544 -27203
rect -86012 -28117 -85936 -27203
rect -85404 -28117 -85328 -27203
rect -84796 -28117 -84720 -27203
rect -84188 -28117 -84112 -27203
rect -83580 -28117 -83504 -27203
rect -82972 -28117 -82896 -27203
rect -82364 -28117 -82288 -27203
rect -81756 -28117 -81680 -27203
rect -81148 -28117 -81072 -27203
rect -80540 -28117 -80464 -27203
rect -79932 -28117 -79856 -27203
rect -79324 -28117 -79248 -27203
rect -78716 -28117 -78640 -27203
rect -77116 -28117 -77040 -27203
rect -76508 -28117 -76432 -27203
rect -75900 -28117 -75824 -27203
rect -75292 -28117 -75216 -27203
rect -74684 -28117 -74608 -27203
rect -74076 -28117 -74000 -27203
rect -73468 -28117 -73392 -27203
rect -72860 -28117 -72784 -27203
rect -72252 -28117 -72176 -27203
rect -71644 -28117 -71568 -27203
rect -71036 -28117 -70960 -27203
rect -70428 -28117 -70352 -27203
rect -69820 -28117 -69744 -27203
rect -69212 -28117 -69136 -27203
rect -68604 -28117 -68528 -27203
rect -67996 -28117 -67920 -27203
rect -67388 -28117 -67312 -27203
rect -66780 -28117 -66704 -27203
rect -66172 -28117 -66096 -27203
rect -65564 -28117 -65488 -27203
rect -64956 -28117 -64880 -27203
rect -64348 -28117 -64272 -27203
rect -63740 -28117 -63664 -27203
rect -63132 -28117 -63056 -27203
rect -62524 -28117 -62448 -27203
rect -61916 -28117 -61840 -27203
rect -61308 -28117 -61232 -27203
rect -60700 -28117 -60624 -27203
rect -60092 -28117 -60016 -27203
rect -59484 -28117 -59408 -27203
rect -58876 -28117 -58800 -27203
rect -58268 -28117 -58192 -27203
rect -57660 -28117 -57584 -27203
rect -57052 -28117 -56976 -27203
rect -56444 -28117 -56368 -27203
rect -55836 -28117 -55760 -27203
rect -55228 -28117 -55152 -27203
rect -54620 -28117 -54544 -27203
rect -54012 -28117 -53936 -27203
rect -53404 -28117 -53328 -27203
rect -52796 -28117 -52720 -27203
rect -52188 -28117 -52112 -27203
rect -51580 -28117 -51504 -27203
rect -50972 -28117 -50896 -27203
rect -50364 -28117 -50288 -27203
rect -49756 -28117 -49680 -27203
rect -49148 -28117 -49072 -27203
rect -48540 -28117 -48464 -27203
rect -47932 -28117 -47856 -27203
rect -47324 -28117 -47248 -27203
rect -46716 -28117 -46640 -27203
rect -45116 -28117 -45040 -27203
rect -44508 -28117 -44432 -27203
rect -43900 -28117 -43824 -27203
rect -43292 -28117 -43216 -27203
rect -42684 -28117 -42608 -27203
rect -42076 -28117 -42000 -27203
rect -41468 -28117 -41392 -27203
rect -40860 -28117 -40784 -27203
rect -40252 -28117 -40176 -27203
rect -39644 -28117 -39568 -27203
rect -39036 -28117 -38960 -27203
rect -38428 -28117 -38352 -27203
rect -37820 -28117 -37744 -27203
rect -37212 -28117 -37136 -27203
rect -36604 -28117 -36528 -27203
rect -35996 -28117 -35920 -27203
rect -35388 -28117 -35312 -27203
rect -34780 -28117 -34704 -27203
rect -34172 -28117 -34096 -27203
rect -33564 -28117 -33488 -27203
rect -32956 -28117 -32880 -27203
rect -32348 -28117 -32272 -27203
rect -31740 -28117 -31664 -27203
rect -31132 -28117 -31056 -27203
rect -30524 -28117 -30448 -27203
rect -29916 -28117 -29840 -27203
rect -29308 -28117 -29232 -27203
rect -28700 -28117 -28624 -27203
rect -28092 -28117 -28016 -27203
rect -27484 -28117 -27408 -27203
rect -26876 -28117 -26800 -27203
rect -26268 -28117 -26192 -27203
rect -25660 -28117 -25584 -27203
rect -25052 -28117 -24976 -27203
rect -24444 -28117 -24368 -27203
rect -23836 -28117 -23760 -27203
rect -23228 -28117 -23152 -27203
rect -22620 -28117 -22544 -27203
rect -22012 -28117 -21936 -27203
rect -21404 -28117 -21328 -27203
rect -20796 -28117 -20720 -27203
rect -20188 -28117 -20112 -27203
rect -19580 -28117 -19504 -27203
rect -18972 -28117 -18896 -27203
rect -18364 -28117 -18288 -27203
rect -17756 -28117 -17680 -27203
rect -17148 -28117 -17072 -27203
rect -16540 -28117 -16464 -27203
rect -15932 -28117 -15856 -27203
rect -15324 -28117 -15248 -27203
rect -14716 -28117 -14640 -27203
rect -13116 -28117 -13040 -27203
rect -12508 -28117 -12432 -27203
rect -11900 -28117 -11824 -27203
rect -11292 -28117 -11216 -27203
rect -10684 -28117 -10608 -27203
rect -10076 -28117 -10000 -27203
rect -9468 -28117 -9392 -27203
rect -8860 -28117 -8784 -27203
rect -8252 -28117 -8176 -27203
rect -7644 -28117 -7568 -27203
rect -7036 -28117 -6960 -27203
rect -6428 -28117 -6352 -27203
rect -5820 -28117 -5744 -27203
rect -5212 -28117 -5136 -27203
rect -4604 -28117 -4528 -27203
rect -3996 -28117 -3920 -27203
rect -3388 -28117 -3312 -27203
rect -2780 -28117 -2704 -27203
rect -2172 -28117 -2096 -27203
rect -1564 -28117 -1488 -27203
rect -956 -28117 -880 -27203
rect -348 -28117 -272 -27203
rect 260 -28117 336 -27203
rect 868 -28117 944 -27203
rect 1476 -28117 1552 -27203
rect 2084 -28117 2160 -27203
rect 2692 -28117 2768 -27203
rect 3300 -28117 3376 -27203
rect 3908 -28117 3984 -27203
rect 4516 -28117 4592 -27203
rect 5124 -28117 5200 -27203
rect 5732 -28117 5808 -27203
rect 6340 -28117 6416 -27203
rect 6948 -28117 7024 -27203
rect 7556 -28117 7632 -27203
rect 8164 -28117 8240 -27203
rect 8772 -28117 8848 -27203
rect 9380 -28117 9456 -27203
rect 9988 -28117 10064 -27203
rect 10596 -28117 10672 -27203
rect 11204 -28117 11280 -27203
rect 11812 -28117 11888 -27203
rect 12420 -28117 12496 -27203
rect 13028 -28117 13104 -27203
rect 13636 -28117 13712 -27203
rect 14244 -28117 14320 -27203
rect 14852 -28117 14928 -27203
rect 15460 -28117 15536 -27203
rect 16068 -28117 16144 -27203
rect 16676 -28117 16752 -27203
rect 17284 -28117 17360 -27203
rect 18884 -28117 18960 -27203
rect 19492 -28117 19568 -27203
rect 20100 -28117 20176 -27203
rect 20708 -28117 20784 -27203
rect 21316 -28117 21392 -27203
rect 21924 -28117 22000 -27203
rect 22532 -28117 22608 -27203
rect 23140 -28117 23216 -27203
rect 23748 -28117 23824 -27203
rect 24356 -28117 24432 -27203
rect 24964 -28117 25040 -27203
rect 25572 -28117 25648 -27203
rect 26180 -28117 26256 -27203
rect 26788 -28117 26864 -27203
rect 27396 -28117 27472 -27203
rect 28004 -28117 28080 -27203
rect 28612 -28117 28688 -27203
rect 29220 -28117 29296 -27203
rect 29828 -28117 29904 -27203
rect 30436 -28117 30512 -27203
rect 31044 -28117 31120 -27203
rect 31652 -28117 31728 -27203
rect 32260 -28117 32336 -27203
rect 32868 -28117 32944 -27203
rect 33476 -28117 33552 -27203
rect 34084 -28117 34160 -27203
rect 34692 -28117 34768 -27203
rect 35300 -28117 35376 -27203
rect 35908 -28117 35984 -27203
rect 36516 -28117 36592 -27203
rect 37124 -28117 37200 -27203
rect 37732 -28117 37808 -27203
rect 38340 -28117 38416 -27203
rect 38948 -28117 39024 -27203
rect 39556 -28117 39632 -27203
rect 40164 -28117 40240 -27203
rect 40772 -28117 40848 -27203
rect 41380 -28117 41456 -27203
rect 41988 -28117 42064 -27203
rect 42596 -28117 42672 -27203
rect 43204 -28117 43280 -27203
rect 43812 -28117 43888 -27203
rect 44420 -28117 44496 -27203
rect 45028 -28117 45104 -27203
rect 45636 -28117 45712 -27203
rect 46244 -28117 46320 -27203
rect 46852 -28117 46928 -27203
rect 47460 -28117 47536 -27203
rect 48068 -28117 48144 -27203
rect 48676 -28117 48752 -27203
rect 49284 -28117 49360 -27203
rect 50884 -28117 50960 -27203
rect 51492 -28117 51568 -27203
rect 52100 -28117 52176 -27203
rect 52708 -28117 52784 -27203
rect 53316 -28117 53392 -27203
rect 53924 -28117 54000 -27203
rect 54532 -28117 54608 -27203
rect 55140 -28117 55216 -27203
rect 55748 -28117 55824 -27203
rect 56356 -28117 56432 -27203
rect 56964 -28117 57040 -27203
rect 57572 -28117 57648 -27203
rect 58180 -28117 58256 -27203
rect 58788 -28117 58864 -27203
rect 59396 -28117 59472 -27203
rect 60004 -28117 60080 -27203
rect 60612 -28117 60688 -27203
rect 61220 -28117 61296 -27203
rect 61828 -28117 61904 -27203
rect 62436 -28117 62512 -27203
rect 63044 -28117 63120 -27203
rect 63652 -28117 63728 -27203
rect 64260 -28117 64336 -27203
rect 64868 -28117 64944 -27203
rect 65476 -28117 65552 -27203
rect 66084 -28117 66160 -27203
rect 66692 -28117 66768 -27203
rect 67300 -28117 67376 -27203
rect 67908 -28117 67984 -27203
rect 68516 -28117 68592 -27203
rect 69124 -28117 69200 -27203
rect 69732 -28117 69808 -27203
rect 70340 -28117 70416 -27203
rect 70948 -28117 71024 -27203
rect 71556 -28117 71632 -27203
rect 72164 -28117 72240 -27203
rect 72772 -28117 72848 -27203
rect 73380 -28117 73456 -27203
rect 73988 -28117 74064 -27203
rect 74596 -28117 74672 -27203
rect 75204 -28117 75280 -27203
rect 75812 -28117 75888 -27203
rect 76420 -28117 76496 -27203
rect 77028 -28117 77104 -27203
rect 77636 -28117 77712 -27203
rect 78244 -28117 78320 -27203
rect 78852 -28117 78928 -27203
rect 79460 -28117 79536 -27203
rect 80068 -28117 80144 -27203
rect 80676 -28117 80752 -27203
rect 81284 -28117 81360 -27203
rect 82884 -28117 82960 -27203
rect 83492 -28117 83568 -27203
rect 84100 -28117 84176 -27203
rect 84708 -28117 84784 -27203
rect 85316 -28117 85392 -27203
rect 85924 -28117 86000 -27203
rect 86532 -28117 86608 -27203
rect 87140 -28117 87216 -27203
rect 87748 -28117 87824 -27203
rect 88356 -28117 88432 -27203
rect 88964 -28117 89040 -27203
rect 89572 -28117 89648 -27203
rect 90180 -28117 90256 -27203
rect 90788 -28117 90864 -27203
rect 91396 -28117 91472 -27203
rect 92004 -28117 92080 -27203
rect 92612 -28117 92688 -27203
rect 93220 -28117 93296 -27203
rect 93828 -28117 93904 -27203
rect 94436 -28117 94512 -27203
rect 95044 -28117 95120 -27203
rect 95652 -28117 95728 -27203
rect 96260 -28117 96336 -27203
rect 96868 -28117 96944 -27203
rect 97476 -28117 97552 -27203
rect 98084 -28117 98160 -27203
rect 98692 -28117 98768 -27203
rect 99300 -28117 99376 -27203
rect 99908 -28117 99984 -27203
rect 100516 -28117 100592 -27203
rect 101124 -28117 101200 -27203
rect 101732 -28117 101808 -27203
rect 102340 -28117 102416 -27203
rect 102948 -28117 103024 -27203
rect 103556 -28117 103632 -27203
rect 104164 -28117 104240 -27203
rect 104772 -28117 104848 -27203
rect 105380 -28117 105456 -27203
rect 105988 -28117 106064 -27203
rect 106596 -28117 106672 -27203
rect 107204 -28117 107280 -27203
rect 107812 -28117 107888 -27203
rect 108420 -28117 108496 -27203
rect 109028 -28117 109104 -27203
rect 109636 -28117 109712 -27203
rect 110244 -28117 110320 -27203
rect 110852 -28117 110928 -27203
rect 111460 -28117 111536 -27203
rect 112068 -28117 112144 -27203
rect 112676 -28117 112752 -27203
rect 113284 -28117 113360 -27203
rect 114884 -28117 114960 -27203
rect 115492 -28117 115568 -27203
rect 116100 -28117 116176 -27203
rect 116708 -28117 116784 -27203
rect 117316 -28117 117392 -27203
rect 117924 -28117 118000 -27203
rect 118532 -28117 118608 -27203
rect 119140 -28117 119216 -27203
rect 119748 -28117 119824 -27203
rect 120356 -28117 120432 -27203
rect 120964 -28117 121040 -27203
rect 121572 -28117 121648 -27203
rect 122180 -28117 122256 -27203
rect 122788 -28117 122864 -27203
rect 123396 -28117 123472 -27203
rect 124004 -28117 124080 -27203
rect 124612 -28117 124688 -27203
rect 125220 -28117 125296 -27203
rect 125828 -28117 125904 -27203
rect 126436 -28117 126512 -27203
rect 127044 -28117 127120 -27203
rect 127652 -28117 127728 -27203
rect 128260 -28117 128336 -27203
rect 128868 -28117 128944 -27203
rect 129476 -28117 129552 -27203
rect 130084 -28117 130160 -27203
rect 130692 -28117 130768 -27203
rect 131300 -28117 131376 -27203
rect 131908 -28117 131984 -27203
rect 132516 -28117 132592 -27203
rect 133124 -28117 133200 -27203
rect 133732 -28117 133808 -27203
rect 134340 -28117 134416 -27203
rect 134948 -28117 135024 -27203
rect 135556 -28117 135632 -27203
rect 136164 -28117 136240 -27203
rect 136772 -28117 136848 -27203
rect 137380 -28117 137456 -27203
rect 137988 -28117 138064 -27203
rect 138596 -28117 138672 -27203
rect 139204 -28117 139280 -27203
rect 139812 -28117 139888 -27203
rect 140420 -28117 140496 -27203
rect 141028 -28117 141104 -27203
rect 141636 -28117 141712 -27203
rect 142244 -28117 142320 -27203
rect 142852 -28117 142928 -27203
rect 143460 -28117 143536 -27203
rect 144068 -28117 144144 -27203
rect 144676 -28117 144752 -27203
rect 145284 -28117 145360 -27203
rect 146884 -28117 146960 -27203
rect 147492 -28117 147568 -27203
rect 148100 -28117 148176 -27203
rect 148708 -28117 148784 -27203
rect 149316 -28117 149392 -27203
rect 149924 -28117 150000 -27203
rect 150532 -28117 150608 -27203
rect 151140 -28117 151216 -27203
rect 151748 -28117 151824 -27203
rect 152356 -28117 152432 -27203
rect 152964 -28117 153040 -27203
rect 153572 -28117 153648 -27203
rect 154180 -28117 154256 -27203
rect 154788 -28117 154864 -27203
rect 155396 -28117 155472 -27203
rect 156004 -28117 156080 -27203
rect 156612 -28117 156688 -27203
rect 157220 -28117 157296 -27203
rect 157828 -28117 157904 -27203
rect 158436 -28117 158512 -27203
rect 159044 -28117 159120 -27203
rect 159652 -28117 159728 -27203
rect 160260 -28117 160336 -27203
rect 160868 -28117 160944 -27203
rect 161476 -28117 161552 -27203
rect 162084 -28117 162160 -27203
rect 162692 -28117 162768 -27203
rect 163300 -28117 163376 -27203
rect 163908 -28117 163984 -27203
rect 164516 -28117 164592 -27203
rect 165124 -28117 165200 -27203
rect 165732 -28117 165808 -27203
rect 166340 -28117 166416 -27203
rect 166948 -28117 167024 -27203
rect 167556 -28117 167632 -27203
rect 168164 -28117 168240 -27203
rect 168772 -28117 168848 -27203
rect 169380 -28117 169456 -27203
rect 169988 -28117 170064 -27203
rect 170596 -28117 170672 -27203
rect 171204 -28117 171280 -27203
rect 171812 -28117 171888 -27203
rect 172420 -28117 172496 -27203
rect 173028 -28117 173104 -27203
rect 173636 -28117 173712 -27203
rect 174244 -28117 174320 -27203
rect 174852 -28117 174928 -27203
rect 175460 -28117 175536 -27203
rect 176068 -28117 176144 -27203
rect 176676 -28117 176752 -27203
rect 177284 -28117 177360 -27203
rect -131554 -34142 -126400 -32005
rect -131554 -35301 -130077 -34142
rect -128909 -35301 -126400 -34142
rect -131554 -38091 -126400 -35301
rect -114442 -171279 -109186 -28119
rect -77274 -48121 -77040 -28119
rect -45274 -48121 -45040 -28119
rect -13274 -48121 -13040 -28119
rect 18726 -48121 18960 -28119
rect 50726 -48121 50960 -28119
rect 82726 -48121 82960 -28119
rect 114726 -48121 114960 -28119
rect 146726 -48121 146960 -28119
rect -108812 -49035 -108736 -48121
rect -108204 -49035 -108128 -48121
rect -107596 -49035 -107520 -48121
rect -106988 -49035 -106912 -48121
rect -106380 -49035 -106304 -48121
rect -105772 -49035 -105696 -48121
rect -105164 -49035 -105088 -48121
rect -104556 -49035 -104480 -48121
rect -103948 -49035 -103872 -48121
rect -103340 -49035 -103264 -48121
rect -102732 -49035 -102656 -48121
rect -102124 -49035 -102048 -48121
rect -101516 -49035 -101440 -48121
rect -100908 -49035 -100832 -48121
rect -100300 -49035 -100224 -48121
rect -99692 -49035 -99616 -48121
rect -99084 -49035 -99008 -48121
rect -98476 -49035 -98400 -48121
rect -97868 -49035 -97792 -48121
rect -97260 -49035 -97184 -48121
rect -96652 -49035 -96576 -48121
rect -96044 -49035 -95968 -48121
rect -95436 -49035 -95360 -48121
rect -94828 -49035 -94752 -48121
rect -94220 -49035 -94144 -48121
rect -93612 -49035 -93536 -48121
rect -93004 -49035 -92928 -48121
rect -92396 -49035 -92320 -48121
rect -91788 -49035 -91712 -48121
rect -91180 -49035 -91104 -48121
rect -90572 -49035 -90496 -48121
rect -89964 -49035 -89888 -48121
rect -89356 -49035 -89280 -48121
rect -88748 -49035 -88672 -48121
rect -88140 -49035 -88064 -48121
rect -87532 -49035 -87456 -48121
rect -86924 -49035 -86848 -48121
rect -86316 -49035 -86240 -48121
rect -85708 -49035 -85632 -48121
rect -85100 -49035 -85024 -48121
rect -84492 -49035 -84416 -48121
rect -83884 -49035 -83808 -48121
rect -83276 -49035 -83200 -48121
rect -82668 -49035 -82592 -48121
rect -82060 -49035 -81984 -48121
rect -81452 -49035 -81376 -48121
rect -80844 -49035 -80768 -48121
rect -80236 -49035 -80160 -48121
rect -79628 -49035 -79552 -48121
rect -79020 -49035 -78944 -48121
rect -76812 -49035 -76736 -48121
rect -76204 -49035 -76128 -48121
rect -75596 -49035 -75520 -48121
rect -74988 -49035 -74912 -48121
rect -74380 -49035 -74304 -48121
rect -73772 -49035 -73696 -48121
rect -73164 -49035 -73088 -48121
rect -72556 -49035 -72480 -48121
rect -71948 -49035 -71872 -48121
rect -71340 -49035 -71264 -48121
rect -70732 -49035 -70656 -48121
rect -70124 -49035 -70048 -48121
rect -69516 -49035 -69440 -48121
rect -68908 -49035 -68832 -48121
rect -68300 -49035 -68224 -48121
rect -67692 -49035 -67616 -48121
rect -67084 -49035 -67008 -48121
rect -66476 -49035 -66400 -48121
rect -65868 -49035 -65792 -48121
rect -65260 -49035 -65184 -48121
rect -64652 -49035 -64576 -48121
rect -64044 -49035 -63968 -48121
rect -63436 -49035 -63360 -48121
rect -62828 -49035 -62752 -48121
rect -62220 -49035 -62144 -48121
rect -61612 -49035 -61536 -48121
rect -61004 -49035 -60928 -48121
rect -60396 -49035 -60320 -48121
rect -59788 -49035 -59712 -48121
rect -59180 -49035 -59104 -48121
rect -58572 -49035 -58496 -48121
rect -57964 -49035 -57888 -48121
rect -57356 -49035 -57280 -48121
rect -56748 -49035 -56672 -48121
rect -56140 -49035 -56064 -48121
rect -55532 -49035 -55456 -48121
rect -54924 -49035 -54848 -48121
rect -54316 -49035 -54240 -48121
rect -53708 -49035 -53632 -48121
rect -53100 -49035 -53024 -48121
rect -52492 -49035 -52416 -48121
rect -51884 -49035 -51808 -48121
rect -51276 -49035 -51200 -48121
rect -50668 -49035 -50592 -48121
rect -50060 -49035 -49984 -48121
rect -49452 -49035 -49376 -48121
rect -48844 -49035 -48768 -48121
rect -48236 -49035 -48160 -48121
rect -47628 -49035 -47552 -48121
rect -47020 -49035 -46944 -48121
rect -44812 -49035 -44736 -48121
rect -44204 -49035 -44128 -48121
rect -43596 -49035 -43520 -48121
rect -42988 -49035 -42912 -48121
rect -42380 -49035 -42304 -48121
rect -41772 -49035 -41696 -48121
rect -41164 -49035 -41088 -48121
rect -40556 -49035 -40480 -48121
rect -39948 -49035 -39872 -48121
rect -39340 -49035 -39264 -48121
rect -38732 -49035 -38656 -48121
rect -38124 -49035 -38048 -48121
rect -37516 -49035 -37440 -48121
rect -36908 -49035 -36832 -48121
rect -36300 -49035 -36224 -48121
rect -35692 -49035 -35616 -48121
rect -35084 -49035 -35008 -48121
rect -34476 -49035 -34400 -48121
rect -33868 -49035 -33792 -48121
rect -33260 -49035 -33184 -48121
rect -32652 -49035 -32576 -48121
rect -32044 -49035 -31968 -48121
rect -31436 -49035 -31360 -48121
rect -30828 -49035 -30752 -48121
rect -30220 -49035 -30144 -48121
rect -29612 -49035 -29536 -48121
rect -29004 -49035 -28928 -48121
rect -28396 -49035 -28320 -48121
rect -27788 -49035 -27712 -48121
rect -27180 -49035 -27104 -48121
rect -26572 -49035 -26496 -48121
rect -25964 -49035 -25888 -48121
rect -25356 -49035 -25280 -48121
rect -24748 -49035 -24672 -48121
rect -24140 -49035 -24064 -48121
rect -23532 -49035 -23456 -48121
rect -22924 -49035 -22848 -48121
rect -22316 -49035 -22240 -48121
rect -21708 -49035 -21632 -48121
rect -21100 -49035 -21024 -48121
rect -20492 -49035 -20416 -48121
rect -19884 -49035 -19808 -48121
rect -19276 -49035 -19200 -48121
rect -18668 -49035 -18592 -48121
rect -18060 -49035 -17984 -48121
rect -17452 -49035 -17376 -48121
rect -16844 -49035 -16768 -48121
rect -16236 -49035 -16160 -48121
rect -15628 -49035 -15552 -48121
rect -15020 -49035 -14944 -48121
rect -12812 -49035 -12736 -48121
rect -12204 -49035 -12128 -48121
rect -11596 -49035 -11520 -48121
rect -10988 -49035 -10912 -48121
rect -10380 -49035 -10304 -48121
rect -9772 -49035 -9696 -48121
rect -9164 -49035 -9088 -48121
rect -8556 -49035 -8480 -48121
rect -7948 -49035 -7872 -48121
rect -7340 -49035 -7264 -48121
rect -6732 -49035 -6656 -48121
rect -6124 -49035 -6048 -48121
rect -5516 -49035 -5440 -48121
rect -4908 -49035 -4832 -48121
rect -4300 -49035 -4224 -48121
rect -3692 -49035 -3616 -48121
rect -3084 -49035 -3008 -48121
rect -2476 -49035 -2400 -48121
rect -1868 -49035 -1792 -48121
rect -1260 -49035 -1184 -48121
rect -652 -49035 -576 -48121
rect -44 -49035 32 -48121
rect 564 -49035 640 -48121
rect 1172 -49035 1248 -48121
rect 1780 -49035 1856 -48121
rect 2388 -49035 2464 -48121
rect 2996 -49035 3072 -48121
rect 3604 -49035 3680 -48121
rect 4212 -49035 4288 -48121
rect 4820 -49035 4896 -48121
rect 5428 -49035 5504 -48121
rect 6036 -49035 6112 -48121
rect 6644 -49035 6720 -48121
rect 7252 -49035 7328 -48121
rect 7860 -49035 7936 -48121
rect 8468 -49035 8544 -48121
rect 9076 -49035 9152 -48121
rect 9684 -49035 9760 -48121
rect 10292 -49035 10368 -48121
rect 10900 -49035 10976 -48121
rect 11508 -49035 11584 -48121
rect 12116 -49035 12192 -48121
rect 12724 -49035 12800 -48121
rect 13332 -49035 13408 -48121
rect 13940 -49035 14016 -48121
rect 14548 -49035 14624 -48121
rect 15156 -49035 15232 -48121
rect 15764 -49035 15840 -48121
rect 16372 -49035 16448 -48121
rect 16980 -49035 17056 -48121
rect 19188 -49035 19264 -48121
rect 19796 -49035 19872 -48121
rect 20404 -49035 20480 -48121
rect 21012 -49035 21088 -48121
rect 21620 -49035 21696 -48121
rect 22228 -49035 22304 -48121
rect 22836 -49035 22912 -48121
rect 23444 -49035 23520 -48121
rect 24052 -49035 24128 -48121
rect 24660 -49035 24736 -48121
rect 25268 -49035 25344 -48121
rect 25876 -49035 25952 -48121
rect 26484 -49035 26560 -48121
rect 27092 -49035 27168 -48121
rect 27700 -49035 27776 -48121
rect 28308 -49035 28384 -48121
rect 28916 -49035 28992 -48121
rect 29524 -49035 29600 -48121
rect 30132 -49035 30208 -48121
rect 30740 -49035 30816 -48121
rect 31348 -49035 31424 -48121
rect 31956 -49035 32032 -48121
rect 32564 -49035 32640 -48121
rect 33172 -49035 33248 -48121
rect 33780 -49035 33856 -48121
rect 34388 -49035 34464 -48121
rect 34996 -49035 35072 -48121
rect 35604 -49035 35680 -48121
rect 36212 -49035 36288 -48121
rect 36820 -49035 36896 -48121
rect 37428 -49035 37504 -48121
rect 38036 -49035 38112 -48121
rect 38644 -49035 38720 -48121
rect 39252 -49035 39328 -48121
rect 39860 -49035 39936 -48121
rect 40468 -49035 40544 -48121
rect 41076 -49035 41152 -48121
rect 41684 -49035 41760 -48121
rect 42292 -49035 42368 -48121
rect 42900 -49035 42976 -48121
rect 43508 -49035 43584 -48121
rect 44116 -49035 44192 -48121
rect 44724 -49035 44800 -48121
rect 45332 -49035 45408 -48121
rect 45940 -49035 46016 -48121
rect 46548 -49035 46624 -48121
rect 47156 -49035 47232 -48121
rect 47764 -49035 47840 -48121
rect 48372 -49035 48448 -48121
rect 48980 -49035 49056 -48121
rect 51188 -49035 51264 -48121
rect 51796 -49035 51872 -48121
rect 52404 -49035 52480 -48121
rect 53012 -49035 53088 -48121
rect 53620 -49035 53696 -48121
rect 54228 -49035 54304 -48121
rect 54836 -49035 54912 -48121
rect 55444 -49035 55520 -48121
rect 56052 -49035 56128 -48121
rect 56660 -49035 56736 -48121
rect 57268 -49035 57344 -48121
rect 57876 -49035 57952 -48121
rect 58484 -49035 58560 -48121
rect 59092 -49035 59168 -48121
rect 59700 -49035 59776 -48121
rect 60308 -49035 60384 -48121
rect 60916 -49035 60992 -48121
rect 61524 -49035 61600 -48121
rect 62132 -49035 62208 -48121
rect 62740 -49035 62816 -48121
rect 63348 -49035 63424 -48121
rect 63956 -49035 64032 -48121
rect 64564 -49035 64640 -48121
rect 65172 -49035 65248 -48121
rect 65780 -49035 65856 -48121
rect 66388 -49035 66464 -48121
rect 66996 -49035 67072 -48121
rect 67604 -49035 67680 -48121
rect 68212 -49035 68288 -48121
rect 68820 -49035 68896 -48121
rect 69428 -49035 69504 -48121
rect 70036 -49035 70112 -48121
rect 70644 -49035 70720 -48121
rect 71252 -49035 71328 -48121
rect 71860 -49035 71936 -48121
rect 72468 -49035 72544 -48121
rect 73076 -49035 73152 -48121
rect 73684 -49035 73760 -48121
rect 74292 -49035 74368 -48121
rect 74900 -49035 74976 -48121
rect 75508 -49035 75584 -48121
rect 76116 -49035 76192 -48121
rect 76724 -49035 76800 -48121
rect 77332 -49035 77408 -48121
rect 77940 -49035 78016 -48121
rect 78548 -49035 78624 -48121
rect 79156 -49035 79232 -48121
rect 79764 -49035 79840 -48121
rect 80372 -49035 80448 -48121
rect 80980 -49035 81056 -48121
rect 83188 -49035 83264 -48121
rect 83796 -49035 83872 -48121
rect 84404 -49035 84480 -48121
rect 85012 -49035 85088 -48121
rect 85620 -49035 85696 -48121
rect 86228 -49035 86304 -48121
rect 86836 -49035 86912 -48121
rect 87444 -49035 87520 -48121
rect 88052 -49035 88128 -48121
rect 88660 -49035 88736 -48121
rect 89268 -49035 89344 -48121
rect 89876 -49035 89952 -48121
rect 90484 -49035 90560 -48121
rect 91092 -49035 91168 -48121
rect 91700 -49035 91776 -48121
rect 92308 -49035 92384 -48121
rect 92916 -49035 92992 -48121
rect 93524 -49035 93600 -48121
rect 94132 -49035 94208 -48121
rect 94740 -49035 94816 -48121
rect 95348 -49035 95424 -48121
rect 95956 -49035 96032 -48121
rect 96564 -49035 96640 -48121
rect 97172 -49035 97248 -48121
rect 97780 -49035 97856 -48121
rect 98388 -49035 98464 -48121
rect 98996 -49035 99072 -48121
rect 99604 -49035 99680 -48121
rect 100212 -49035 100288 -48121
rect 100820 -49035 100896 -48121
rect 101428 -49035 101504 -48121
rect 102036 -49035 102112 -48121
rect 102644 -49035 102720 -48121
rect 103252 -49035 103328 -48121
rect 103860 -49035 103936 -48121
rect 104468 -49035 104544 -48121
rect 105076 -49035 105152 -48121
rect 105684 -49035 105760 -48121
rect 106292 -49035 106368 -48121
rect 106900 -49035 106976 -48121
rect 107508 -49035 107584 -48121
rect 108116 -49035 108192 -48121
rect 108724 -49035 108800 -48121
rect 109332 -49035 109408 -48121
rect 109940 -49035 110016 -48121
rect 110548 -49035 110624 -48121
rect 111156 -49035 111232 -48121
rect 111764 -49035 111840 -48121
rect 112372 -49035 112448 -48121
rect 112980 -49035 113056 -48121
rect 115188 -49035 115264 -48121
rect 115796 -49035 115872 -48121
rect 116404 -49035 116480 -48121
rect 117012 -49035 117088 -48121
rect 117620 -49035 117696 -48121
rect 118228 -49035 118304 -48121
rect 118836 -49035 118912 -48121
rect 119444 -49035 119520 -48121
rect 120052 -49035 120128 -48121
rect 120660 -49035 120736 -48121
rect 121268 -49035 121344 -48121
rect 121876 -49035 121952 -48121
rect 122484 -49035 122560 -48121
rect 123092 -49035 123168 -48121
rect 123700 -49035 123776 -48121
rect 124308 -49035 124384 -48121
rect 124916 -49035 124992 -48121
rect 125524 -49035 125600 -48121
rect 126132 -49035 126208 -48121
rect 126740 -49035 126816 -48121
rect 127348 -49035 127424 -48121
rect 127956 -49035 128032 -48121
rect 128564 -49035 128640 -48121
rect 129172 -49035 129248 -48121
rect 129780 -49035 129856 -48121
rect 130388 -49035 130464 -48121
rect 130996 -49035 131072 -48121
rect 131604 -49035 131680 -48121
rect 132212 -49035 132288 -48121
rect 132820 -49035 132896 -48121
rect 133428 -49035 133504 -48121
rect 134036 -49035 134112 -48121
rect 134644 -49035 134720 -48121
rect 135252 -49035 135328 -48121
rect 135860 -49035 135936 -48121
rect 136468 -49035 136544 -48121
rect 137076 -49035 137152 -48121
rect 137684 -49035 137760 -48121
rect 138292 -49035 138368 -48121
rect 138900 -49035 138976 -48121
rect 139508 -49035 139584 -48121
rect 140116 -49035 140192 -48121
rect 140724 -49035 140800 -48121
rect 141332 -49035 141408 -48121
rect 141940 -49035 142016 -48121
rect 142548 -49035 142624 -48121
rect 143156 -49035 143232 -48121
rect 143764 -49035 143840 -48121
rect 144372 -49035 144448 -48121
rect 144980 -49035 145056 -48121
rect 147188 -49035 147264 -48121
rect 147796 -49035 147872 -48121
rect 148404 -49035 148480 -48121
rect 149012 -49035 149088 -48121
rect 149620 -49035 149696 -48121
rect 150228 -49035 150304 -48121
rect 150836 -49035 150912 -48121
rect 151444 -49035 151520 -48121
rect 152052 -49035 152128 -48121
rect 152660 -49035 152736 -48121
rect 153268 -49035 153344 -48121
rect 153876 -49035 153952 -48121
rect 154484 -49035 154560 -48121
rect 155092 -49035 155168 -48121
rect 155700 -49035 155776 -48121
rect 156308 -49035 156384 -48121
rect 156916 -49035 156992 -48121
rect 157524 -49035 157600 -48121
rect 158132 -49035 158208 -48121
rect 158740 -49035 158816 -48121
rect 159348 -49035 159424 -48121
rect 159956 -49035 160032 -48121
rect 160564 -49035 160640 -48121
rect 161172 -49035 161248 -48121
rect 161780 -49035 161856 -48121
rect 162388 -49035 162464 -48121
rect 162996 -49035 163072 -48121
rect 163604 -49035 163680 -48121
rect 164212 -49035 164288 -48121
rect 164820 -49035 164896 -48121
rect 165428 -49035 165504 -48121
rect 166036 -49035 166112 -48121
rect 166644 -49035 166720 -48121
rect 167252 -49035 167328 -48121
rect 167860 -49035 167936 -48121
rect 168468 -49035 168544 -48121
rect 169076 -49035 169152 -48121
rect 169684 -49035 169760 -48121
rect 170292 -49035 170368 -48121
rect 170900 -49035 170976 -48121
rect 171508 -49035 171584 -48121
rect 172116 -49035 172192 -48121
rect 172724 -49035 172800 -48121
rect 173332 -49035 173408 -48121
rect 173940 -49035 174016 -48121
rect 174548 -49035 174624 -48121
rect 175156 -49035 175232 -48121
rect 175764 -49035 175840 -48121
rect 176372 -49035 176448 -48121
rect 176980 -49035 177056 -48121
rect -108812 -49602 178308 -49035
rect 108496 -51137 117196 -50572
rect 108496 -51181 109305 -51137
rect 109349 -51181 109405 -51137
rect 109449 -51181 109505 -51137
rect 109549 -51181 109605 -51137
rect 109649 -51181 109705 -51137
rect 109749 -51181 109805 -51137
rect 109849 -51181 109905 -51137
rect 109949 -51181 110005 -51137
rect 110049 -51181 110105 -51137
rect 110149 -51181 110205 -51137
rect 110249 -51181 110305 -51137
rect 110349 -51181 110405 -51137
rect 110449 -51181 110505 -51137
rect 110549 -51181 110605 -51137
rect 110649 -51181 110705 -51137
rect 110749 -51181 110805 -51137
rect 110849 -51181 111305 -51137
rect 111349 -51181 111405 -51137
rect 111449 -51181 111505 -51137
rect 111549 -51181 111605 -51137
rect 111649 -51181 111705 -51137
rect 111749 -51181 111805 -51137
rect 111849 -51181 111905 -51137
rect 111949 -51181 112005 -51137
rect 112049 -51181 112105 -51137
rect 112149 -51181 112205 -51137
rect 112249 -51181 112305 -51137
rect 112349 -51181 112405 -51137
rect 112449 -51181 112505 -51137
rect 112549 -51181 112605 -51137
rect 112649 -51181 112705 -51137
rect 112749 -51181 112805 -51137
rect 112849 -51181 113305 -51137
rect 113349 -51181 113405 -51137
rect 113449 -51181 113505 -51137
rect 113549 -51181 113605 -51137
rect 113649 -51181 113705 -51137
rect 113749 -51181 113805 -51137
rect 113849 -51181 113905 -51137
rect 113949 -51181 114005 -51137
rect 114049 -51181 114105 -51137
rect 114149 -51181 114205 -51137
rect 114249 -51181 114305 -51137
rect 114349 -51181 114405 -51137
rect 114449 -51181 114505 -51137
rect 114549 -51181 114605 -51137
rect 114649 -51181 114705 -51137
rect 114749 -51181 114805 -51137
rect 114849 -51181 115305 -51137
rect 115349 -51181 115405 -51137
rect 115449 -51181 115505 -51137
rect 115549 -51181 115605 -51137
rect 115649 -51181 115705 -51137
rect 115749 -51181 115805 -51137
rect 115849 -51181 115905 -51137
rect 115949 -51181 116005 -51137
rect 116049 -51181 116105 -51137
rect 116149 -51181 116205 -51137
rect 116249 -51181 116305 -51137
rect 116349 -51181 116405 -51137
rect 116449 -51181 116505 -51137
rect 116549 -51181 116605 -51137
rect 116649 -51181 116705 -51137
rect 116749 -51181 116805 -51137
rect 116849 -51181 117196 -51137
rect 108496 -51237 117196 -51181
rect 108496 -51281 109305 -51237
rect 109349 -51281 109405 -51237
rect 109449 -51281 109505 -51237
rect 109549 -51281 109605 -51237
rect 109649 -51281 109705 -51237
rect 109749 -51281 109805 -51237
rect 109849 -51281 109905 -51237
rect 109949 -51281 110005 -51237
rect 110049 -51281 110105 -51237
rect 110149 -51281 110205 -51237
rect 110249 -51281 110305 -51237
rect 110349 -51281 110405 -51237
rect 110449 -51281 110505 -51237
rect 110549 -51281 110605 -51237
rect 110649 -51281 110705 -51237
rect 110749 -51281 110805 -51237
rect 110849 -51281 111305 -51237
rect 111349 -51281 111405 -51237
rect 111449 -51281 111505 -51237
rect 111549 -51281 111605 -51237
rect 111649 -51281 111705 -51237
rect 111749 -51281 111805 -51237
rect 111849 -51281 111905 -51237
rect 111949 -51281 112005 -51237
rect 112049 -51281 112105 -51237
rect 112149 -51281 112205 -51237
rect 112249 -51281 112305 -51237
rect 112349 -51281 112405 -51237
rect 112449 -51281 112505 -51237
rect 112549 -51281 112605 -51237
rect 112649 -51281 112705 -51237
rect 112749 -51281 112805 -51237
rect 112849 -51281 113305 -51237
rect 113349 -51281 113405 -51237
rect 113449 -51281 113505 -51237
rect 113549 -51281 113605 -51237
rect 113649 -51281 113705 -51237
rect 113749 -51281 113805 -51237
rect 113849 -51281 113905 -51237
rect 113949 -51281 114005 -51237
rect 114049 -51281 114105 -51237
rect 114149 -51281 114205 -51237
rect 114249 -51281 114305 -51237
rect 114349 -51281 114405 -51237
rect 114449 -51281 114505 -51237
rect 114549 -51281 114605 -51237
rect 114649 -51281 114705 -51237
rect 114749 -51281 114805 -51237
rect 114849 -51281 115305 -51237
rect 115349 -51281 115405 -51237
rect 115449 -51281 115505 -51237
rect 115549 -51281 115605 -51237
rect 115649 -51281 115705 -51237
rect 115749 -51281 115805 -51237
rect 115849 -51281 115905 -51237
rect 115949 -51281 116005 -51237
rect 116049 -51281 116105 -51237
rect 116149 -51281 116205 -51237
rect 116249 -51281 116305 -51237
rect 116349 -51281 116405 -51237
rect 116449 -51281 116505 -51237
rect 116549 -51281 116605 -51237
rect 116649 -51281 116705 -51237
rect 116749 -51281 116805 -51237
rect 116849 -51281 117196 -51237
rect 108496 -51337 117196 -51281
rect 108496 -51381 109305 -51337
rect 109349 -51381 109405 -51337
rect 109449 -51381 109505 -51337
rect 109549 -51381 109605 -51337
rect 109649 -51381 109705 -51337
rect 109749 -51381 109805 -51337
rect 109849 -51381 109905 -51337
rect 109949 -51381 110005 -51337
rect 110049 -51381 110105 -51337
rect 110149 -51381 110205 -51337
rect 110249 -51381 110305 -51337
rect 110349 -51381 110405 -51337
rect 110449 -51381 110505 -51337
rect 110549 -51381 110605 -51337
rect 110649 -51381 110705 -51337
rect 110749 -51381 110805 -51337
rect 110849 -51381 111305 -51337
rect 111349 -51381 111405 -51337
rect 111449 -51381 111505 -51337
rect 111549 -51381 111605 -51337
rect 111649 -51381 111705 -51337
rect 111749 -51381 111805 -51337
rect 111849 -51381 111905 -51337
rect 111949 -51381 112005 -51337
rect 112049 -51381 112105 -51337
rect 112149 -51381 112205 -51337
rect 112249 -51381 112305 -51337
rect 112349 -51381 112405 -51337
rect 112449 -51381 112505 -51337
rect 112549 -51381 112605 -51337
rect 112649 -51381 112705 -51337
rect 112749 -51381 112805 -51337
rect 112849 -51381 113305 -51337
rect 113349 -51381 113405 -51337
rect 113449 -51381 113505 -51337
rect 113549 -51381 113605 -51337
rect 113649 -51381 113705 -51337
rect 113749 -51381 113805 -51337
rect 113849 -51381 113905 -51337
rect 113949 -51381 114005 -51337
rect 114049 -51381 114105 -51337
rect 114149 -51381 114205 -51337
rect 114249 -51381 114305 -51337
rect 114349 -51381 114405 -51337
rect 114449 -51381 114505 -51337
rect 114549 -51381 114605 -51337
rect 114649 -51381 114705 -51337
rect 114749 -51381 114805 -51337
rect 114849 -51381 115305 -51337
rect 115349 -51381 115405 -51337
rect 115449 -51381 115505 -51337
rect 115549 -51381 115605 -51337
rect 115649 -51381 115705 -51337
rect 115749 -51381 115805 -51337
rect 115849 -51381 115905 -51337
rect 115949 -51381 116005 -51337
rect 116049 -51381 116105 -51337
rect 116149 -51381 116205 -51337
rect 116249 -51381 116305 -51337
rect 116349 -51381 116405 -51337
rect 116449 -51381 116505 -51337
rect 116549 -51381 116605 -51337
rect 116649 -51381 116705 -51337
rect 116749 -51381 116805 -51337
rect 116849 -51381 117196 -51337
rect 108496 -51437 117196 -51381
rect 108496 -51481 109305 -51437
rect 109349 -51481 109405 -51437
rect 109449 -51481 109505 -51437
rect 109549 -51481 109605 -51437
rect 109649 -51481 109705 -51437
rect 109749 -51481 109805 -51437
rect 109849 -51481 109905 -51437
rect 109949 -51481 110005 -51437
rect 110049 -51481 110105 -51437
rect 110149 -51481 110205 -51437
rect 110249 -51481 110305 -51437
rect 110349 -51481 110405 -51437
rect 110449 -51481 110505 -51437
rect 110549 -51481 110605 -51437
rect 110649 -51481 110705 -51437
rect 110749 -51481 110805 -51437
rect 110849 -51481 111305 -51437
rect 111349 -51481 111405 -51437
rect 111449 -51481 111505 -51437
rect 111549 -51481 111605 -51437
rect 111649 -51481 111705 -51437
rect 111749 -51481 111805 -51437
rect 111849 -51481 111905 -51437
rect 111949 -51481 112005 -51437
rect 112049 -51481 112105 -51437
rect 112149 -51481 112205 -51437
rect 112249 -51481 112305 -51437
rect 112349 -51481 112405 -51437
rect 112449 -51481 112505 -51437
rect 112549 -51481 112605 -51437
rect 112649 -51481 112705 -51437
rect 112749 -51481 112805 -51437
rect 112849 -51481 113305 -51437
rect 113349 -51481 113405 -51437
rect 113449 -51481 113505 -51437
rect 113549 -51481 113605 -51437
rect 113649 -51481 113705 -51437
rect 113749 -51481 113805 -51437
rect 113849 -51481 113905 -51437
rect 113949 -51481 114005 -51437
rect 114049 -51481 114105 -51437
rect 114149 -51481 114205 -51437
rect 114249 -51481 114305 -51437
rect 114349 -51481 114405 -51437
rect 114449 -51481 114505 -51437
rect 114549 -51481 114605 -51437
rect 114649 -51481 114705 -51437
rect 114749 -51481 114805 -51437
rect 114849 -51481 115305 -51437
rect 115349 -51481 115405 -51437
rect 115449 -51481 115505 -51437
rect 115549 -51481 115605 -51437
rect 115649 -51481 115705 -51437
rect 115749 -51481 115805 -51437
rect 115849 -51481 115905 -51437
rect 115949 -51481 116005 -51437
rect 116049 -51481 116105 -51437
rect 116149 -51481 116205 -51437
rect 116249 -51481 116305 -51437
rect 116349 -51481 116405 -51437
rect 116449 -51481 116505 -51437
rect 116549 -51481 116605 -51437
rect 116649 -51481 116705 -51437
rect 116749 -51481 116805 -51437
rect 116849 -51481 117196 -51437
rect 108496 -51537 117196 -51481
rect 108496 -51581 109305 -51537
rect 109349 -51581 109405 -51537
rect 109449 -51581 109505 -51537
rect 109549 -51581 109605 -51537
rect 109649 -51581 109705 -51537
rect 109749 -51581 109805 -51537
rect 109849 -51581 109905 -51537
rect 109949 -51581 110005 -51537
rect 110049 -51581 110105 -51537
rect 110149 -51581 110205 -51537
rect 110249 -51581 110305 -51537
rect 110349 -51581 110405 -51537
rect 110449 -51581 110505 -51537
rect 110549 -51581 110605 -51537
rect 110649 -51581 110705 -51537
rect 110749 -51581 110805 -51537
rect 110849 -51581 111305 -51537
rect 111349 -51581 111405 -51537
rect 111449 -51581 111505 -51537
rect 111549 -51581 111605 -51537
rect 111649 -51581 111705 -51537
rect 111749 -51581 111805 -51537
rect 111849 -51581 111905 -51537
rect 111949 -51581 112005 -51537
rect 112049 -51581 112105 -51537
rect 112149 -51581 112205 -51537
rect 112249 -51581 112305 -51537
rect 112349 -51581 112405 -51537
rect 112449 -51581 112505 -51537
rect 112549 -51581 112605 -51537
rect 112649 -51581 112705 -51537
rect 112749 -51581 112805 -51537
rect 112849 -51581 113305 -51537
rect 113349 -51581 113405 -51537
rect 113449 -51581 113505 -51537
rect 113549 -51581 113605 -51537
rect 113649 -51581 113705 -51537
rect 113749 -51581 113805 -51537
rect 113849 -51581 113905 -51537
rect 113949 -51581 114005 -51537
rect 114049 -51581 114105 -51537
rect 114149 -51581 114205 -51537
rect 114249 -51581 114305 -51537
rect 114349 -51581 114405 -51537
rect 114449 -51581 114505 -51537
rect 114549 -51581 114605 -51537
rect 114649 -51581 114705 -51537
rect 114749 -51581 114805 -51537
rect 114849 -51581 115305 -51537
rect 115349 -51581 115405 -51537
rect 115449 -51581 115505 -51537
rect 115549 -51581 115605 -51537
rect 115649 -51581 115705 -51537
rect 115749 -51581 115805 -51537
rect 115849 -51581 115905 -51537
rect 115949 -51581 116005 -51537
rect 116049 -51581 116105 -51537
rect 116149 -51581 116205 -51537
rect 116249 -51581 116305 -51537
rect 116349 -51581 116405 -51537
rect 116449 -51581 116505 -51537
rect 116549 -51581 116605 -51537
rect 116649 -51581 116705 -51537
rect 116749 -51581 116805 -51537
rect 116849 -51581 117196 -51537
rect 108496 -51637 117196 -51581
rect 108496 -51681 109305 -51637
rect 109349 -51681 109405 -51637
rect 109449 -51681 109505 -51637
rect 109549 -51681 109605 -51637
rect 109649 -51681 109705 -51637
rect 109749 -51681 109805 -51637
rect 109849 -51681 109905 -51637
rect 109949 -51681 110005 -51637
rect 110049 -51681 110105 -51637
rect 110149 -51681 110205 -51637
rect 110249 -51681 110305 -51637
rect 110349 -51681 110405 -51637
rect 110449 -51681 110505 -51637
rect 110549 -51681 110605 -51637
rect 110649 -51681 110705 -51637
rect 110749 -51681 110805 -51637
rect 110849 -51681 111305 -51637
rect 111349 -51681 111405 -51637
rect 111449 -51681 111505 -51637
rect 111549 -51681 111605 -51637
rect 111649 -51681 111705 -51637
rect 111749 -51681 111805 -51637
rect 111849 -51681 111905 -51637
rect 111949 -51681 112005 -51637
rect 112049 -51681 112105 -51637
rect 112149 -51681 112205 -51637
rect 112249 -51681 112305 -51637
rect 112349 -51681 112405 -51637
rect 112449 -51681 112505 -51637
rect 112549 -51681 112605 -51637
rect 112649 -51681 112705 -51637
rect 112749 -51681 112805 -51637
rect 112849 -51681 113305 -51637
rect 113349 -51681 113405 -51637
rect 113449 -51681 113505 -51637
rect 113549 -51681 113605 -51637
rect 113649 -51681 113705 -51637
rect 113749 -51681 113805 -51637
rect 113849 -51681 113905 -51637
rect 113949 -51681 114005 -51637
rect 114049 -51681 114105 -51637
rect 114149 -51681 114205 -51637
rect 114249 -51681 114305 -51637
rect 114349 -51681 114405 -51637
rect 114449 -51681 114505 -51637
rect 114549 -51681 114605 -51637
rect 114649 -51681 114705 -51637
rect 114749 -51681 114805 -51637
rect 114849 -51681 115305 -51637
rect 115349 -51681 115405 -51637
rect 115449 -51681 115505 -51637
rect 115549 -51681 115605 -51637
rect 115649 -51681 115705 -51637
rect 115749 -51681 115805 -51637
rect 115849 -51681 115905 -51637
rect 115949 -51681 116005 -51637
rect 116049 -51681 116105 -51637
rect 116149 -51681 116205 -51637
rect 116249 -51681 116305 -51637
rect 116349 -51681 116405 -51637
rect 116449 -51681 116505 -51637
rect 116549 -51681 116605 -51637
rect 116649 -51681 116705 -51637
rect 116749 -51681 116805 -51637
rect 116849 -51681 117196 -51637
rect 108496 -51737 117196 -51681
rect 108496 -51781 109305 -51737
rect 109349 -51781 109405 -51737
rect 109449 -51781 109505 -51737
rect 109549 -51781 109605 -51737
rect 109649 -51781 109705 -51737
rect 109749 -51781 109805 -51737
rect 109849 -51781 109905 -51737
rect 109949 -51781 110005 -51737
rect 110049 -51781 110105 -51737
rect 110149 -51781 110205 -51737
rect 110249 -51781 110305 -51737
rect 110349 -51781 110405 -51737
rect 110449 -51781 110505 -51737
rect 110549 -51781 110605 -51737
rect 110649 -51781 110705 -51737
rect 110749 -51781 110805 -51737
rect 110849 -51781 111305 -51737
rect 111349 -51781 111405 -51737
rect 111449 -51781 111505 -51737
rect 111549 -51781 111605 -51737
rect 111649 -51781 111705 -51737
rect 111749 -51781 111805 -51737
rect 111849 -51781 111905 -51737
rect 111949 -51781 112005 -51737
rect 112049 -51781 112105 -51737
rect 112149 -51781 112205 -51737
rect 112249 -51781 112305 -51737
rect 112349 -51781 112405 -51737
rect 112449 -51781 112505 -51737
rect 112549 -51781 112605 -51737
rect 112649 -51781 112705 -51737
rect 112749 -51781 112805 -51737
rect 112849 -51781 113305 -51737
rect 113349 -51781 113405 -51737
rect 113449 -51781 113505 -51737
rect 113549 -51781 113605 -51737
rect 113649 -51781 113705 -51737
rect 113749 -51781 113805 -51737
rect 113849 -51781 113905 -51737
rect 113949 -51781 114005 -51737
rect 114049 -51781 114105 -51737
rect 114149 -51781 114205 -51737
rect 114249 -51781 114305 -51737
rect 114349 -51781 114405 -51737
rect 114449 -51781 114505 -51737
rect 114549 -51781 114605 -51737
rect 114649 -51781 114705 -51737
rect 114749 -51781 114805 -51737
rect 114849 -51781 115305 -51737
rect 115349 -51781 115405 -51737
rect 115449 -51781 115505 -51737
rect 115549 -51781 115605 -51737
rect 115649 -51781 115705 -51737
rect 115749 -51781 115805 -51737
rect 115849 -51781 115905 -51737
rect 115949 -51781 116005 -51737
rect 116049 -51781 116105 -51737
rect 116149 -51781 116205 -51737
rect 116249 -51781 116305 -51737
rect 116349 -51781 116405 -51737
rect 116449 -51781 116505 -51737
rect 116549 -51781 116605 -51737
rect 116649 -51781 116705 -51737
rect 116749 -51781 116805 -51737
rect 116849 -51781 117196 -51737
rect 108496 -51837 117196 -51781
rect 108496 -51881 109305 -51837
rect 109349 -51881 109405 -51837
rect 109449 -51881 109505 -51837
rect 109549 -51881 109605 -51837
rect 109649 -51881 109705 -51837
rect 109749 -51881 109805 -51837
rect 109849 -51881 109905 -51837
rect 109949 -51881 110005 -51837
rect 110049 -51881 110105 -51837
rect 110149 -51881 110205 -51837
rect 110249 -51881 110305 -51837
rect 110349 -51881 110405 -51837
rect 110449 -51881 110505 -51837
rect 110549 -51881 110605 -51837
rect 110649 -51881 110705 -51837
rect 110749 -51881 110805 -51837
rect 110849 -51881 111305 -51837
rect 111349 -51881 111405 -51837
rect 111449 -51881 111505 -51837
rect 111549 -51881 111605 -51837
rect 111649 -51881 111705 -51837
rect 111749 -51881 111805 -51837
rect 111849 -51881 111905 -51837
rect 111949 -51881 112005 -51837
rect 112049 -51881 112105 -51837
rect 112149 -51881 112205 -51837
rect 112249 -51881 112305 -51837
rect 112349 -51881 112405 -51837
rect 112449 -51881 112505 -51837
rect 112549 -51881 112605 -51837
rect 112649 -51881 112705 -51837
rect 112749 -51881 112805 -51837
rect 112849 -51881 113305 -51837
rect 113349 -51881 113405 -51837
rect 113449 -51881 113505 -51837
rect 113549 -51881 113605 -51837
rect 113649 -51881 113705 -51837
rect 113749 -51881 113805 -51837
rect 113849 -51881 113905 -51837
rect 113949 -51881 114005 -51837
rect 114049 -51881 114105 -51837
rect 114149 -51881 114205 -51837
rect 114249 -51881 114305 -51837
rect 114349 -51881 114405 -51837
rect 114449 -51881 114505 -51837
rect 114549 -51881 114605 -51837
rect 114649 -51881 114705 -51837
rect 114749 -51881 114805 -51837
rect 114849 -51881 115305 -51837
rect 115349 -51881 115405 -51837
rect 115449 -51881 115505 -51837
rect 115549 -51881 115605 -51837
rect 115649 -51881 115705 -51837
rect 115749 -51881 115805 -51837
rect 115849 -51881 115905 -51837
rect 115949 -51881 116005 -51837
rect 116049 -51881 116105 -51837
rect 116149 -51881 116205 -51837
rect 116249 -51881 116305 -51837
rect 116349 -51881 116405 -51837
rect 116449 -51881 116505 -51837
rect 116549 -51881 116605 -51837
rect 116649 -51881 116705 -51837
rect 116749 -51881 116805 -51837
rect 116849 -51881 117196 -51837
rect 108496 -51937 117196 -51881
rect 108496 -51981 109305 -51937
rect 109349 -51981 109405 -51937
rect 109449 -51981 109505 -51937
rect 109549 -51981 109605 -51937
rect 109649 -51981 109705 -51937
rect 109749 -51981 109805 -51937
rect 109849 -51981 109905 -51937
rect 109949 -51981 110005 -51937
rect 110049 -51981 110105 -51937
rect 110149 -51981 110205 -51937
rect 110249 -51981 110305 -51937
rect 110349 -51981 110405 -51937
rect 110449 -51981 110505 -51937
rect 110549 -51981 110605 -51937
rect 110649 -51981 110705 -51937
rect 110749 -51981 110805 -51937
rect 110849 -51981 111305 -51937
rect 111349 -51981 111405 -51937
rect 111449 -51981 111505 -51937
rect 111549 -51981 111605 -51937
rect 111649 -51981 111705 -51937
rect 111749 -51981 111805 -51937
rect 111849 -51981 111905 -51937
rect 111949 -51981 112005 -51937
rect 112049 -51981 112105 -51937
rect 112149 -51981 112205 -51937
rect 112249 -51981 112305 -51937
rect 112349 -51981 112405 -51937
rect 112449 -51981 112505 -51937
rect 112549 -51981 112605 -51937
rect 112649 -51981 112705 -51937
rect 112749 -51981 112805 -51937
rect 112849 -51981 113305 -51937
rect 113349 -51981 113405 -51937
rect 113449 -51981 113505 -51937
rect 113549 -51981 113605 -51937
rect 113649 -51981 113705 -51937
rect 113749 -51981 113805 -51937
rect 113849 -51981 113905 -51937
rect 113949 -51981 114005 -51937
rect 114049 -51981 114105 -51937
rect 114149 -51981 114205 -51937
rect 114249 -51981 114305 -51937
rect 114349 -51981 114405 -51937
rect 114449 -51981 114505 -51937
rect 114549 -51981 114605 -51937
rect 114649 -51981 114705 -51937
rect 114749 -51981 114805 -51937
rect 114849 -51981 115305 -51937
rect 115349 -51981 115405 -51937
rect 115449 -51981 115505 -51937
rect 115549 -51981 115605 -51937
rect 115649 -51981 115705 -51937
rect 115749 -51981 115805 -51937
rect 115849 -51981 115905 -51937
rect 115949 -51981 116005 -51937
rect 116049 -51981 116105 -51937
rect 116149 -51981 116205 -51937
rect 116249 -51981 116305 -51937
rect 116349 -51981 116405 -51937
rect 116449 -51981 116505 -51937
rect 116549 -51981 116605 -51937
rect 116649 -51981 116705 -51937
rect 116749 -51981 116805 -51937
rect 116849 -51981 117196 -51937
rect 108496 -52037 117196 -51981
rect 108496 -52081 109305 -52037
rect 109349 -52081 109405 -52037
rect 109449 -52081 109505 -52037
rect 109549 -52081 109605 -52037
rect 109649 -52081 109705 -52037
rect 109749 -52081 109805 -52037
rect 109849 -52081 109905 -52037
rect 109949 -52081 110005 -52037
rect 110049 -52081 110105 -52037
rect 110149 -52081 110205 -52037
rect 110249 -52081 110305 -52037
rect 110349 -52081 110405 -52037
rect 110449 -52081 110505 -52037
rect 110549 -52081 110605 -52037
rect 110649 -52081 110705 -52037
rect 110749 -52081 110805 -52037
rect 110849 -52081 111305 -52037
rect 111349 -52081 111405 -52037
rect 111449 -52081 111505 -52037
rect 111549 -52081 111605 -52037
rect 111649 -52081 111705 -52037
rect 111749 -52081 111805 -52037
rect 111849 -52081 111905 -52037
rect 111949 -52081 112005 -52037
rect 112049 -52081 112105 -52037
rect 112149 -52081 112205 -52037
rect 112249 -52081 112305 -52037
rect 112349 -52081 112405 -52037
rect 112449 -52081 112505 -52037
rect 112549 -52081 112605 -52037
rect 112649 -52081 112705 -52037
rect 112749 -52081 112805 -52037
rect 112849 -52081 113305 -52037
rect 113349 -52081 113405 -52037
rect 113449 -52081 113505 -52037
rect 113549 -52081 113605 -52037
rect 113649 -52081 113705 -52037
rect 113749 -52081 113805 -52037
rect 113849 -52081 113905 -52037
rect 113949 -52081 114005 -52037
rect 114049 -52081 114105 -52037
rect 114149 -52081 114205 -52037
rect 114249 -52081 114305 -52037
rect 114349 -52081 114405 -52037
rect 114449 -52081 114505 -52037
rect 114549 -52081 114605 -52037
rect 114649 -52081 114705 -52037
rect 114749 -52081 114805 -52037
rect 114849 -52081 115305 -52037
rect 115349 -52081 115405 -52037
rect 115449 -52081 115505 -52037
rect 115549 -52081 115605 -52037
rect 115649 -52081 115705 -52037
rect 115749 -52081 115805 -52037
rect 115849 -52081 115905 -52037
rect 115949 -52081 116005 -52037
rect 116049 -52081 116105 -52037
rect 116149 -52081 116205 -52037
rect 116249 -52081 116305 -52037
rect 116349 -52081 116405 -52037
rect 116449 -52081 116505 -52037
rect 116549 -52081 116605 -52037
rect 116649 -52081 116705 -52037
rect 116749 -52081 116805 -52037
rect 116849 -52081 117196 -52037
rect 108496 -52137 117196 -52081
rect 108496 -52181 109305 -52137
rect 109349 -52181 109405 -52137
rect 109449 -52181 109505 -52137
rect 109549 -52181 109605 -52137
rect 109649 -52181 109705 -52137
rect 109749 -52181 109805 -52137
rect 109849 -52181 109905 -52137
rect 109949 -52181 110005 -52137
rect 110049 -52181 110105 -52137
rect 110149 -52181 110205 -52137
rect 110249 -52181 110305 -52137
rect 110349 -52181 110405 -52137
rect 110449 -52181 110505 -52137
rect 110549 -52181 110605 -52137
rect 110649 -52181 110705 -52137
rect 110749 -52181 110805 -52137
rect 110849 -52181 111305 -52137
rect 111349 -52181 111405 -52137
rect 111449 -52181 111505 -52137
rect 111549 -52181 111605 -52137
rect 111649 -52181 111705 -52137
rect 111749 -52181 111805 -52137
rect 111849 -52181 111905 -52137
rect 111949 -52181 112005 -52137
rect 112049 -52181 112105 -52137
rect 112149 -52181 112205 -52137
rect 112249 -52181 112305 -52137
rect 112349 -52181 112405 -52137
rect 112449 -52181 112505 -52137
rect 112549 -52181 112605 -52137
rect 112649 -52181 112705 -52137
rect 112749 -52181 112805 -52137
rect 112849 -52181 113305 -52137
rect 113349 -52181 113405 -52137
rect 113449 -52181 113505 -52137
rect 113549 -52181 113605 -52137
rect 113649 -52181 113705 -52137
rect 113749 -52181 113805 -52137
rect 113849 -52181 113905 -52137
rect 113949 -52181 114005 -52137
rect 114049 -52181 114105 -52137
rect 114149 -52181 114205 -52137
rect 114249 -52181 114305 -52137
rect 114349 -52181 114405 -52137
rect 114449 -52181 114505 -52137
rect 114549 -52181 114605 -52137
rect 114649 -52181 114705 -52137
rect 114749 -52181 114805 -52137
rect 114849 -52181 115305 -52137
rect 115349 -52181 115405 -52137
rect 115449 -52181 115505 -52137
rect 115549 -52181 115605 -52137
rect 115649 -52181 115705 -52137
rect 115749 -52181 115805 -52137
rect 115849 -52181 115905 -52137
rect 115949 -52181 116005 -52137
rect 116049 -52181 116105 -52137
rect 116149 -52181 116205 -52137
rect 116249 -52181 116305 -52137
rect 116349 -52181 116405 -52137
rect 116449 -52181 116505 -52137
rect 116549 -52181 116605 -52137
rect 116649 -52181 116705 -52137
rect 116749 -52181 116805 -52137
rect 116849 -52181 117196 -52137
rect 108496 -52237 117196 -52181
rect 108496 -52281 109305 -52237
rect 109349 -52281 109405 -52237
rect 109449 -52281 109505 -52237
rect 109549 -52281 109605 -52237
rect 109649 -52281 109705 -52237
rect 109749 -52281 109805 -52237
rect 109849 -52281 109905 -52237
rect 109949 -52281 110005 -52237
rect 110049 -52281 110105 -52237
rect 110149 -52281 110205 -52237
rect 110249 -52281 110305 -52237
rect 110349 -52281 110405 -52237
rect 110449 -52281 110505 -52237
rect 110549 -52281 110605 -52237
rect 110649 -52281 110705 -52237
rect 110749 -52281 110805 -52237
rect 110849 -52281 111305 -52237
rect 111349 -52281 111405 -52237
rect 111449 -52281 111505 -52237
rect 111549 -52281 111605 -52237
rect 111649 -52281 111705 -52237
rect 111749 -52281 111805 -52237
rect 111849 -52281 111905 -52237
rect 111949 -52281 112005 -52237
rect 112049 -52281 112105 -52237
rect 112149 -52281 112205 -52237
rect 112249 -52281 112305 -52237
rect 112349 -52281 112405 -52237
rect 112449 -52281 112505 -52237
rect 112549 -52281 112605 -52237
rect 112649 -52281 112705 -52237
rect 112749 -52281 112805 -52237
rect 112849 -52281 113305 -52237
rect 113349 -52281 113405 -52237
rect 113449 -52281 113505 -52237
rect 113549 -52281 113605 -52237
rect 113649 -52281 113705 -52237
rect 113749 -52281 113805 -52237
rect 113849 -52281 113905 -52237
rect 113949 -52281 114005 -52237
rect 114049 -52281 114105 -52237
rect 114149 -52281 114205 -52237
rect 114249 -52281 114305 -52237
rect 114349 -52281 114405 -52237
rect 114449 -52281 114505 -52237
rect 114549 -52281 114605 -52237
rect 114649 -52281 114705 -52237
rect 114749 -52281 114805 -52237
rect 114849 -52281 115305 -52237
rect 115349 -52281 115405 -52237
rect 115449 -52281 115505 -52237
rect 115549 -52281 115605 -52237
rect 115649 -52281 115705 -52237
rect 115749 -52281 115805 -52237
rect 115849 -52281 115905 -52237
rect 115949 -52281 116005 -52237
rect 116049 -52281 116105 -52237
rect 116149 -52281 116205 -52237
rect 116249 -52281 116305 -52237
rect 116349 -52281 116405 -52237
rect 116449 -52281 116505 -52237
rect 116549 -52281 116605 -52237
rect 116649 -52281 116705 -52237
rect 116749 -52281 116805 -52237
rect 116849 -52281 117196 -52237
rect 108496 -52337 117196 -52281
rect 108496 -52381 109305 -52337
rect 109349 -52381 109405 -52337
rect 109449 -52381 109505 -52337
rect 109549 -52381 109605 -52337
rect 109649 -52381 109705 -52337
rect 109749 -52381 109805 -52337
rect 109849 -52381 109905 -52337
rect 109949 -52381 110005 -52337
rect 110049 -52381 110105 -52337
rect 110149 -52381 110205 -52337
rect 110249 -52381 110305 -52337
rect 110349 -52381 110405 -52337
rect 110449 -52381 110505 -52337
rect 110549 -52381 110605 -52337
rect 110649 -52381 110705 -52337
rect 110749 -52381 110805 -52337
rect 110849 -52381 111305 -52337
rect 111349 -52381 111405 -52337
rect 111449 -52381 111505 -52337
rect 111549 -52381 111605 -52337
rect 111649 -52381 111705 -52337
rect 111749 -52381 111805 -52337
rect 111849 -52381 111905 -52337
rect 111949 -52381 112005 -52337
rect 112049 -52381 112105 -52337
rect 112149 -52381 112205 -52337
rect 112249 -52381 112305 -52337
rect 112349 -52381 112405 -52337
rect 112449 -52381 112505 -52337
rect 112549 -52381 112605 -52337
rect 112649 -52381 112705 -52337
rect 112749 -52381 112805 -52337
rect 112849 -52381 113305 -52337
rect 113349 -52381 113405 -52337
rect 113449 -52381 113505 -52337
rect 113549 -52381 113605 -52337
rect 113649 -52381 113705 -52337
rect 113749 -52381 113805 -52337
rect 113849 -52381 113905 -52337
rect 113949 -52381 114005 -52337
rect 114049 -52381 114105 -52337
rect 114149 -52381 114205 -52337
rect 114249 -52381 114305 -52337
rect 114349 -52381 114405 -52337
rect 114449 -52381 114505 -52337
rect 114549 -52381 114605 -52337
rect 114649 -52381 114705 -52337
rect 114749 -52381 114805 -52337
rect 114849 -52381 115305 -52337
rect 115349 -52381 115405 -52337
rect 115449 -52381 115505 -52337
rect 115549 -52381 115605 -52337
rect 115649 -52381 115705 -52337
rect 115749 -52381 115805 -52337
rect 115849 -52381 115905 -52337
rect 115949 -52381 116005 -52337
rect 116049 -52381 116105 -52337
rect 116149 -52381 116205 -52337
rect 116249 -52381 116305 -52337
rect 116349 -52381 116405 -52337
rect 116449 -52381 116505 -52337
rect 116549 -52381 116605 -52337
rect 116649 -52381 116705 -52337
rect 116749 -52381 116805 -52337
rect 116849 -52381 117196 -52337
rect 108496 -52437 117196 -52381
rect 108496 -52481 109305 -52437
rect 109349 -52481 109405 -52437
rect 109449 -52481 109505 -52437
rect 109549 -52481 109605 -52437
rect 109649 -52481 109705 -52437
rect 109749 -52481 109805 -52437
rect 109849 -52481 109905 -52437
rect 109949 -52481 110005 -52437
rect 110049 -52481 110105 -52437
rect 110149 -52481 110205 -52437
rect 110249 -52481 110305 -52437
rect 110349 -52481 110405 -52437
rect 110449 -52481 110505 -52437
rect 110549 -52481 110605 -52437
rect 110649 -52481 110705 -52437
rect 110749 -52481 110805 -52437
rect 110849 -52481 111305 -52437
rect 111349 -52481 111405 -52437
rect 111449 -52481 111505 -52437
rect 111549 -52481 111605 -52437
rect 111649 -52481 111705 -52437
rect 111749 -52481 111805 -52437
rect 111849 -52481 111905 -52437
rect 111949 -52481 112005 -52437
rect 112049 -52481 112105 -52437
rect 112149 -52481 112205 -52437
rect 112249 -52481 112305 -52437
rect 112349 -52481 112405 -52437
rect 112449 -52481 112505 -52437
rect 112549 -52481 112605 -52437
rect 112649 -52481 112705 -52437
rect 112749 -52481 112805 -52437
rect 112849 -52481 113305 -52437
rect 113349 -52481 113405 -52437
rect 113449 -52481 113505 -52437
rect 113549 -52481 113605 -52437
rect 113649 -52481 113705 -52437
rect 113749 -52481 113805 -52437
rect 113849 -52481 113905 -52437
rect 113949 -52481 114005 -52437
rect 114049 -52481 114105 -52437
rect 114149 -52481 114205 -52437
rect 114249 -52481 114305 -52437
rect 114349 -52481 114405 -52437
rect 114449 -52481 114505 -52437
rect 114549 -52481 114605 -52437
rect 114649 -52481 114705 -52437
rect 114749 -52481 114805 -52437
rect 114849 -52481 115305 -52437
rect 115349 -52481 115405 -52437
rect 115449 -52481 115505 -52437
rect 115549 -52481 115605 -52437
rect 115649 -52481 115705 -52437
rect 115749 -52481 115805 -52437
rect 115849 -52481 115905 -52437
rect 115949 -52481 116005 -52437
rect 116049 -52481 116105 -52437
rect 116149 -52481 116205 -52437
rect 116249 -52481 116305 -52437
rect 116349 -52481 116405 -52437
rect 116449 -52481 116505 -52437
rect 116549 -52481 116605 -52437
rect 116649 -52481 116705 -52437
rect 116749 -52481 116805 -52437
rect 116849 -52481 117196 -52437
rect 108496 -52537 117196 -52481
rect 108496 -52581 109305 -52537
rect 109349 -52581 109405 -52537
rect 109449 -52581 109505 -52537
rect 109549 -52581 109605 -52537
rect 109649 -52581 109705 -52537
rect 109749 -52581 109805 -52537
rect 109849 -52581 109905 -52537
rect 109949 -52581 110005 -52537
rect 110049 -52581 110105 -52537
rect 110149 -52581 110205 -52537
rect 110249 -52581 110305 -52537
rect 110349 -52581 110405 -52537
rect 110449 -52581 110505 -52537
rect 110549 -52581 110605 -52537
rect 110649 -52581 110705 -52537
rect 110749 -52581 110805 -52537
rect 110849 -52581 111305 -52537
rect 111349 -52581 111405 -52537
rect 111449 -52581 111505 -52537
rect 111549 -52581 111605 -52537
rect 111649 -52581 111705 -52537
rect 111749 -52581 111805 -52537
rect 111849 -52581 111905 -52537
rect 111949 -52581 112005 -52537
rect 112049 -52581 112105 -52537
rect 112149 -52581 112205 -52537
rect 112249 -52581 112305 -52537
rect 112349 -52581 112405 -52537
rect 112449 -52581 112505 -52537
rect 112549 -52581 112605 -52537
rect 112649 -52581 112705 -52537
rect 112749 -52581 112805 -52537
rect 112849 -52581 113305 -52537
rect 113349 -52581 113405 -52537
rect 113449 -52581 113505 -52537
rect 113549 -52581 113605 -52537
rect 113649 -52581 113705 -52537
rect 113749 -52581 113805 -52537
rect 113849 -52581 113905 -52537
rect 113949 -52581 114005 -52537
rect 114049 -52581 114105 -52537
rect 114149 -52581 114205 -52537
rect 114249 -52581 114305 -52537
rect 114349 -52581 114405 -52537
rect 114449 -52581 114505 -52537
rect 114549 -52581 114605 -52537
rect 114649 -52581 114705 -52537
rect 114749 -52581 114805 -52537
rect 114849 -52581 115305 -52537
rect 115349 -52581 115405 -52537
rect 115449 -52581 115505 -52537
rect 115549 -52581 115605 -52537
rect 115649 -52581 115705 -52537
rect 115749 -52581 115805 -52537
rect 115849 -52581 115905 -52537
rect 115949 -52581 116005 -52537
rect 116049 -52581 116105 -52537
rect 116149 -52581 116205 -52537
rect 116249 -52581 116305 -52537
rect 116349 -52581 116405 -52537
rect 116449 -52581 116505 -52537
rect 116549 -52581 116605 -52537
rect 116649 -52581 116705 -52537
rect 116749 -52581 116805 -52537
rect 116849 -52581 117196 -52537
rect 108496 -52636 117196 -52581
rect -109116 -52637 177360 -52636
rect -109116 -52681 109305 -52637
rect 109349 -52681 109405 -52637
rect 109449 -52681 109505 -52637
rect 109549 -52681 109605 -52637
rect 109649 -52681 109705 -52637
rect 109749 -52681 109805 -52637
rect 109849 -52681 109905 -52637
rect 109949 -52681 110005 -52637
rect 110049 -52681 110105 -52637
rect 110149 -52681 110205 -52637
rect 110249 -52681 110305 -52637
rect 110349 -52681 110405 -52637
rect 110449 -52681 110505 -52637
rect 110549 -52681 110605 -52637
rect 110649 -52681 110705 -52637
rect 110749 -52681 110805 -52637
rect 110849 -52681 111305 -52637
rect 111349 -52681 111405 -52637
rect 111449 -52681 111505 -52637
rect 111549 -52681 111605 -52637
rect 111649 -52681 111705 -52637
rect 111749 -52681 111805 -52637
rect 111849 -52681 111905 -52637
rect 111949 -52681 112005 -52637
rect 112049 -52681 112105 -52637
rect 112149 -52681 112205 -52637
rect 112249 -52681 112305 -52637
rect 112349 -52681 112405 -52637
rect 112449 -52681 112505 -52637
rect 112549 -52681 112605 -52637
rect 112649 -52681 112705 -52637
rect 112749 -52681 112805 -52637
rect 112849 -52681 113305 -52637
rect 113349 -52681 113405 -52637
rect 113449 -52681 113505 -52637
rect 113549 -52681 113605 -52637
rect 113649 -52681 113705 -52637
rect 113749 -52681 113805 -52637
rect 113849 -52681 113905 -52637
rect 113949 -52681 114005 -52637
rect 114049 -52681 114105 -52637
rect 114149 -52681 114205 -52637
rect 114249 -52681 114305 -52637
rect 114349 -52681 114405 -52637
rect 114449 -52681 114505 -52637
rect 114549 -52681 114605 -52637
rect 114649 -52681 114705 -52637
rect 114749 -52681 114805 -52637
rect 114849 -52681 115305 -52637
rect 115349 -52681 115405 -52637
rect 115449 -52681 115505 -52637
rect 115549 -52681 115605 -52637
rect 115649 -52681 115705 -52637
rect 115749 -52681 115805 -52637
rect 115849 -52681 115905 -52637
rect 115949 -52681 116005 -52637
rect 116049 -52681 116105 -52637
rect 116149 -52681 116205 -52637
rect 116249 -52681 116305 -52637
rect 116349 -52681 116405 -52637
rect 116449 -52681 116505 -52637
rect 116549 -52681 116605 -52637
rect 116649 -52681 116705 -52637
rect 116749 -52681 116805 -52637
rect 116849 -52681 177360 -52637
rect -109116 -53203 177360 -52681
rect -109116 -54117 -109040 -53203
rect -108508 -54117 -108432 -53203
rect -107900 -54117 -107824 -53203
rect -107292 -54117 -107216 -53203
rect -106684 -54117 -106608 -53203
rect -106076 -54117 -106000 -53203
rect -105468 -54117 -105392 -53203
rect -104860 -54117 -104784 -53203
rect -104252 -54117 -104176 -53203
rect -103644 -54117 -103568 -53203
rect -103036 -54117 -102960 -53203
rect -102428 -54117 -102352 -53203
rect -101820 -54117 -101744 -53203
rect -101212 -54117 -101136 -53203
rect -100604 -54117 -100528 -53203
rect -99996 -54117 -99920 -53203
rect -99388 -54117 -99312 -53203
rect -98780 -54117 -98704 -53203
rect -98172 -54117 -98096 -53203
rect -97564 -54117 -97488 -53203
rect -96956 -54117 -96880 -53203
rect -96348 -54117 -96272 -53203
rect -95740 -54117 -95664 -53203
rect -95132 -54117 -95056 -53203
rect -94524 -54117 -94448 -53203
rect -93916 -54117 -93840 -53203
rect -93308 -54117 -93232 -53203
rect -92700 -54117 -92624 -53203
rect -92092 -54117 -92016 -53203
rect -91484 -54117 -91408 -53203
rect -90876 -54117 -90800 -53203
rect -90268 -54117 -90192 -53203
rect -89660 -54117 -89584 -53203
rect -89052 -54117 -88976 -53203
rect -88444 -54117 -88368 -53203
rect -87836 -54117 -87760 -53203
rect -87228 -54117 -87152 -53203
rect -86620 -54117 -86544 -53203
rect -86012 -54117 -85936 -53203
rect -85404 -54117 -85328 -53203
rect -84796 -54117 -84720 -53203
rect -84188 -54117 -84112 -53203
rect -83580 -54117 -83504 -53203
rect -82972 -54117 -82896 -53203
rect -82364 -54117 -82288 -53203
rect -81756 -54117 -81680 -53203
rect -81148 -54117 -81072 -53203
rect -80540 -54117 -80464 -53203
rect -79932 -54117 -79856 -53203
rect -79324 -54117 -79248 -53203
rect -78716 -54117 -78640 -53203
rect -77116 -54117 -77040 -53203
rect -76508 -54117 -76432 -53203
rect -75900 -54117 -75824 -53203
rect -75292 -54117 -75216 -53203
rect -74684 -54117 -74608 -53203
rect -74076 -54117 -74000 -53203
rect -73468 -54117 -73392 -53203
rect -72860 -54117 -72784 -53203
rect -72252 -54117 -72176 -53203
rect -71644 -54117 -71568 -53203
rect -71036 -54117 -70960 -53203
rect -70428 -54117 -70352 -53203
rect -69820 -54117 -69744 -53203
rect -69212 -54117 -69136 -53203
rect -68604 -54117 -68528 -53203
rect -67996 -54117 -67920 -53203
rect -67388 -54117 -67312 -53203
rect -66780 -54117 -66704 -53203
rect -66172 -54117 -66096 -53203
rect -65564 -54117 -65488 -53203
rect -64956 -54117 -64880 -53203
rect -64348 -54117 -64272 -53203
rect -63740 -54117 -63664 -53203
rect -63132 -54117 -63056 -53203
rect -62524 -54117 -62448 -53203
rect -61916 -54117 -61840 -53203
rect -61308 -54117 -61232 -53203
rect -60700 -54117 -60624 -53203
rect -60092 -54117 -60016 -53203
rect -59484 -54117 -59408 -53203
rect -58876 -54117 -58800 -53203
rect -58268 -54117 -58192 -53203
rect -57660 -54117 -57584 -53203
rect -57052 -54117 -56976 -53203
rect -56444 -54117 -56368 -53203
rect -55836 -54117 -55760 -53203
rect -55228 -54117 -55152 -53203
rect -54620 -54117 -54544 -53203
rect -54012 -54117 -53936 -53203
rect -53404 -54117 -53328 -53203
rect -52796 -54117 -52720 -53203
rect -52188 -54117 -52112 -53203
rect -51580 -54117 -51504 -53203
rect -50972 -54117 -50896 -53203
rect -50364 -54117 -50288 -53203
rect -49756 -54117 -49680 -53203
rect -49148 -54117 -49072 -53203
rect -48540 -54117 -48464 -53203
rect -47932 -54117 -47856 -53203
rect -47324 -54117 -47248 -53203
rect -46716 -54117 -46640 -53203
rect -45116 -54117 -45040 -53203
rect -44508 -54117 -44432 -53203
rect -43900 -54117 -43824 -53203
rect -43292 -54117 -43216 -53203
rect -42684 -54117 -42608 -53203
rect -42076 -54117 -42000 -53203
rect -41468 -54117 -41392 -53203
rect -40860 -54117 -40784 -53203
rect -40252 -54117 -40176 -53203
rect -39644 -54117 -39568 -53203
rect -39036 -54117 -38960 -53203
rect -38428 -54117 -38352 -53203
rect -37820 -54117 -37744 -53203
rect -37212 -54117 -37136 -53203
rect -36604 -54117 -36528 -53203
rect -35996 -54117 -35920 -53203
rect -35388 -54117 -35312 -53203
rect -34780 -54117 -34704 -53203
rect -34172 -54117 -34096 -53203
rect -33564 -54117 -33488 -53203
rect -32956 -54117 -32880 -53203
rect -32348 -54117 -32272 -53203
rect -31740 -54117 -31664 -53203
rect -31132 -54117 -31056 -53203
rect -30524 -54117 -30448 -53203
rect -29916 -54117 -29840 -53203
rect -29308 -54117 -29232 -53203
rect -28700 -54117 -28624 -53203
rect -28092 -54117 -28016 -53203
rect -27484 -54117 -27408 -53203
rect -26876 -54117 -26800 -53203
rect -26268 -54117 -26192 -53203
rect -25660 -54117 -25584 -53203
rect -25052 -54117 -24976 -53203
rect -24444 -54117 -24368 -53203
rect -23836 -54117 -23760 -53203
rect -23228 -54117 -23152 -53203
rect -22620 -54117 -22544 -53203
rect -22012 -54117 -21936 -53203
rect -21404 -54117 -21328 -53203
rect -20796 -54117 -20720 -53203
rect -20188 -54117 -20112 -53203
rect -19580 -54117 -19504 -53203
rect -18972 -54117 -18896 -53203
rect -18364 -54117 -18288 -53203
rect -17756 -54117 -17680 -53203
rect -17148 -54117 -17072 -53203
rect -16540 -54117 -16464 -53203
rect -15932 -54117 -15856 -53203
rect -15324 -54117 -15248 -53203
rect -14716 -54117 -14640 -53203
rect -13116 -54117 -13040 -53203
rect -12508 -54117 -12432 -53203
rect -11900 -54117 -11824 -53203
rect -11292 -54117 -11216 -53203
rect -10684 -54117 -10608 -53203
rect -10076 -54117 -10000 -53203
rect -9468 -54117 -9392 -53203
rect -8860 -54117 -8784 -53203
rect -8252 -54117 -8176 -53203
rect -7644 -54117 -7568 -53203
rect -7036 -54117 -6960 -53203
rect -6428 -54117 -6352 -53203
rect -5820 -54117 -5744 -53203
rect -5212 -54117 -5136 -53203
rect -4604 -54117 -4528 -53203
rect -3996 -54117 -3920 -53203
rect -3388 -54117 -3312 -53203
rect -2780 -54117 -2704 -53203
rect -2172 -54117 -2096 -53203
rect -1564 -54117 -1488 -53203
rect -956 -54117 -880 -53203
rect -348 -54117 -272 -53203
rect 260 -54117 336 -53203
rect 868 -54117 944 -53203
rect 1476 -54117 1552 -53203
rect 2084 -54117 2160 -53203
rect 2692 -54117 2768 -53203
rect 3300 -54117 3376 -53203
rect 3908 -54117 3984 -53203
rect 4516 -54117 4592 -53203
rect 5124 -54117 5200 -53203
rect 5732 -54117 5808 -53203
rect 6340 -54117 6416 -53203
rect 6948 -54117 7024 -53203
rect 7556 -54117 7632 -53203
rect 8164 -54117 8240 -53203
rect 8772 -54117 8848 -53203
rect 9380 -54117 9456 -53203
rect 9988 -54117 10064 -53203
rect 10596 -54117 10672 -53203
rect 11204 -54117 11280 -53203
rect 11812 -54117 11888 -53203
rect 12420 -54117 12496 -53203
rect 13028 -54117 13104 -53203
rect 13636 -54117 13712 -53203
rect 14244 -54117 14320 -53203
rect 14852 -54117 14928 -53203
rect 15460 -54117 15536 -53203
rect 16068 -54117 16144 -53203
rect 16676 -54117 16752 -53203
rect 17284 -54117 17360 -53203
rect 18884 -54117 18960 -53203
rect 19492 -54117 19568 -53203
rect 20100 -54117 20176 -53203
rect 20708 -54117 20784 -53203
rect 21316 -54117 21392 -53203
rect 21924 -54117 22000 -53203
rect 22532 -54117 22608 -53203
rect 23140 -54117 23216 -53203
rect 23748 -54117 23824 -53203
rect 24356 -54117 24432 -53203
rect 24964 -54117 25040 -53203
rect 25572 -54117 25648 -53203
rect 26180 -54117 26256 -53203
rect 26788 -54117 26864 -53203
rect 27396 -54117 27472 -53203
rect 28004 -54117 28080 -53203
rect 28612 -54117 28688 -53203
rect 29220 -54117 29296 -53203
rect 29828 -54117 29904 -53203
rect 30436 -54117 30512 -53203
rect 31044 -54117 31120 -53203
rect 31652 -54117 31728 -53203
rect 32260 -54117 32336 -53203
rect 32868 -54117 32944 -53203
rect 33476 -54117 33552 -53203
rect 34084 -54117 34160 -53203
rect 34692 -54117 34768 -53203
rect 35300 -54117 35376 -53203
rect 35908 -54117 35984 -53203
rect 36516 -54117 36592 -53203
rect 37124 -54117 37200 -53203
rect 37732 -54117 37808 -53203
rect 38340 -54117 38416 -53203
rect 38948 -54117 39024 -53203
rect 39556 -54117 39632 -53203
rect 40164 -54117 40240 -53203
rect 40772 -54117 40848 -53203
rect 41380 -54117 41456 -53203
rect 41988 -54117 42064 -53203
rect 42596 -54117 42672 -53203
rect 43204 -54117 43280 -53203
rect 43812 -54117 43888 -53203
rect 44420 -54117 44496 -53203
rect 45028 -54117 45104 -53203
rect 45636 -54117 45712 -53203
rect 46244 -54117 46320 -53203
rect 46852 -54117 46928 -53203
rect 47460 -54117 47536 -53203
rect 48068 -54117 48144 -53203
rect 48676 -54117 48752 -53203
rect 49284 -54117 49360 -53203
rect 50884 -54117 50960 -53203
rect 51492 -54117 51568 -53203
rect 52100 -54117 52176 -53203
rect 52708 -54117 52784 -53203
rect 53316 -54117 53392 -53203
rect 53924 -54117 54000 -53203
rect 54532 -54117 54608 -53203
rect 55140 -54117 55216 -53203
rect 55748 -54117 55824 -53203
rect 56356 -54117 56432 -53203
rect 56964 -54117 57040 -53203
rect 57572 -54117 57648 -53203
rect 58180 -54117 58256 -53203
rect 58788 -54117 58864 -53203
rect 59396 -54117 59472 -53203
rect 60004 -54117 60080 -53203
rect 60612 -54117 60688 -53203
rect 61220 -54117 61296 -53203
rect 61828 -54117 61904 -53203
rect 62436 -54117 62512 -53203
rect 63044 -54117 63120 -53203
rect 63652 -54117 63728 -53203
rect 64260 -54117 64336 -53203
rect 64868 -54117 64944 -53203
rect 65476 -54117 65552 -53203
rect 66084 -54117 66160 -53203
rect 66692 -54117 66768 -53203
rect 67300 -54117 67376 -53203
rect 67908 -54117 67984 -53203
rect 68516 -54117 68592 -53203
rect 69124 -54117 69200 -53203
rect 69732 -54117 69808 -53203
rect 70340 -54117 70416 -53203
rect 70948 -54117 71024 -53203
rect 71556 -54117 71632 -53203
rect 72164 -54117 72240 -53203
rect 72772 -54117 72848 -53203
rect 73380 -54117 73456 -53203
rect 73988 -54117 74064 -53203
rect 74596 -54117 74672 -53203
rect 75204 -54117 75280 -53203
rect 75812 -54117 75888 -53203
rect 76420 -54117 76496 -53203
rect 77028 -54117 77104 -53203
rect 77636 -54117 77712 -53203
rect 78244 -54117 78320 -53203
rect 78852 -54117 78928 -53203
rect 79460 -54117 79536 -53203
rect 80068 -54117 80144 -53203
rect 80676 -54117 80752 -53203
rect 81284 -54117 81360 -53203
rect 82884 -54117 82960 -53203
rect 83492 -54117 83568 -53203
rect 84100 -54117 84176 -53203
rect 84708 -54117 84784 -53203
rect 85316 -54117 85392 -53203
rect 85924 -54117 86000 -53203
rect 86532 -54117 86608 -53203
rect 87140 -54117 87216 -53203
rect 87748 -54117 87824 -53203
rect 88356 -54117 88432 -53203
rect 88964 -54117 89040 -53203
rect 89572 -54117 89648 -53203
rect 90180 -54117 90256 -53203
rect 90788 -54117 90864 -53203
rect 91396 -54117 91472 -53203
rect 92004 -54117 92080 -53203
rect 92612 -54117 92688 -53203
rect 93220 -54117 93296 -53203
rect 93828 -54117 93904 -53203
rect 94436 -54117 94512 -53203
rect 95044 -54117 95120 -53203
rect 95652 -54117 95728 -53203
rect 96260 -54117 96336 -53203
rect 96868 -54117 96944 -53203
rect 97476 -54117 97552 -53203
rect 98084 -54117 98160 -53203
rect 98692 -54117 98768 -53203
rect 99300 -54117 99376 -53203
rect 99908 -54117 99984 -53203
rect 100516 -54117 100592 -53203
rect 101124 -54117 101200 -53203
rect 101732 -54117 101808 -53203
rect 102340 -54117 102416 -53203
rect 102948 -54117 103024 -53203
rect 103556 -54117 103632 -53203
rect 104164 -54117 104240 -53203
rect 104772 -54117 104848 -53203
rect 105380 -54117 105456 -53203
rect 105988 -54117 106064 -53203
rect 106596 -54117 106672 -53203
rect 107204 -54117 107280 -53203
rect 107812 -54117 107888 -53203
rect 108420 -54117 108496 -53203
rect 109028 -54117 109104 -53203
rect 109636 -54117 109712 -53203
rect 110244 -54117 110320 -53203
rect 110852 -54117 110928 -53203
rect 111460 -54117 111536 -53203
rect 112068 -54117 112144 -53203
rect 112676 -54117 112752 -53203
rect 113284 -54117 113360 -53203
rect 114884 -54117 114960 -53203
rect 115492 -54117 115568 -53203
rect 116100 -54117 116176 -53203
rect 116708 -54117 116784 -53203
rect 117316 -54117 117392 -53203
rect 117924 -54117 118000 -53203
rect 118532 -54117 118608 -53203
rect 119140 -54117 119216 -53203
rect 119748 -54117 119824 -53203
rect 120356 -54117 120432 -53203
rect 120964 -54117 121040 -53203
rect 121572 -54117 121648 -53203
rect 122180 -54117 122256 -53203
rect 122788 -54117 122864 -53203
rect 123396 -54117 123472 -53203
rect 124004 -54117 124080 -53203
rect 124612 -54117 124688 -53203
rect 125220 -54117 125296 -53203
rect 125828 -54117 125904 -53203
rect 126436 -54117 126512 -53203
rect 127044 -54117 127120 -53203
rect 127652 -54117 127728 -53203
rect 128260 -54117 128336 -53203
rect 128868 -54117 128944 -53203
rect 129476 -54117 129552 -53203
rect 130084 -54117 130160 -53203
rect 130692 -54117 130768 -53203
rect 131300 -54117 131376 -53203
rect 131908 -54117 131984 -53203
rect 132516 -54117 132592 -53203
rect 133124 -54117 133200 -53203
rect 133732 -54117 133808 -53203
rect 134340 -54117 134416 -53203
rect 134948 -54117 135024 -53203
rect 135556 -54117 135632 -53203
rect 136164 -54117 136240 -53203
rect 136772 -54117 136848 -53203
rect 137380 -54117 137456 -53203
rect 137988 -54117 138064 -53203
rect 138596 -54117 138672 -53203
rect 139204 -54117 139280 -53203
rect 139812 -54117 139888 -53203
rect 140420 -54117 140496 -53203
rect 141028 -54117 141104 -53203
rect 141636 -54117 141712 -53203
rect 142244 -54117 142320 -53203
rect 142852 -54117 142928 -53203
rect 143460 -54117 143536 -53203
rect 144068 -54117 144144 -53203
rect 144676 -54117 144752 -53203
rect 145284 -54117 145360 -53203
rect 146884 -54117 146960 -53203
rect 147492 -54117 147568 -53203
rect 148100 -54117 148176 -53203
rect 148708 -54117 148784 -53203
rect 149316 -54117 149392 -53203
rect 149924 -54117 150000 -53203
rect 150532 -54117 150608 -53203
rect 151140 -54117 151216 -53203
rect 151748 -54117 151824 -53203
rect 152356 -54117 152432 -53203
rect 152964 -54117 153040 -53203
rect 153572 -54117 153648 -53203
rect 154180 -54117 154256 -53203
rect 154788 -54117 154864 -53203
rect 155396 -54117 155472 -53203
rect 156004 -54117 156080 -53203
rect 156612 -54117 156688 -53203
rect 157220 -54117 157296 -53203
rect 157828 -54117 157904 -53203
rect 158436 -54117 158512 -53203
rect 159044 -54117 159120 -53203
rect 159652 -54117 159728 -53203
rect 160260 -54117 160336 -53203
rect 160868 -54117 160944 -53203
rect 161476 -54117 161552 -53203
rect 162084 -54117 162160 -53203
rect 162692 -54117 162768 -53203
rect 163300 -54117 163376 -53203
rect 163908 -54117 163984 -53203
rect 164516 -54117 164592 -53203
rect 165124 -54117 165200 -53203
rect 165732 -54117 165808 -53203
rect 166340 -54117 166416 -53203
rect 166948 -54117 167024 -53203
rect 167556 -54117 167632 -53203
rect 168164 -54117 168240 -53203
rect 168772 -54117 168848 -53203
rect 169380 -54117 169456 -53203
rect 169988 -54117 170064 -53203
rect 170596 -54117 170672 -53203
rect 171204 -54117 171280 -53203
rect 171812 -54117 171888 -53203
rect 172420 -54117 172496 -53203
rect 173028 -54117 173104 -53203
rect 173636 -54117 173712 -53203
rect 174244 -54117 174320 -53203
rect 174852 -54117 174928 -53203
rect 175460 -54117 175536 -53203
rect 176068 -54117 176144 -53203
rect 176676 -54117 176752 -53203
rect 177284 -54117 177360 -53203
rect -77274 -74121 -77040 -54119
rect -45274 -74121 -45040 -54119
rect -13274 -74121 -13040 -54119
rect 18726 -74121 18960 -54119
rect 50726 -74121 50960 -54119
rect 82726 -74121 82960 -54119
rect 114726 -74121 114960 -54119
rect 146726 -74121 146960 -54119
rect -108812 -75035 -108736 -74121
rect -108204 -75035 -108128 -74121
rect -107596 -75035 -107520 -74121
rect -106988 -75035 -106912 -74121
rect -106380 -75035 -106304 -74121
rect -105772 -75035 -105696 -74121
rect -105164 -75035 -105088 -74121
rect -104556 -75035 -104480 -74121
rect -103948 -75035 -103872 -74121
rect -103340 -75035 -103264 -74121
rect -102732 -75035 -102656 -74121
rect -102124 -75035 -102048 -74121
rect -101516 -75035 -101440 -74121
rect -100908 -75035 -100832 -74121
rect -100300 -75035 -100224 -74121
rect -99692 -75035 -99616 -74121
rect -99084 -75035 -99008 -74121
rect -98476 -75035 -98400 -74121
rect -97868 -75035 -97792 -74121
rect -97260 -75035 -97184 -74121
rect -96652 -75035 -96576 -74121
rect -96044 -75035 -95968 -74121
rect -95436 -75035 -95360 -74121
rect -94828 -75035 -94752 -74121
rect -94220 -75035 -94144 -74121
rect -93612 -75035 -93536 -74121
rect -93004 -75035 -92928 -74121
rect -92396 -75035 -92320 -74121
rect -91788 -75035 -91712 -74121
rect -91180 -75035 -91104 -74121
rect -90572 -75035 -90496 -74121
rect -89964 -75035 -89888 -74121
rect -89356 -75035 -89280 -74121
rect -88748 -75035 -88672 -74121
rect -88140 -75035 -88064 -74121
rect -87532 -75035 -87456 -74121
rect -86924 -75035 -86848 -74121
rect -86316 -75035 -86240 -74121
rect -85708 -75035 -85632 -74121
rect -85100 -75035 -85024 -74121
rect -84492 -75035 -84416 -74121
rect -83884 -75035 -83808 -74121
rect -83276 -75035 -83200 -74121
rect -82668 -75035 -82592 -74121
rect -82060 -75035 -81984 -74121
rect -81452 -75035 -81376 -74121
rect -80844 -75035 -80768 -74121
rect -80236 -75035 -80160 -74121
rect -79628 -75035 -79552 -74121
rect -79020 -75035 -78944 -74121
rect -76812 -75035 -76736 -74121
rect -76204 -75035 -76128 -74121
rect -75596 -75035 -75520 -74121
rect -74988 -75035 -74912 -74121
rect -74380 -75035 -74304 -74121
rect -73772 -75035 -73696 -74121
rect -73164 -75035 -73088 -74121
rect -72556 -75035 -72480 -74121
rect -71948 -75035 -71872 -74121
rect -71340 -75035 -71264 -74121
rect -70732 -75035 -70656 -74121
rect -70124 -75035 -70048 -74121
rect -69516 -75035 -69440 -74121
rect -68908 -75035 -68832 -74121
rect -68300 -75035 -68224 -74121
rect -67692 -75035 -67616 -74121
rect -67084 -75035 -67008 -74121
rect -66476 -75035 -66400 -74121
rect -65868 -75035 -65792 -74121
rect -65260 -75035 -65184 -74121
rect -64652 -75035 -64576 -74121
rect -64044 -75035 -63968 -74121
rect -63436 -75035 -63360 -74121
rect -62828 -75035 -62752 -74121
rect -62220 -75035 -62144 -74121
rect -61612 -75035 -61536 -74121
rect -61004 -75035 -60928 -74121
rect -60396 -75035 -60320 -74121
rect -59788 -75035 -59712 -74121
rect -59180 -75035 -59104 -74121
rect -58572 -75035 -58496 -74121
rect -57964 -75035 -57888 -74121
rect -57356 -75035 -57280 -74121
rect -56748 -75035 -56672 -74121
rect -56140 -75035 -56064 -74121
rect -55532 -75035 -55456 -74121
rect -54924 -75035 -54848 -74121
rect -54316 -75035 -54240 -74121
rect -53708 -75035 -53632 -74121
rect -53100 -75035 -53024 -74121
rect -52492 -75035 -52416 -74121
rect -51884 -75035 -51808 -74121
rect -51276 -75035 -51200 -74121
rect -50668 -75035 -50592 -74121
rect -50060 -75035 -49984 -74121
rect -49452 -75035 -49376 -74121
rect -48844 -75035 -48768 -74121
rect -48236 -75035 -48160 -74121
rect -47628 -75035 -47552 -74121
rect -47020 -75035 -46944 -74121
rect -44812 -75035 -44736 -74121
rect -44204 -75035 -44128 -74121
rect -43596 -75035 -43520 -74121
rect -42988 -75035 -42912 -74121
rect -42380 -75035 -42304 -74121
rect -41772 -75035 -41696 -74121
rect -41164 -75035 -41088 -74121
rect -40556 -75035 -40480 -74121
rect -39948 -75035 -39872 -74121
rect -39340 -75035 -39264 -74121
rect -38732 -75035 -38656 -74121
rect -38124 -75035 -38048 -74121
rect -37516 -75035 -37440 -74121
rect -36908 -75035 -36832 -74121
rect -36300 -75035 -36224 -74121
rect -35692 -75035 -35616 -74121
rect -35084 -75035 -35008 -74121
rect -34476 -75035 -34400 -74121
rect -33868 -75035 -33792 -74121
rect -33260 -75035 -33184 -74121
rect -32652 -75035 -32576 -74121
rect -32044 -75035 -31968 -74121
rect -31436 -75035 -31360 -74121
rect -30828 -75035 -30752 -74121
rect -30220 -75035 -30144 -74121
rect -29612 -75035 -29536 -74121
rect -29004 -75035 -28928 -74121
rect -28396 -75035 -28320 -74121
rect -27788 -75035 -27712 -74121
rect -27180 -75035 -27104 -74121
rect -26572 -75035 -26496 -74121
rect -25964 -75035 -25888 -74121
rect -25356 -75035 -25280 -74121
rect -24748 -75035 -24672 -74121
rect -24140 -75035 -24064 -74121
rect -23532 -75035 -23456 -74121
rect -22924 -75035 -22848 -74121
rect -22316 -75035 -22240 -74121
rect -21708 -75035 -21632 -74121
rect -21100 -75035 -21024 -74121
rect -20492 -75035 -20416 -74121
rect -19884 -75035 -19808 -74121
rect -19276 -75035 -19200 -74121
rect -18668 -75035 -18592 -74121
rect -18060 -75035 -17984 -74121
rect -17452 -75035 -17376 -74121
rect -16844 -75035 -16768 -74121
rect -16236 -75035 -16160 -74121
rect -15628 -75035 -15552 -74121
rect -15020 -75035 -14944 -74121
rect -12812 -75035 -12736 -74121
rect -12204 -75035 -12128 -74121
rect -11596 -75035 -11520 -74121
rect -10988 -75035 -10912 -74121
rect -10380 -75035 -10304 -74121
rect -9772 -75035 -9696 -74121
rect -9164 -75035 -9088 -74121
rect -8556 -75035 -8480 -74121
rect -7948 -75035 -7872 -74121
rect -7340 -75035 -7264 -74121
rect -6732 -75035 -6656 -74121
rect -6124 -75035 -6048 -74121
rect -5516 -75035 -5440 -74121
rect -4908 -75035 -4832 -74121
rect -4300 -75035 -4224 -74121
rect -3692 -75035 -3616 -74121
rect -3084 -75035 -3008 -74121
rect -2476 -75035 -2400 -74121
rect -1868 -75035 -1792 -74121
rect -1260 -75035 -1184 -74121
rect -652 -75035 -576 -74121
rect -44 -75035 32 -74121
rect 564 -75035 640 -74121
rect 1172 -75035 1248 -74121
rect 1780 -75035 1856 -74121
rect 2388 -75035 2464 -74121
rect 2996 -75035 3072 -74121
rect 3604 -75035 3680 -74121
rect 4212 -75035 4288 -74121
rect 4820 -75035 4896 -74121
rect 5428 -75035 5504 -74121
rect 6036 -75035 6112 -74121
rect 6644 -75035 6720 -74121
rect 7252 -75035 7328 -74121
rect 7860 -75035 7936 -74121
rect 8468 -75035 8544 -74121
rect 9076 -75035 9152 -74121
rect 9684 -75035 9760 -74121
rect 10292 -75035 10368 -74121
rect 10900 -75035 10976 -74121
rect 11508 -75035 11584 -74121
rect 12116 -75035 12192 -74121
rect 12724 -75035 12800 -74121
rect 13332 -75035 13408 -74121
rect 13940 -75035 14016 -74121
rect 14548 -75035 14624 -74121
rect 15156 -75035 15232 -74121
rect 15764 -75035 15840 -74121
rect 16372 -75035 16448 -74121
rect 16980 -75035 17056 -74121
rect 19188 -75035 19264 -74121
rect 19796 -75035 19872 -74121
rect 20404 -75035 20480 -74121
rect 21012 -75035 21088 -74121
rect 21620 -75035 21696 -74121
rect 22228 -75035 22304 -74121
rect 22836 -75035 22912 -74121
rect 23444 -75035 23520 -74121
rect 24052 -75035 24128 -74121
rect 24660 -75035 24736 -74121
rect 25268 -75035 25344 -74121
rect 25876 -75035 25952 -74121
rect 26484 -75035 26560 -74121
rect 27092 -75035 27168 -74121
rect 27700 -75035 27776 -74121
rect 28308 -75035 28384 -74121
rect 28916 -75035 28992 -74121
rect 29524 -75035 29600 -74121
rect 30132 -75035 30208 -74121
rect 30740 -75035 30816 -74121
rect 31348 -75035 31424 -74121
rect 31956 -75035 32032 -74121
rect 32564 -75035 32640 -74121
rect 33172 -75035 33248 -74121
rect 33780 -75035 33856 -74121
rect 34388 -75035 34464 -74121
rect 34996 -75035 35072 -74121
rect 35604 -75035 35680 -74121
rect 36212 -75035 36288 -74121
rect 36820 -75035 36896 -74121
rect 37428 -75035 37504 -74121
rect 38036 -75035 38112 -74121
rect 38644 -75035 38720 -74121
rect 39252 -75035 39328 -74121
rect 39860 -75035 39936 -74121
rect 40468 -75035 40544 -74121
rect 41076 -75035 41152 -74121
rect 41684 -75035 41760 -74121
rect 42292 -75035 42368 -74121
rect 42900 -75035 42976 -74121
rect 43508 -75035 43584 -74121
rect 44116 -75035 44192 -74121
rect 44724 -75035 44800 -74121
rect 45332 -75035 45408 -74121
rect 45940 -75035 46016 -74121
rect 46548 -75035 46624 -74121
rect 47156 -75035 47232 -74121
rect 47764 -75035 47840 -74121
rect 48372 -75035 48448 -74121
rect 48980 -75035 49056 -74121
rect 51188 -75035 51264 -74121
rect 51796 -75035 51872 -74121
rect 52404 -75035 52480 -74121
rect 53012 -75035 53088 -74121
rect 53620 -75035 53696 -74121
rect 54228 -75035 54304 -74121
rect 54836 -75035 54912 -74121
rect 55444 -75035 55520 -74121
rect 56052 -75035 56128 -74121
rect 56660 -75035 56736 -74121
rect 57268 -75035 57344 -74121
rect 57876 -75035 57952 -74121
rect 58484 -75035 58560 -74121
rect 59092 -75035 59168 -74121
rect 59700 -75035 59776 -74121
rect 60308 -75035 60384 -74121
rect 60916 -75035 60992 -74121
rect 61524 -75035 61600 -74121
rect 62132 -75035 62208 -74121
rect 62740 -75035 62816 -74121
rect 63348 -75035 63424 -74121
rect 63956 -75035 64032 -74121
rect 64564 -75035 64640 -74121
rect 65172 -75035 65248 -74121
rect 65780 -75035 65856 -74121
rect 66388 -75035 66464 -74121
rect 66996 -75035 67072 -74121
rect 67604 -75035 67680 -74121
rect 68212 -75035 68288 -74121
rect 68820 -75035 68896 -74121
rect 69428 -75035 69504 -74121
rect 70036 -75035 70112 -74121
rect 70644 -75035 70720 -74121
rect 71252 -75035 71328 -74121
rect 71860 -75035 71936 -74121
rect 72468 -75035 72544 -74121
rect 73076 -75035 73152 -74121
rect 73684 -75035 73760 -74121
rect 74292 -75035 74368 -74121
rect 74900 -75035 74976 -74121
rect 75508 -75035 75584 -74121
rect 76116 -75035 76192 -74121
rect 76724 -75035 76800 -74121
rect 77332 -75035 77408 -74121
rect 77940 -75035 78016 -74121
rect 78548 -75035 78624 -74121
rect 79156 -75035 79232 -74121
rect 79764 -75035 79840 -74121
rect 80372 -75035 80448 -74121
rect 80980 -75035 81056 -74121
rect 83188 -75035 83264 -74121
rect 83796 -75035 83872 -74121
rect 84404 -75035 84480 -74121
rect 85012 -75035 85088 -74121
rect 85620 -75035 85696 -74121
rect 86228 -75035 86304 -74121
rect 86836 -75035 86912 -74121
rect 87444 -75035 87520 -74121
rect 88052 -75035 88128 -74121
rect 88660 -75035 88736 -74121
rect 89268 -75035 89344 -74121
rect 89876 -75035 89952 -74121
rect 90484 -75035 90560 -74121
rect 91092 -75035 91168 -74121
rect 91700 -75035 91776 -74121
rect 92308 -75035 92384 -74121
rect 92916 -75035 92992 -74121
rect 93524 -75035 93600 -74121
rect 94132 -75035 94208 -74121
rect 94740 -75035 94816 -74121
rect 95348 -75035 95424 -74121
rect 95956 -75035 96032 -74121
rect 96564 -75035 96640 -74121
rect 97172 -75035 97248 -74121
rect 97780 -75035 97856 -74121
rect 98388 -75035 98464 -74121
rect 98996 -75035 99072 -74121
rect 99604 -75035 99680 -74121
rect 100212 -75035 100288 -74121
rect 100820 -75035 100896 -74121
rect 101428 -75035 101504 -74121
rect 102036 -75035 102112 -74121
rect 102644 -75035 102720 -74121
rect 103252 -75035 103328 -74121
rect 103860 -75035 103936 -74121
rect 104468 -75035 104544 -74121
rect 105076 -75035 105152 -74121
rect 105684 -75035 105760 -74121
rect 106292 -75035 106368 -74121
rect 106900 -75035 106976 -74121
rect 107508 -75035 107584 -74121
rect 108116 -75035 108192 -74121
rect 108724 -75035 108800 -74121
rect 109332 -75035 109408 -74121
rect 109940 -75035 110016 -74121
rect 110548 -75035 110624 -74121
rect 111156 -75035 111232 -74121
rect 111764 -75035 111840 -74121
rect 112372 -75035 112448 -74121
rect 112980 -75035 113056 -74121
rect 115188 -75035 115264 -74121
rect 115796 -75035 115872 -74121
rect 116404 -75035 116480 -74121
rect 117012 -75035 117088 -74121
rect 117620 -75035 117696 -74121
rect 118228 -75035 118304 -74121
rect 118836 -75035 118912 -74121
rect 119444 -75035 119520 -74121
rect 120052 -75035 120128 -74121
rect 120660 -75035 120736 -74121
rect 121268 -75035 121344 -74121
rect 121876 -75035 121952 -74121
rect 122484 -75035 122560 -74121
rect 123092 -75035 123168 -74121
rect 123700 -75035 123776 -74121
rect 124308 -75035 124384 -74121
rect 124916 -75035 124992 -74121
rect 125524 -75035 125600 -74121
rect 126132 -75035 126208 -74121
rect 126740 -75035 126816 -74121
rect 127348 -75035 127424 -74121
rect 127956 -75035 128032 -74121
rect 128564 -75035 128640 -74121
rect 129172 -75035 129248 -74121
rect 129780 -75035 129856 -74121
rect 130388 -75035 130464 -74121
rect 130996 -75035 131072 -74121
rect 131604 -75035 131680 -74121
rect 132212 -75035 132288 -74121
rect 132820 -75035 132896 -74121
rect 133428 -75035 133504 -74121
rect 134036 -75035 134112 -74121
rect 134644 -75035 134720 -74121
rect 135252 -75035 135328 -74121
rect 135860 -75035 135936 -74121
rect 136468 -75035 136544 -74121
rect 137076 -75035 137152 -74121
rect 137684 -75035 137760 -74121
rect 138292 -75035 138368 -74121
rect 138900 -75035 138976 -74121
rect 139508 -75035 139584 -74121
rect 140116 -75035 140192 -74121
rect 140724 -75035 140800 -74121
rect 141332 -75035 141408 -74121
rect 141940 -75035 142016 -74121
rect 142548 -75035 142624 -74121
rect 143156 -75035 143232 -74121
rect 143764 -75035 143840 -74121
rect 144372 -75035 144448 -74121
rect 144980 -75035 145056 -74121
rect 147188 -75035 147264 -74121
rect 147796 -75035 147872 -74121
rect 148404 -75035 148480 -74121
rect 149012 -75035 149088 -74121
rect 149620 -75035 149696 -74121
rect 150228 -75035 150304 -74121
rect 150836 -75035 150912 -74121
rect 151444 -75035 151520 -74121
rect 152052 -75035 152128 -74121
rect 152660 -75035 152736 -74121
rect 153268 -75035 153344 -74121
rect 153876 -75035 153952 -74121
rect 154484 -75035 154560 -74121
rect 155092 -75035 155168 -74121
rect 155700 -75035 155776 -74121
rect 156308 -75035 156384 -74121
rect 156916 -75035 156992 -74121
rect 157524 -75035 157600 -74121
rect 158132 -75035 158208 -74121
rect 158740 -75035 158816 -74121
rect 159348 -75035 159424 -74121
rect 159956 -75035 160032 -74121
rect 160564 -75035 160640 -74121
rect 161172 -75035 161248 -74121
rect 161780 -75035 161856 -74121
rect 162388 -75035 162464 -74121
rect 162996 -75035 163072 -74121
rect 163604 -75035 163680 -74121
rect 164212 -75035 164288 -74121
rect 164820 -75035 164896 -74121
rect 165428 -75035 165504 -74121
rect 166036 -75035 166112 -74121
rect 166644 -75035 166720 -74121
rect 167252 -75035 167328 -74121
rect 167860 -75035 167936 -74121
rect 168468 -75035 168544 -74121
rect 169076 -75035 169152 -74121
rect 169684 -75035 169760 -74121
rect 170292 -75035 170368 -74121
rect 170900 -75035 170976 -74121
rect 171508 -75035 171584 -74121
rect 172116 -75035 172192 -74121
rect 172724 -75035 172800 -74121
rect 173332 -75035 173408 -74121
rect 173940 -75035 174016 -74121
rect 174548 -75035 174624 -74121
rect 175156 -75035 175232 -74121
rect 175764 -75035 175840 -74121
rect 176372 -75035 176448 -74121
rect 176980 -75035 177056 -74121
rect 177664 -75035 178308 -49602
rect -108812 -75188 178308 -75035
rect -108812 -75232 9236 -75188
rect 9280 -75232 9336 -75188
rect 9380 -75232 9436 -75188
rect 9480 -75232 9536 -75188
rect 9580 -75232 9636 -75188
rect 9680 -75232 9736 -75188
rect 9780 -75232 9836 -75188
rect 9880 -75232 9936 -75188
rect 9980 -75232 10036 -75188
rect 10080 -75232 10136 -75188
rect 10180 -75232 10236 -75188
rect 10280 -75232 10336 -75188
rect 10380 -75232 10436 -75188
rect 10480 -75232 10536 -75188
rect 10580 -75232 10636 -75188
rect 10680 -75232 10736 -75188
rect 10780 -75232 11236 -75188
rect 11280 -75232 11336 -75188
rect 11380 -75232 11436 -75188
rect 11480 -75232 11536 -75188
rect 11580 -75232 11636 -75188
rect 11680 -75232 11736 -75188
rect 11780 -75232 11836 -75188
rect 11880 -75232 11936 -75188
rect 11980 -75232 12036 -75188
rect 12080 -75232 12136 -75188
rect 12180 -75232 12236 -75188
rect 12280 -75232 12336 -75188
rect 12380 -75232 12436 -75188
rect 12480 -75232 12536 -75188
rect 12580 -75232 12636 -75188
rect 12680 -75232 12736 -75188
rect 12780 -75232 13236 -75188
rect 13280 -75232 13336 -75188
rect 13380 -75232 13436 -75188
rect 13480 -75232 13536 -75188
rect 13580 -75232 13636 -75188
rect 13680 -75232 13736 -75188
rect 13780 -75232 13836 -75188
rect 13880 -75232 13936 -75188
rect 13980 -75232 14036 -75188
rect 14080 -75232 14136 -75188
rect 14180 -75232 14236 -75188
rect 14280 -75232 14336 -75188
rect 14380 -75232 14436 -75188
rect 14480 -75232 14536 -75188
rect 14580 -75232 14636 -75188
rect 14680 -75232 14736 -75188
rect 14780 -75232 15236 -75188
rect 15280 -75232 15336 -75188
rect 15380 -75232 15436 -75188
rect 15480 -75232 15536 -75188
rect 15580 -75232 15636 -75188
rect 15680 -75232 15736 -75188
rect 15780 -75232 15836 -75188
rect 15880 -75232 15936 -75188
rect 15980 -75232 16036 -75188
rect 16080 -75232 16136 -75188
rect 16180 -75232 16236 -75188
rect 16280 -75232 16336 -75188
rect 16380 -75232 16436 -75188
rect 16480 -75232 16536 -75188
rect 16580 -75232 16636 -75188
rect 16680 -75232 16736 -75188
rect 16780 -75232 178308 -75188
rect -108812 -75288 178308 -75232
rect -108812 -75332 9236 -75288
rect 9280 -75332 9336 -75288
rect 9380 -75332 9436 -75288
rect 9480 -75332 9536 -75288
rect 9580 -75332 9636 -75288
rect 9680 -75332 9736 -75288
rect 9780 -75332 9836 -75288
rect 9880 -75332 9936 -75288
rect 9980 -75332 10036 -75288
rect 10080 -75332 10136 -75288
rect 10180 -75332 10236 -75288
rect 10280 -75332 10336 -75288
rect 10380 -75332 10436 -75288
rect 10480 -75332 10536 -75288
rect 10580 -75332 10636 -75288
rect 10680 -75332 10736 -75288
rect 10780 -75332 11236 -75288
rect 11280 -75332 11336 -75288
rect 11380 -75332 11436 -75288
rect 11480 -75332 11536 -75288
rect 11580 -75332 11636 -75288
rect 11680 -75332 11736 -75288
rect 11780 -75332 11836 -75288
rect 11880 -75332 11936 -75288
rect 11980 -75332 12036 -75288
rect 12080 -75332 12136 -75288
rect 12180 -75332 12236 -75288
rect 12280 -75332 12336 -75288
rect 12380 -75332 12436 -75288
rect 12480 -75332 12536 -75288
rect 12580 -75332 12636 -75288
rect 12680 -75332 12736 -75288
rect 12780 -75332 13236 -75288
rect 13280 -75332 13336 -75288
rect 13380 -75332 13436 -75288
rect 13480 -75332 13536 -75288
rect 13580 -75332 13636 -75288
rect 13680 -75332 13736 -75288
rect 13780 -75332 13836 -75288
rect 13880 -75332 13936 -75288
rect 13980 -75332 14036 -75288
rect 14080 -75332 14136 -75288
rect 14180 -75332 14236 -75288
rect 14280 -75332 14336 -75288
rect 14380 -75332 14436 -75288
rect 14480 -75332 14536 -75288
rect 14580 -75332 14636 -75288
rect 14680 -75332 14736 -75288
rect 14780 -75332 15236 -75288
rect 15280 -75332 15336 -75288
rect 15380 -75332 15436 -75288
rect 15480 -75332 15536 -75288
rect 15580 -75332 15636 -75288
rect 15680 -75332 15736 -75288
rect 15780 -75332 15836 -75288
rect 15880 -75332 15936 -75288
rect 15980 -75332 16036 -75288
rect 16080 -75332 16136 -75288
rect 16180 -75332 16236 -75288
rect 16280 -75332 16336 -75288
rect 16380 -75332 16436 -75288
rect 16480 -75332 16536 -75288
rect 16580 -75332 16636 -75288
rect 16680 -75332 16736 -75288
rect 16780 -75332 178308 -75288
rect -108812 -75388 178308 -75332
rect -108812 -75432 9236 -75388
rect 9280 -75432 9336 -75388
rect 9380 -75432 9436 -75388
rect 9480 -75432 9536 -75388
rect 9580 -75432 9636 -75388
rect 9680 -75432 9736 -75388
rect 9780 -75432 9836 -75388
rect 9880 -75432 9936 -75388
rect 9980 -75432 10036 -75388
rect 10080 -75432 10136 -75388
rect 10180 -75432 10236 -75388
rect 10280 -75432 10336 -75388
rect 10380 -75432 10436 -75388
rect 10480 -75432 10536 -75388
rect 10580 -75432 10636 -75388
rect 10680 -75432 10736 -75388
rect 10780 -75432 11236 -75388
rect 11280 -75432 11336 -75388
rect 11380 -75432 11436 -75388
rect 11480 -75432 11536 -75388
rect 11580 -75432 11636 -75388
rect 11680 -75432 11736 -75388
rect 11780 -75432 11836 -75388
rect 11880 -75432 11936 -75388
rect 11980 -75432 12036 -75388
rect 12080 -75432 12136 -75388
rect 12180 -75432 12236 -75388
rect 12280 -75432 12336 -75388
rect 12380 -75432 12436 -75388
rect 12480 -75432 12536 -75388
rect 12580 -75432 12636 -75388
rect 12680 -75432 12736 -75388
rect 12780 -75432 13236 -75388
rect 13280 -75432 13336 -75388
rect 13380 -75432 13436 -75388
rect 13480 -75432 13536 -75388
rect 13580 -75432 13636 -75388
rect 13680 -75432 13736 -75388
rect 13780 -75432 13836 -75388
rect 13880 -75432 13936 -75388
rect 13980 -75432 14036 -75388
rect 14080 -75432 14136 -75388
rect 14180 -75432 14236 -75388
rect 14280 -75432 14336 -75388
rect 14380 -75432 14436 -75388
rect 14480 -75432 14536 -75388
rect 14580 -75432 14636 -75388
rect 14680 -75432 14736 -75388
rect 14780 -75432 15236 -75388
rect 15280 -75432 15336 -75388
rect 15380 -75432 15436 -75388
rect 15480 -75432 15536 -75388
rect 15580 -75432 15636 -75388
rect 15680 -75432 15736 -75388
rect 15780 -75432 15836 -75388
rect 15880 -75432 15936 -75388
rect 15980 -75432 16036 -75388
rect 16080 -75432 16136 -75388
rect 16180 -75432 16236 -75388
rect 16280 -75432 16336 -75388
rect 16380 -75432 16436 -75388
rect 16480 -75432 16536 -75388
rect 16580 -75432 16636 -75388
rect 16680 -75432 16736 -75388
rect 16780 -75432 178308 -75388
rect -108812 -75488 178308 -75432
rect -108812 -75532 9236 -75488
rect 9280 -75532 9336 -75488
rect 9380 -75532 9436 -75488
rect 9480 -75532 9536 -75488
rect 9580 -75532 9636 -75488
rect 9680 -75532 9736 -75488
rect 9780 -75532 9836 -75488
rect 9880 -75532 9936 -75488
rect 9980 -75532 10036 -75488
rect 10080 -75532 10136 -75488
rect 10180 -75532 10236 -75488
rect 10280 -75532 10336 -75488
rect 10380 -75532 10436 -75488
rect 10480 -75532 10536 -75488
rect 10580 -75532 10636 -75488
rect 10680 -75532 10736 -75488
rect 10780 -75532 11236 -75488
rect 11280 -75532 11336 -75488
rect 11380 -75532 11436 -75488
rect 11480 -75532 11536 -75488
rect 11580 -75532 11636 -75488
rect 11680 -75532 11736 -75488
rect 11780 -75532 11836 -75488
rect 11880 -75532 11936 -75488
rect 11980 -75532 12036 -75488
rect 12080 -75532 12136 -75488
rect 12180 -75532 12236 -75488
rect 12280 -75532 12336 -75488
rect 12380 -75532 12436 -75488
rect 12480 -75532 12536 -75488
rect 12580 -75532 12636 -75488
rect 12680 -75532 12736 -75488
rect 12780 -75532 13236 -75488
rect 13280 -75532 13336 -75488
rect 13380 -75532 13436 -75488
rect 13480 -75532 13536 -75488
rect 13580 -75532 13636 -75488
rect 13680 -75532 13736 -75488
rect 13780 -75532 13836 -75488
rect 13880 -75532 13936 -75488
rect 13980 -75532 14036 -75488
rect 14080 -75532 14136 -75488
rect 14180 -75532 14236 -75488
rect 14280 -75532 14336 -75488
rect 14380 -75532 14436 -75488
rect 14480 -75532 14536 -75488
rect 14580 -75532 14636 -75488
rect 14680 -75532 14736 -75488
rect 14780 -75532 15236 -75488
rect 15280 -75532 15336 -75488
rect 15380 -75532 15436 -75488
rect 15480 -75532 15536 -75488
rect 15580 -75532 15636 -75488
rect 15680 -75532 15736 -75488
rect 15780 -75532 15836 -75488
rect 15880 -75532 15936 -75488
rect 15980 -75532 16036 -75488
rect 16080 -75532 16136 -75488
rect 16180 -75532 16236 -75488
rect 16280 -75532 16336 -75488
rect 16380 -75532 16436 -75488
rect 16480 -75532 16536 -75488
rect 16580 -75532 16636 -75488
rect 16680 -75532 16736 -75488
rect 16780 -75532 178308 -75488
rect -108812 -75588 178308 -75532
rect -108812 -75632 9236 -75588
rect 9280 -75632 9336 -75588
rect 9380 -75632 9436 -75588
rect 9480 -75632 9536 -75588
rect 9580 -75632 9636 -75588
rect 9680 -75632 9736 -75588
rect 9780 -75632 9836 -75588
rect 9880 -75632 9936 -75588
rect 9980 -75632 10036 -75588
rect 10080 -75632 10136 -75588
rect 10180 -75632 10236 -75588
rect 10280 -75632 10336 -75588
rect 10380 -75632 10436 -75588
rect 10480 -75632 10536 -75588
rect 10580 -75632 10636 -75588
rect 10680 -75632 10736 -75588
rect 10780 -75632 11236 -75588
rect 11280 -75632 11336 -75588
rect 11380 -75632 11436 -75588
rect 11480 -75632 11536 -75588
rect 11580 -75632 11636 -75588
rect 11680 -75632 11736 -75588
rect 11780 -75632 11836 -75588
rect 11880 -75632 11936 -75588
rect 11980 -75632 12036 -75588
rect 12080 -75632 12136 -75588
rect 12180 -75632 12236 -75588
rect 12280 -75632 12336 -75588
rect 12380 -75632 12436 -75588
rect 12480 -75632 12536 -75588
rect 12580 -75632 12636 -75588
rect 12680 -75632 12736 -75588
rect 12780 -75632 13236 -75588
rect 13280 -75632 13336 -75588
rect 13380 -75632 13436 -75588
rect 13480 -75632 13536 -75588
rect 13580 -75632 13636 -75588
rect 13680 -75632 13736 -75588
rect 13780 -75632 13836 -75588
rect 13880 -75632 13936 -75588
rect 13980 -75632 14036 -75588
rect 14080 -75632 14136 -75588
rect 14180 -75632 14236 -75588
rect 14280 -75632 14336 -75588
rect 14380 -75632 14436 -75588
rect 14480 -75632 14536 -75588
rect 14580 -75632 14636 -75588
rect 14680 -75632 14736 -75588
rect 14780 -75632 15236 -75588
rect 15280 -75632 15336 -75588
rect 15380 -75632 15436 -75588
rect 15480 -75632 15536 -75588
rect 15580 -75632 15636 -75588
rect 15680 -75632 15736 -75588
rect 15780 -75632 15836 -75588
rect 15880 -75632 15936 -75588
rect 15980 -75632 16036 -75588
rect 16080 -75632 16136 -75588
rect 16180 -75632 16236 -75588
rect 16280 -75632 16336 -75588
rect 16380 -75632 16436 -75588
rect 16480 -75632 16536 -75588
rect 16580 -75632 16636 -75588
rect 16680 -75632 16736 -75588
rect 16780 -75602 178308 -75588
rect 16780 -75632 177664 -75602
rect -108812 -75688 177664 -75632
rect -108812 -75732 9236 -75688
rect 9280 -75732 9336 -75688
rect 9380 -75732 9436 -75688
rect 9480 -75732 9536 -75688
rect 9580 -75732 9636 -75688
rect 9680 -75732 9736 -75688
rect 9780 -75732 9836 -75688
rect 9880 -75732 9936 -75688
rect 9980 -75732 10036 -75688
rect 10080 -75732 10136 -75688
rect 10180 -75732 10236 -75688
rect 10280 -75732 10336 -75688
rect 10380 -75732 10436 -75688
rect 10480 -75732 10536 -75688
rect 10580 -75732 10636 -75688
rect 10680 -75732 10736 -75688
rect 10780 -75732 11236 -75688
rect 11280 -75732 11336 -75688
rect 11380 -75732 11436 -75688
rect 11480 -75732 11536 -75688
rect 11580 -75732 11636 -75688
rect 11680 -75732 11736 -75688
rect 11780 -75732 11836 -75688
rect 11880 -75732 11936 -75688
rect 11980 -75732 12036 -75688
rect 12080 -75732 12136 -75688
rect 12180 -75732 12236 -75688
rect 12280 -75732 12336 -75688
rect 12380 -75732 12436 -75688
rect 12480 -75732 12536 -75688
rect 12580 -75732 12636 -75688
rect 12680 -75732 12736 -75688
rect 12780 -75732 13236 -75688
rect 13280 -75732 13336 -75688
rect 13380 -75732 13436 -75688
rect 13480 -75732 13536 -75688
rect 13580 -75732 13636 -75688
rect 13680 -75732 13736 -75688
rect 13780 -75732 13836 -75688
rect 13880 -75732 13936 -75688
rect 13980 -75732 14036 -75688
rect 14080 -75732 14136 -75688
rect 14180 -75732 14236 -75688
rect 14280 -75732 14336 -75688
rect 14380 -75732 14436 -75688
rect 14480 -75732 14536 -75688
rect 14580 -75732 14636 -75688
rect 14680 -75732 14736 -75688
rect 14780 -75732 15236 -75688
rect 15280 -75732 15336 -75688
rect 15380 -75732 15436 -75688
rect 15480 -75732 15536 -75688
rect 15580 -75732 15636 -75688
rect 15680 -75732 15736 -75688
rect 15780 -75732 15836 -75688
rect 15880 -75732 15936 -75688
rect 15980 -75732 16036 -75688
rect 16080 -75732 16136 -75688
rect 16180 -75732 16236 -75688
rect 16280 -75732 16336 -75688
rect 16380 -75732 16436 -75688
rect 16480 -75732 16536 -75688
rect 16580 -75732 16636 -75688
rect 16680 -75732 16736 -75688
rect 16780 -75732 177664 -75688
rect -108812 -75788 177664 -75732
rect -108812 -75832 9236 -75788
rect 9280 -75832 9336 -75788
rect 9380 -75832 9436 -75788
rect 9480 -75832 9536 -75788
rect 9580 -75832 9636 -75788
rect 9680 -75832 9736 -75788
rect 9780 -75832 9836 -75788
rect 9880 -75832 9936 -75788
rect 9980 -75832 10036 -75788
rect 10080 -75832 10136 -75788
rect 10180 -75832 10236 -75788
rect 10280 -75832 10336 -75788
rect 10380 -75832 10436 -75788
rect 10480 -75832 10536 -75788
rect 10580 -75832 10636 -75788
rect 10680 -75832 10736 -75788
rect 10780 -75832 11236 -75788
rect 11280 -75832 11336 -75788
rect 11380 -75832 11436 -75788
rect 11480 -75832 11536 -75788
rect 11580 -75832 11636 -75788
rect 11680 -75832 11736 -75788
rect 11780 -75832 11836 -75788
rect 11880 -75832 11936 -75788
rect 11980 -75832 12036 -75788
rect 12080 -75832 12136 -75788
rect 12180 -75832 12236 -75788
rect 12280 -75832 12336 -75788
rect 12380 -75832 12436 -75788
rect 12480 -75832 12536 -75788
rect 12580 -75832 12636 -75788
rect 12680 -75832 12736 -75788
rect 12780 -75832 13236 -75788
rect 13280 -75832 13336 -75788
rect 13380 -75832 13436 -75788
rect 13480 -75832 13536 -75788
rect 13580 -75832 13636 -75788
rect 13680 -75832 13736 -75788
rect 13780 -75832 13836 -75788
rect 13880 -75832 13936 -75788
rect 13980 -75832 14036 -75788
rect 14080 -75832 14136 -75788
rect 14180 -75832 14236 -75788
rect 14280 -75832 14336 -75788
rect 14380 -75832 14436 -75788
rect 14480 -75832 14536 -75788
rect 14580 -75832 14636 -75788
rect 14680 -75832 14736 -75788
rect 14780 -75832 15236 -75788
rect 15280 -75832 15336 -75788
rect 15380 -75832 15436 -75788
rect 15480 -75832 15536 -75788
rect 15580 -75832 15636 -75788
rect 15680 -75832 15736 -75788
rect 15780 -75832 15836 -75788
rect 15880 -75832 15936 -75788
rect 15980 -75832 16036 -75788
rect 16080 -75832 16136 -75788
rect 16180 -75832 16236 -75788
rect 16280 -75832 16336 -75788
rect 16380 -75832 16436 -75788
rect 16480 -75832 16536 -75788
rect 16580 -75832 16636 -75788
rect 16680 -75832 16736 -75788
rect 16780 -75832 177664 -75788
rect -108812 -75888 177664 -75832
rect -108812 -75932 9236 -75888
rect 9280 -75932 9336 -75888
rect 9380 -75932 9436 -75888
rect 9480 -75932 9536 -75888
rect 9580 -75932 9636 -75888
rect 9680 -75932 9736 -75888
rect 9780 -75932 9836 -75888
rect 9880 -75932 9936 -75888
rect 9980 -75932 10036 -75888
rect 10080 -75932 10136 -75888
rect 10180 -75932 10236 -75888
rect 10280 -75932 10336 -75888
rect 10380 -75932 10436 -75888
rect 10480 -75932 10536 -75888
rect 10580 -75932 10636 -75888
rect 10680 -75932 10736 -75888
rect 10780 -75932 11236 -75888
rect 11280 -75932 11336 -75888
rect 11380 -75932 11436 -75888
rect 11480 -75932 11536 -75888
rect 11580 -75932 11636 -75888
rect 11680 -75932 11736 -75888
rect 11780 -75932 11836 -75888
rect 11880 -75932 11936 -75888
rect 11980 -75932 12036 -75888
rect 12080 -75932 12136 -75888
rect 12180 -75932 12236 -75888
rect 12280 -75932 12336 -75888
rect 12380 -75932 12436 -75888
rect 12480 -75932 12536 -75888
rect 12580 -75932 12636 -75888
rect 12680 -75932 12736 -75888
rect 12780 -75932 13236 -75888
rect 13280 -75932 13336 -75888
rect 13380 -75932 13436 -75888
rect 13480 -75932 13536 -75888
rect 13580 -75932 13636 -75888
rect 13680 -75932 13736 -75888
rect 13780 -75932 13836 -75888
rect 13880 -75932 13936 -75888
rect 13980 -75932 14036 -75888
rect 14080 -75932 14136 -75888
rect 14180 -75932 14236 -75888
rect 14280 -75932 14336 -75888
rect 14380 -75932 14436 -75888
rect 14480 -75932 14536 -75888
rect 14580 -75932 14636 -75888
rect 14680 -75932 14736 -75888
rect 14780 -75932 15236 -75888
rect 15280 -75932 15336 -75888
rect 15380 -75932 15436 -75888
rect 15480 -75932 15536 -75888
rect 15580 -75932 15636 -75888
rect 15680 -75932 15736 -75888
rect 15780 -75932 15836 -75888
rect 15880 -75932 15936 -75888
rect 15980 -75932 16036 -75888
rect 16080 -75932 16136 -75888
rect 16180 -75932 16236 -75888
rect 16280 -75932 16336 -75888
rect 16380 -75932 16436 -75888
rect 16480 -75932 16536 -75888
rect 16580 -75932 16636 -75888
rect 16680 -75932 16736 -75888
rect 16780 -75932 177664 -75888
rect -108812 -75988 177664 -75932
rect -108812 -76032 9236 -75988
rect 9280 -76032 9336 -75988
rect 9380 -76032 9436 -75988
rect 9480 -76032 9536 -75988
rect 9580 -76032 9636 -75988
rect 9680 -76032 9736 -75988
rect 9780 -76032 9836 -75988
rect 9880 -76032 9936 -75988
rect 9980 -76032 10036 -75988
rect 10080 -76032 10136 -75988
rect 10180 -76032 10236 -75988
rect 10280 -76032 10336 -75988
rect 10380 -76032 10436 -75988
rect 10480 -76032 10536 -75988
rect 10580 -76032 10636 -75988
rect 10680 -76032 10736 -75988
rect 10780 -76032 11236 -75988
rect 11280 -76032 11336 -75988
rect 11380 -76032 11436 -75988
rect 11480 -76032 11536 -75988
rect 11580 -76032 11636 -75988
rect 11680 -76032 11736 -75988
rect 11780 -76032 11836 -75988
rect 11880 -76032 11936 -75988
rect 11980 -76032 12036 -75988
rect 12080 -76032 12136 -75988
rect 12180 -76032 12236 -75988
rect 12280 -76032 12336 -75988
rect 12380 -76032 12436 -75988
rect 12480 -76032 12536 -75988
rect 12580 -76032 12636 -75988
rect 12680 -76032 12736 -75988
rect 12780 -76032 13236 -75988
rect 13280 -76032 13336 -75988
rect 13380 -76032 13436 -75988
rect 13480 -76032 13536 -75988
rect 13580 -76032 13636 -75988
rect 13680 -76032 13736 -75988
rect 13780 -76032 13836 -75988
rect 13880 -76032 13936 -75988
rect 13980 -76032 14036 -75988
rect 14080 -76032 14136 -75988
rect 14180 -76032 14236 -75988
rect 14280 -76032 14336 -75988
rect 14380 -76032 14436 -75988
rect 14480 -76032 14536 -75988
rect 14580 -76032 14636 -75988
rect 14680 -76032 14736 -75988
rect 14780 -76032 15236 -75988
rect 15280 -76032 15336 -75988
rect 15380 -76032 15436 -75988
rect 15480 -76032 15536 -75988
rect 15580 -76032 15636 -75988
rect 15680 -76032 15736 -75988
rect 15780 -76032 15836 -75988
rect 15880 -76032 15936 -75988
rect 15980 -76032 16036 -75988
rect 16080 -76032 16136 -75988
rect 16180 -76032 16236 -75988
rect 16280 -76032 16336 -75988
rect 16380 -76032 16436 -75988
rect 16480 -76032 16536 -75988
rect 16580 -76032 16636 -75988
rect 16680 -76032 16736 -75988
rect 16780 -76032 177664 -75988
rect -108812 -76088 177664 -76032
rect -108812 -76132 9236 -76088
rect 9280 -76132 9336 -76088
rect 9380 -76132 9436 -76088
rect 9480 -76132 9536 -76088
rect 9580 -76132 9636 -76088
rect 9680 -76132 9736 -76088
rect 9780 -76132 9836 -76088
rect 9880 -76132 9936 -76088
rect 9980 -76132 10036 -76088
rect 10080 -76132 10136 -76088
rect 10180 -76132 10236 -76088
rect 10280 -76132 10336 -76088
rect 10380 -76132 10436 -76088
rect 10480 -76132 10536 -76088
rect 10580 -76132 10636 -76088
rect 10680 -76132 10736 -76088
rect 10780 -76132 11236 -76088
rect 11280 -76132 11336 -76088
rect 11380 -76132 11436 -76088
rect 11480 -76132 11536 -76088
rect 11580 -76132 11636 -76088
rect 11680 -76132 11736 -76088
rect 11780 -76132 11836 -76088
rect 11880 -76132 11936 -76088
rect 11980 -76132 12036 -76088
rect 12080 -76132 12136 -76088
rect 12180 -76132 12236 -76088
rect 12280 -76132 12336 -76088
rect 12380 -76132 12436 -76088
rect 12480 -76132 12536 -76088
rect 12580 -76132 12636 -76088
rect 12680 -76132 12736 -76088
rect 12780 -76132 13236 -76088
rect 13280 -76132 13336 -76088
rect 13380 -76132 13436 -76088
rect 13480 -76132 13536 -76088
rect 13580 -76132 13636 -76088
rect 13680 -76132 13736 -76088
rect 13780 -76132 13836 -76088
rect 13880 -76132 13936 -76088
rect 13980 -76132 14036 -76088
rect 14080 -76132 14136 -76088
rect 14180 -76132 14236 -76088
rect 14280 -76132 14336 -76088
rect 14380 -76132 14436 -76088
rect 14480 -76132 14536 -76088
rect 14580 -76132 14636 -76088
rect 14680 -76132 14736 -76088
rect 14780 -76132 15236 -76088
rect 15280 -76132 15336 -76088
rect 15380 -76132 15436 -76088
rect 15480 -76132 15536 -76088
rect 15580 -76132 15636 -76088
rect 15680 -76132 15736 -76088
rect 15780 -76132 15836 -76088
rect 15880 -76132 15936 -76088
rect 15980 -76132 16036 -76088
rect 16080 -76132 16136 -76088
rect 16180 -76132 16236 -76088
rect 16280 -76132 16336 -76088
rect 16380 -76132 16436 -76088
rect 16480 -76132 16536 -76088
rect 16580 -76132 16636 -76088
rect 16680 -76132 16736 -76088
rect 16780 -76132 177664 -76088
rect -108812 -76188 177664 -76132
rect -108812 -76232 9236 -76188
rect 9280 -76232 9336 -76188
rect 9380 -76232 9436 -76188
rect 9480 -76232 9536 -76188
rect 9580 -76232 9636 -76188
rect 9680 -76232 9736 -76188
rect 9780 -76232 9836 -76188
rect 9880 -76232 9936 -76188
rect 9980 -76232 10036 -76188
rect 10080 -76232 10136 -76188
rect 10180 -76232 10236 -76188
rect 10280 -76232 10336 -76188
rect 10380 -76232 10436 -76188
rect 10480 -76232 10536 -76188
rect 10580 -76232 10636 -76188
rect 10680 -76232 10736 -76188
rect 10780 -76232 11236 -76188
rect 11280 -76232 11336 -76188
rect 11380 -76232 11436 -76188
rect 11480 -76232 11536 -76188
rect 11580 -76232 11636 -76188
rect 11680 -76232 11736 -76188
rect 11780 -76232 11836 -76188
rect 11880 -76232 11936 -76188
rect 11980 -76232 12036 -76188
rect 12080 -76232 12136 -76188
rect 12180 -76232 12236 -76188
rect 12280 -76232 12336 -76188
rect 12380 -76232 12436 -76188
rect 12480 -76232 12536 -76188
rect 12580 -76232 12636 -76188
rect 12680 -76232 12736 -76188
rect 12780 -76232 13236 -76188
rect 13280 -76232 13336 -76188
rect 13380 -76232 13436 -76188
rect 13480 -76232 13536 -76188
rect 13580 -76232 13636 -76188
rect 13680 -76232 13736 -76188
rect 13780 -76232 13836 -76188
rect 13880 -76232 13936 -76188
rect 13980 -76232 14036 -76188
rect 14080 -76232 14136 -76188
rect 14180 -76232 14236 -76188
rect 14280 -76232 14336 -76188
rect 14380 -76232 14436 -76188
rect 14480 -76232 14536 -76188
rect 14580 -76232 14636 -76188
rect 14680 -76232 14736 -76188
rect 14780 -76232 15236 -76188
rect 15280 -76232 15336 -76188
rect 15380 -76232 15436 -76188
rect 15480 -76232 15536 -76188
rect 15580 -76232 15636 -76188
rect 15680 -76232 15736 -76188
rect 15780 -76232 15836 -76188
rect 15880 -76232 15936 -76188
rect 15980 -76232 16036 -76188
rect 16080 -76232 16136 -76188
rect 16180 -76232 16236 -76188
rect 16280 -76232 16336 -76188
rect 16380 -76232 16436 -76188
rect 16480 -76232 16536 -76188
rect 16580 -76232 16636 -76188
rect 16680 -76232 16736 -76188
rect 16780 -76232 177664 -76188
rect -108812 -76288 177664 -76232
rect -108812 -76332 9236 -76288
rect 9280 -76332 9336 -76288
rect 9380 -76332 9436 -76288
rect 9480 -76332 9536 -76288
rect 9580 -76332 9636 -76288
rect 9680 -76332 9736 -76288
rect 9780 -76332 9836 -76288
rect 9880 -76332 9936 -76288
rect 9980 -76332 10036 -76288
rect 10080 -76332 10136 -76288
rect 10180 -76332 10236 -76288
rect 10280 -76332 10336 -76288
rect 10380 -76332 10436 -76288
rect 10480 -76332 10536 -76288
rect 10580 -76332 10636 -76288
rect 10680 -76332 10736 -76288
rect 10780 -76332 11236 -76288
rect 11280 -76332 11336 -76288
rect 11380 -76332 11436 -76288
rect 11480 -76332 11536 -76288
rect 11580 -76332 11636 -76288
rect 11680 -76332 11736 -76288
rect 11780 -76332 11836 -76288
rect 11880 -76332 11936 -76288
rect 11980 -76332 12036 -76288
rect 12080 -76332 12136 -76288
rect 12180 -76332 12236 -76288
rect 12280 -76332 12336 -76288
rect 12380 -76332 12436 -76288
rect 12480 -76332 12536 -76288
rect 12580 -76332 12636 -76288
rect 12680 -76332 12736 -76288
rect 12780 -76332 13236 -76288
rect 13280 -76332 13336 -76288
rect 13380 -76332 13436 -76288
rect 13480 -76332 13536 -76288
rect 13580 -76332 13636 -76288
rect 13680 -76332 13736 -76288
rect 13780 -76332 13836 -76288
rect 13880 -76332 13936 -76288
rect 13980 -76332 14036 -76288
rect 14080 -76332 14136 -76288
rect 14180 -76332 14236 -76288
rect 14280 -76332 14336 -76288
rect 14380 -76332 14436 -76288
rect 14480 -76332 14536 -76288
rect 14580 -76332 14636 -76288
rect 14680 -76332 14736 -76288
rect 14780 -76332 15236 -76288
rect 15280 -76332 15336 -76288
rect 15380 -76332 15436 -76288
rect 15480 -76332 15536 -76288
rect 15580 -76332 15636 -76288
rect 15680 -76332 15736 -76288
rect 15780 -76332 15836 -76288
rect 15880 -76332 15936 -76288
rect 15980 -76332 16036 -76288
rect 16080 -76332 16136 -76288
rect 16180 -76332 16236 -76288
rect 16280 -76332 16336 -76288
rect 16380 -76332 16436 -76288
rect 16480 -76332 16536 -76288
rect 16580 -76332 16636 -76288
rect 16680 -76332 16736 -76288
rect 16780 -76332 177664 -76288
rect -108812 -76388 177664 -76332
rect -108812 -76432 9236 -76388
rect 9280 -76432 9336 -76388
rect 9380 -76432 9436 -76388
rect 9480 -76432 9536 -76388
rect 9580 -76432 9636 -76388
rect 9680 -76432 9736 -76388
rect 9780 -76432 9836 -76388
rect 9880 -76432 9936 -76388
rect 9980 -76432 10036 -76388
rect 10080 -76432 10136 -76388
rect 10180 -76432 10236 -76388
rect 10280 -76432 10336 -76388
rect 10380 -76432 10436 -76388
rect 10480 -76432 10536 -76388
rect 10580 -76432 10636 -76388
rect 10680 -76432 10736 -76388
rect 10780 -76432 11236 -76388
rect 11280 -76432 11336 -76388
rect 11380 -76432 11436 -76388
rect 11480 -76432 11536 -76388
rect 11580 -76432 11636 -76388
rect 11680 -76432 11736 -76388
rect 11780 -76432 11836 -76388
rect 11880 -76432 11936 -76388
rect 11980 -76432 12036 -76388
rect 12080 -76432 12136 -76388
rect 12180 -76432 12236 -76388
rect 12280 -76432 12336 -76388
rect 12380 -76432 12436 -76388
rect 12480 -76432 12536 -76388
rect 12580 -76432 12636 -76388
rect 12680 -76432 12736 -76388
rect 12780 -76432 13236 -76388
rect 13280 -76432 13336 -76388
rect 13380 -76432 13436 -76388
rect 13480 -76432 13536 -76388
rect 13580 -76432 13636 -76388
rect 13680 -76432 13736 -76388
rect 13780 -76432 13836 -76388
rect 13880 -76432 13936 -76388
rect 13980 -76432 14036 -76388
rect 14080 -76432 14136 -76388
rect 14180 -76432 14236 -76388
rect 14280 -76432 14336 -76388
rect 14380 -76432 14436 -76388
rect 14480 -76432 14536 -76388
rect 14580 -76432 14636 -76388
rect 14680 -76432 14736 -76388
rect 14780 -76432 15236 -76388
rect 15280 -76432 15336 -76388
rect 15380 -76432 15436 -76388
rect 15480 -76432 15536 -76388
rect 15580 -76432 15636 -76388
rect 15680 -76432 15736 -76388
rect 15780 -76432 15836 -76388
rect 15880 -76432 15936 -76388
rect 15980 -76432 16036 -76388
rect 16080 -76432 16136 -76388
rect 16180 -76432 16236 -76388
rect 16280 -76432 16336 -76388
rect 16380 -76432 16436 -76388
rect 16480 -76432 16536 -76388
rect 16580 -76432 16636 -76388
rect 16680 -76432 16736 -76388
rect 16780 -76432 177664 -76388
rect -108812 -76488 177664 -76432
rect -108812 -76532 9236 -76488
rect 9280 -76532 9336 -76488
rect 9380 -76532 9436 -76488
rect 9480 -76532 9536 -76488
rect 9580 -76532 9636 -76488
rect 9680 -76532 9736 -76488
rect 9780 -76532 9836 -76488
rect 9880 -76532 9936 -76488
rect 9980 -76532 10036 -76488
rect 10080 -76532 10136 -76488
rect 10180 -76532 10236 -76488
rect 10280 -76532 10336 -76488
rect 10380 -76532 10436 -76488
rect 10480 -76532 10536 -76488
rect 10580 -76532 10636 -76488
rect 10680 -76532 10736 -76488
rect 10780 -76532 11236 -76488
rect 11280 -76532 11336 -76488
rect 11380 -76532 11436 -76488
rect 11480 -76532 11536 -76488
rect 11580 -76532 11636 -76488
rect 11680 -76532 11736 -76488
rect 11780 -76532 11836 -76488
rect 11880 -76532 11936 -76488
rect 11980 -76532 12036 -76488
rect 12080 -76532 12136 -76488
rect 12180 -76532 12236 -76488
rect 12280 -76532 12336 -76488
rect 12380 -76532 12436 -76488
rect 12480 -76532 12536 -76488
rect 12580 -76532 12636 -76488
rect 12680 -76532 12736 -76488
rect 12780 -76532 13236 -76488
rect 13280 -76532 13336 -76488
rect 13380 -76532 13436 -76488
rect 13480 -76532 13536 -76488
rect 13580 -76532 13636 -76488
rect 13680 -76532 13736 -76488
rect 13780 -76532 13836 -76488
rect 13880 -76532 13936 -76488
rect 13980 -76532 14036 -76488
rect 14080 -76532 14136 -76488
rect 14180 -76532 14236 -76488
rect 14280 -76532 14336 -76488
rect 14380 -76532 14436 -76488
rect 14480 -76532 14536 -76488
rect 14580 -76532 14636 -76488
rect 14680 -76532 14736 -76488
rect 14780 -76532 15236 -76488
rect 15280 -76532 15336 -76488
rect 15380 -76532 15436 -76488
rect 15480 -76532 15536 -76488
rect 15580 -76532 15636 -76488
rect 15680 -76532 15736 -76488
rect 15780 -76532 15836 -76488
rect 15880 -76532 15936 -76488
rect 15980 -76532 16036 -76488
rect 16080 -76532 16136 -76488
rect 16180 -76532 16236 -76488
rect 16280 -76532 16336 -76488
rect 16380 -76532 16436 -76488
rect 16480 -76532 16536 -76488
rect 16580 -76532 16636 -76488
rect 16680 -76532 16736 -76488
rect 16780 -76532 177664 -76488
rect -108812 -76588 177664 -76532
rect -108812 -76632 9236 -76588
rect 9280 -76632 9336 -76588
rect 9380 -76632 9436 -76588
rect 9480 -76632 9536 -76588
rect 9580 -76632 9636 -76588
rect 9680 -76632 9736 -76588
rect 9780 -76632 9836 -76588
rect 9880 -76632 9936 -76588
rect 9980 -76632 10036 -76588
rect 10080 -76632 10136 -76588
rect 10180 -76632 10236 -76588
rect 10280 -76632 10336 -76588
rect 10380 -76632 10436 -76588
rect 10480 -76632 10536 -76588
rect 10580 -76632 10636 -76588
rect 10680 -76632 10736 -76588
rect 10780 -76632 11236 -76588
rect 11280 -76632 11336 -76588
rect 11380 -76632 11436 -76588
rect 11480 -76632 11536 -76588
rect 11580 -76632 11636 -76588
rect 11680 -76632 11736 -76588
rect 11780 -76632 11836 -76588
rect 11880 -76632 11936 -76588
rect 11980 -76632 12036 -76588
rect 12080 -76632 12136 -76588
rect 12180 -76632 12236 -76588
rect 12280 -76632 12336 -76588
rect 12380 -76632 12436 -76588
rect 12480 -76632 12536 -76588
rect 12580 -76632 12636 -76588
rect 12680 -76632 12736 -76588
rect 12780 -76632 13236 -76588
rect 13280 -76632 13336 -76588
rect 13380 -76632 13436 -76588
rect 13480 -76632 13536 -76588
rect 13580 -76632 13636 -76588
rect 13680 -76632 13736 -76588
rect 13780 -76632 13836 -76588
rect 13880 -76632 13936 -76588
rect 13980 -76632 14036 -76588
rect 14080 -76632 14136 -76588
rect 14180 -76632 14236 -76588
rect 14280 -76632 14336 -76588
rect 14380 -76632 14436 -76588
rect 14480 -76632 14536 -76588
rect 14580 -76632 14636 -76588
rect 14680 -76632 14736 -76588
rect 14780 -76632 15236 -76588
rect 15280 -76632 15336 -76588
rect 15380 -76632 15436 -76588
rect 15480 -76632 15536 -76588
rect 15580 -76632 15636 -76588
rect 15680 -76632 15736 -76588
rect 15780 -76632 15836 -76588
rect 15880 -76632 15936 -76588
rect 15980 -76632 16036 -76588
rect 16080 -76632 16136 -76588
rect 16180 -76632 16236 -76588
rect 16280 -76632 16336 -76588
rect 16380 -76632 16436 -76588
rect 16480 -76632 16536 -76588
rect 16580 -76632 16636 -76588
rect 16680 -76632 16736 -76588
rect 16780 -76632 177664 -76588
rect -108812 -76688 177664 -76632
rect -108812 -76732 9236 -76688
rect 9280 -76732 9336 -76688
rect 9380 -76732 9436 -76688
rect 9480 -76732 9536 -76688
rect 9580 -76732 9636 -76688
rect 9680 -76732 9736 -76688
rect 9780 -76732 9836 -76688
rect 9880 -76732 9936 -76688
rect 9980 -76732 10036 -76688
rect 10080 -76732 10136 -76688
rect 10180 -76732 10236 -76688
rect 10280 -76732 10336 -76688
rect 10380 -76732 10436 -76688
rect 10480 -76732 10536 -76688
rect 10580 -76732 10636 -76688
rect 10680 -76732 10736 -76688
rect 10780 -76732 11236 -76688
rect 11280 -76732 11336 -76688
rect 11380 -76732 11436 -76688
rect 11480 -76732 11536 -76688
rect 11580 -76732 11636 -76688
rect 11680 -76732 11736 -76688
rect 11780 -76732 11836 -76688
rect 11880 -76732 11936 -76688
rect 11980 -76732 12036 -76688
rect 12080 -76732 12136 -76688
rect 12180 -76732 12236 -76688
rect 12280 -76732 12336 -76688
rect 12380 -76732 12436 -76688
rect 12480 -76732 12536 -76688
rect 12580 -76732 12636 -76688
rect 12680 -76732 12736 -76688
rect 12780 -76732 13236 -76688
rect 13280 -76732 13336 -76688
rect 13380 -76732 13436 -76688
rect 13480 -76732 13536 -76688
rect 13580 -76732 13636 -76688
rect 13680 -76732 13736 -76688
rect 13780 -76732 13836 -76688
rect 13880 -76732 13936 -76688
rect 13980 -76732 14036 -76688
rect 14080 -76732 14136 -76688
rect 14180 -76732 14236 -76688
rect 14280 -76732 14336 -76688
rect 14380 -76732 14436 -76688
rect 14480 -76732 14536 -76688
rect 14580 -76732 14636 -76688
rect 14680 -76732 14736 -76688
rect 14780 -76732 15236 -76688
rect 15280 -76732 15336 -76688
rect 15380 -76732 15436 -76688
rect 15480 -76732 15536 -76688
rect 15580 -76732 15636 -76688
rect 15680 -76732 15736 -76688
rect 15780 -76732 15836 -76688
rect 15880 -76732 15936 -76688
rect 15980 -76732 16036 -76688
rect 16080 -76732 16136 -76688
rect 16180 -76732 16236 -76688
rect 16280 -76732 16336 -76688
rect 16380 -76732 16436 -76688
rect 16480 -76732 16536 -76688
rect 16580 -76732 16636 -76688
rect 16680 -76732 16736 -76688
rect 16780 -76732 177664 -76688
rect -108812 -76921 177664 -76732
rect -109116 -80455 177360 -80270
rect -109116 -80459 80737 -80455
rect -109116 -80503 -82968 -80459
rect -82924 -80503 -82868 -80459
rect -82824 -80503 -82768 -80459
rect -82724 -80503 -82668 -80459
rect -82624 -80503 -82568 -80459
rect -82524 -80503 -82468 -80459
rect -82424 -80503 -82368 -80459
rect -82324 -80503 -82268 -80459
rect -82224 -80503 -82168 -80459
rect -82124 -80503 -82068 -80459
rect -82024 -80503 -81968 -80459
rect -81924 -80503 -81868 -80459
rect -81824 -80503 -81768 -80459
rect -81724 -80503 -81668 -80459
rect -81624 -80503 -81568 -80459
rect -81524 -80503 -81468 -80459
rect -81424 -80503 -80968 -80459
rect -80924 -80503 -80868 -80459
rect -80824 -80503 -80768 -80459
rect -80724 -80503 -80668 -80459
rect -80624 -80503 -80568 -80459
rect -80524 -80503 -80468 -80459
rect -80424 -80503 -80368 -80459
rect -80324 -80503 -80268 -80459
rect -80224 -80503 -80168 -80459
rect -80124 -80503 -80068 -80459
rect -80024 -80503 -79968 -80459
rect -79924 -80503 -79868 -80459
rect -79824 -80503 -79768 -80459
rect -79724 -80503 -79668 -80459
rect -79624 -80503 -79568 -80459
rect -79524 -80503 -79468 -80459
rect -79424 -80503 -78968 -80459
rect -78924 -80503 -78868 -80459
rect -78824 -80503 -78768 -80459
rect -78724 -80503 -78668 -80459
rect -78624 -80503 -78568 -80459
rect -78524 -80503 -78468 -80459
rect -78424 -80503 -78368 -80459
rect -78324 -80503 -78268 -80459
rect -78224 -80503 -78168 -80459
rect -78124 -80503 -78068 -80459
rect -78024 -80503 -77968 -80459
rect -77924 -80503 -77868 -80459
rect -77824 -80503 -77768 -80459
rect -77724 -80503 -77668 -80459
rect -77624 -80503 -77568 -80459
rect -77524 -80503 -77468 -80459
rect -77424 -80503 -76968 -80459
rect -76924 -80503 -76868 -80459
rect -76824 -80503 -76768 -80459
rect -76724 -80503 -76668 -80459
rect -76624 -80503 -76568 -80459
rect -76524 -80503 -76468 -80459
rect -76424 -80503 -76368 -80459
rect -76324 -80503 -76268 -80459
rect -76224 -80503 -76168 -80459
rect -76124 -80503 -76068 -80459
rect -76024 -80503 -75968 -80459
rect -75924 -80503 -75868 -80459
rect -75824 -80503 -75768 -80459
rect -75724 -80503 -75668 -80459
rect -75624 -80503 -75568 -80459
rect -75524 -80503 -75468 -80459
rect -75424 -80461 80737 -80459
rect -75424 -80503 -50017 -80461
rect -109116 -80505 -50017 -80503
rect -49973 -80505 -49917 -80461
rect -49873 -80505 -49817 -80461
rect -49773 -80505 -49717 -80461
rect -49673 -80505 -49617 -80461
rect -49573 -80505 -49517 -80461
rect -49473 -80505 -49417 -80461
rect -49373 -80505 -49317 -80461
rect -49273 -80505 -49217 -80461
rect -49173 -80505 -49117 -80461
rect -49073 -80505 -49017 -80461
rect -48973 -80505 -48917 -80461
rect -48873 -80505 -48817 -80461
rect -48773 -80505 -48717 -80461
rect -48673 -80505 -48617 -80461
rect -48573 -80505 -48517 -80461
rect -48473 -80505 -48017 -80461
rect -47973 -80505 -47917 -80461
rect -47873 -80505 -47817 -80461
rect -47773 -80505 -47717 -80461
rect -47673 -80505 -47617 -80461
rect -47573 -80505 -47517 -80461
rect -47473 -80505 -47417 -80461
rect -47373 -80505 -47317 -80461
rect -47273 -80505 -47217 -80461
rect -47173 -80505 -47117 -80461
rect -47073 -80505 -47017 -80461
rect -46973 -80505 -46917 -80461
rect -46873 -80505 -46817 -80461
rect -46773 -80505 -46717 -80461
rect -46673 -80505 -46617 -80461
rect -46573 -80505 -46517 -80461
rect -46473 -80505 -46017 -80461
rect -45973 -80505 -45917 -80461
rect -45873 -80505 -45817 -80461
rect -45773 -80505 -45717 -80461
rect -45673 -80505 -45617 -80461
rect -45573 -80505 -45517 -80461
rect -45473 -80505 -45417 -80461
rect -45373 -80505 -45317 -80461
rect -45273 -80505 -45217 -80461
rect -45173 -80505 -45117 -80461
rect -45073 -80505 -45017 -80461
rect -44973 -80505 -44917 -80461
rect -44873 -80505 -44817 -80461
rect -44773 -80505 -44717 -80461
rect -44673 -80505 -44617 -80461
rect -44573 -80505 -44517 -80461
rect -44473 -80505 -44017 -80461
rect -43973 -80505 -43917 -80461
rect -43873 -80505 -43817 -80461
rect -43773 -80505 -43717 -80461
rect -43673 -80505 -43617 -80461
rect -43573 -80505 -43517 -80461
rect -43473 -80505 -43417 -80461
rect -43373 -80505 -43317 -80461
rect -43273 -80505 -43217 -80461
rect -43173 -80505 -43117 -80461
rect -43073 -80505 -43017 -80461
rect -42973 -80505 -42917 -80461
rect -42873 -80505 -42817 -80461
rect -42773 -80505 -42717 -80461
rect -42673 -80505 -42617 -80461
rect -42573 -80505 -42517 -80461
rect -42473 -80499 80737 -80461
rect 80781 -80499 80837 -80455
rect 80881 -80499 80937 -80455
rect 80981 -80499 81037 -80455
rect 81081 -80499 81137 -80455
rect 81181 -80499 81237 -80455
rect 81281 -80499 81337 -80455
rect 81381 -80499 81437 -80455
rect 81481 -80499 81537 -80455
rect 81581 -80499 81637 -80455
rect 81681 -80499 81737 -80455
rect 81781 -80499 81837 -80455
rect 81881 -80499 81937 -80455
rect 81981 -80499 82037 -80455
rect 82081 -80499 82137 -80455
rect 82181 -80499 82237 -80455
rect 82281 -80499 82737 -80455
rect 82781 -80499 82837 -80455
rect 82881 -80499 82937 -80455
rect 82981 -80499 83037 -80455
rect 83081 -80499 83137 -80455
rect 83181 -80499 83237 -80455
rect 83281 -80499 83337 -80455
rect 83381 -80499 83437 -80455
rect 83481 -80499 83537 -80455
rect 83581 -80499 83637 -80455
rect 83681 -80499 83737 -80455
rect 83781 -80499 83837 -80455
rect 83881 -80499 83937 -80455
rect 83981 -80499 84037 -80455
rect 84081 -80499 84137 -80455
rect 84181 -80499 84237 -80455
rect 84281 -80499 84737 -80455
rect 84781 -80499 84837 -80455
rect 84881 -80499 84937 -80455
rect 84981 -80499 85037 -80455
rect 85081 -80499 85137 -80455
rect 85181 -80499 85237 -80455
rect 85281 -80499 85337 -80455
rect 85381 -80499 85437 -80455
rect 85481 -80499 85537 -80455
rect 85581 -80499 85637 -80455
rect 85681 -80499 85737 -80455
rect 85781 -80499 85837 -80455
rect 85881 -80499 85937 -80455
rect 85981 -80499 86037 -80455
rect 86081 -80499 86137 -80455
rect 86181 -80499 86237 -80455
rect 86281 -80499 86737 -80455
rect 86781 -80499 86837 -80455
rect 86881 -80499 86937 -80455
rect 86981 -80499 87037 -80455
rect 87081 -80499 87137 -80455
rect 87181 -80499 87237 -80455
rect 87281 -80499 87337 -80455
rect 87381 -80499 87437 -80455
rect 87481 -80499 87537 -80455
rect 87581 -80499 87637 -80455
rect 87681 -80499 87737 -80455
rect 87781 -80499 87837 -80455
rect 87881 -80499 87937 -80455
rect 87981 -80499 88037 -80455
rect 88081 -80499 88137 -80455
rect 88181 -80499 88237 -80455
rect 88281 -80499 177360 -80455
rect -42473 -80505 177360 -80499
rect -109116 -80555 177360 -80505
rect -109116 -80559 80737 -80555
rect -109116 -80603 -82968 -80559
rect -82924 -80603 -82868 -80559
rect -82824 -80603 -82768 -80559
rect -82724 -80603 -82668 -80559
rect -82624 -80603 -82568 -80559
rect -82524 -80603 -82468 -80559
rect -82424 -80603 -82368 -80559
rect -82324 -80603 -82268 -80559
rect -82224 -80603 -82168 -80559
rect -82124 -80603 -82068 -80559
rect -82024 -80603 -81968 -80559
rect -81924 -80603 -81868 -80559
rect -81824 -80603 -81768 -80559
rect -81724 -80603 -81668 -80559
rect -81624 -80603 -81568 -80559
rect -81524 -80603 -81468 -80559
rect -81424 -80603 -80968 -80559
rect -80924 -80603 -80868 -80559
rect -80824 -80603 -80768 -80559
rect -80724 -80603 -80668 -80559
rect -80624 -80603 -80568 -80559
rect -80524 -80603 -80468 -80559
rect -80424 -80603 -80368 -80559
rect -80324 -80603 -80268 -80559
rect -80224 -80603 -80168 -80559
rect -80124 -80603 -80068 -80559
rect -80024 -80603 -79968 -80559
rect -79924 -80603 -79868 -80559
rect -79824 -80603 -79768 -80559
rect -79724 -80603 -79668 -80559
rect -79624 -80603 -79568 -80559
rect -79524 -80603 -79468 -80559
rect -79424 -80603 -78968 -80559
rect -78924 -80603 -78868 -80559
rect -78824 -80603 -78768 -80559
rect -78724 -80603 -78668 -80559
rect -78624 -80603 -78568 -80559
rect -78524 -80603 -78468 -80559
rect -78424 -80603 -78368 -80559
rect -78324 -80603 -78268 -80559
rect -78224 -80603 -78168 -80559
rect -78124 -80603 -78068 -80559
rect -78024 -80603 -77968 -80559
rect -77924 -80603 -77868 -80559
rect -77824 -80603 -77768 -80559
rect -77724 -80603 -77668 -80559
rect -77624 -80603 -77568 -80559
rect -77524 -80603 -77468 -80559
rect -77424 -80603 -76968 -80559
rect -76924 -80603 -76868 -80559
rect -76824 -80603 -76768 -80559
rect -76724 -80603 -76668 -80559
rect -76624 -80603 -76568 -80559
rect -76524 -80603 -76468 -80559
rect -76424 -80603 -76368 -80559
rect -76324 -80603 -76268 -80559
rect -76224 -80603 -76168 -80559
rect -76124 -80603 -76068 -80559
rect -76024 -80603 -75968 -80559
rect -75924 -80603 -75868 -80559
rect -75824 -80603 -75768 -80559
rect -75724 -80603 -75668 -80559
rect -75624 -80603 -75568 -80559
rect -75524 -80603 -75468 -80559
rect -75424 -80561 80737 -80559
rect -75424 -80603 -50017 -80561
rect -109116 -80605 -50017 -80603
rect -49973 -80605 -49917 -80561
rect -49873 -80605 -49817 -80561
rect -49773 -80605 -49717 -80561
rect -49673 -80605 -49617 -80561
rect -49573 -80605 -49517 -80561
rect -49473 -80605 -49417 -80561
rect -49373 -80605 -49317 -80561
rect -49273 -80605 -49217 -80561
rect -49173 -80605 -49117 -80561
rect -49073 -80605 -49017 -80561
rect -48973 -80605 -48917 -80561
rect -48873 -80605 -48817 -80561
rect -48773 -80605 -48717 -80561
rect -48673 -80605 -48617 -80561
rect -48573 -80605 -48517 -80561
rect -48473 -80605 -48017 -80561
rect -47973 -80605 -47917 -80561
rect -47873 -80605 -47817 -80561
rect -47773 -80605 -47717 -80561
rect -47673 -80605 -47617 -80561
rect -47573 -80605 -47517 -80561
rect -47473 -80605 -47417 -80561
rect -47373 -80605 -47317 -80561
rect -47273 -80605 -47217 -80561
rect -47173 -80605 -47117 -80561
rect -47073 -80605 -47017 -80561
rect -46973 -80605 -46917 -80561
rect -46873 -80605 -46817 -80561
rect -46773 -80605 -46717 -80561
rect -46673 -80605 -46617 -80561
rect -46573 -80605 -46517 -80561
rect -46473 -80605 -46017 -80561
rect -45973 -80605 -45917 -80561
rect -45873 -80605 -45817 -80561
rect -45773 -80605 -45717 -80561
rect -45673 -80605 -45617 -80561
rect -45573 -80605 -45517 -80561
rect -45473 -80605 -45417 -80561
rect -45373 -80605 -45317 -80561
rect -45273 -80605 -45217 -80561
rect -45173 -80605 -45117 -80561
rect -45073 -80605 -45017 -80561
rect -44973 -80605 -44917 -80561
rect -44873 -80605 -44817 -80561
rect -44773 -80605 -44717 -80561
rect -44673 -80605 -44617 -80561
rect -44573 -80605 -44517 -80561
rect -44473 -80605 -44017 -80561
rect -43973 -80605 -43917 -80561
rect -43873 -80605 -43817 -80561
rect -43773 -80605 -43717 -80561
rect -43673 -80605 -43617 -80561
rect -43573 -80605 -43517 -80561
rect -43473 -80605 -43417 -80561
rect -43373 -80605 -43317 -80561
rect -43273 -80605 -43217 -80561
rect -43173 -80605 -43117 -80561
rect -43073 -80605 -43017 -80561
rect -42973 -80605 -42917 -80561
rect -42873 -80605 -42817 -80561
rect -42773 -80605 -42717 -80561
rect -42673 -80605 -42617 -80561
rect -42573 -80605 -42517 -80561
rect -42473 -80599 80737 -80561
rect 80781 -80599 80837 -80555
rect 80881 -80599 80937 -80555
rect 80981 -80599 81037 -80555
rect 81081 -80599 81137 -80555
rect 81181 -80599 81237 -80555
rect 81281 -80599 81337 -80555
rect 81381 -80599 81437 -80555
rect 81481 -80599 81537 -80555
rect 81581 -80599 81637 -80555
rect 81681 -80599 81737 -80555
rect 81781 -80599 81837 -80555
rect 81881 -80599 81937 -80555
rect 81981 -80599 82037 -80555
rect 82081 -80599 82137 -80555
rect 82181 -80599 82237 -80555
rect 82281 -80599 82737 -80555
rect 82781 -80599 82837 -80555
rect 82881 -80599 82937 -80555
rect 82981 -80599 83037 -80555
rect 83081 -80599 83137 -80555
rect 83181 -80599 83237 -80555
rect 83281 -80599 83337 -80555
rect 83381 -80599 83437 -80555
rect 83481 -80599 83537 -80555
rect 83581 -80599 83637 -80555
rect 83681 -80599 83737 -80555
rect 83781 -80599 83837 -80555
rect 83881 -80599 83937 -80555
rect 83981 -80599 84037 -80555
rect 84081 -80599 84137 -80555
rect 84181 -80599 84237 -80555
rect 84281 -80599 84737 -80555
rect 84781 -80599 84837 -80555
rect 84881 -80599 84937 -80555
rect 84981 -80599 85037 -80555
rect 85081 -80599 85137 -80555
rect 85181 -80599 85237 -80555
rect 85281 -80599 85337 -80555
rect 85381 -80599 85437 -80555
rect 85481 -80599 85537 -80555
rect 85581 -80599 85637 -80555
rect 85681 -80599 85737 -80555
rect 85781 -80599 85837 -80555
rect 85881 -80599 85937 -80555
rect 85981 -80599 86037 -80555
rect 86081 -80599 86137 -80555
rect 86181 -80599 86237 -80555
rect 86281 -80599 86737 -80555
rect 86781 -80599 86837 -80555
rect 86881 -80599 86937 -80555
rect 86981 -80599 87037 -80555
rect 87081 -80599 87137 -80555
rect 87181 -80599 87237 -80555
rect 87281 -80599 87337 -80555
rect 87381 -80599 87437 -80555
rect 87481 -80599 87537 -80555
rect 87581 -80599 87637 -80555
rect 87681 -80599 87737 -80555
rect 87781 -80599 87837 -80555
rect 87881 -80599 87937 -80555
rect 87981 -80599 88037 -80555
rect 88081 -80599 88137 -80555
rect 88181 -80599 88237 -80555
rect 88281 -80599 177360 -80555
rect -42473 -80605 177360 -80599
rect -109116 -80655 177360 -80605
rect -109116 -80659 80737 -80655
rect -109116 -80703 -82968 -80659
rect -82924 -80703 -82868 -80659
rect -82824 -80703 -82768 -80659
rect -82724 -80703 -82668 -80659
rect -82624 -80703 -82568 -80659
rect -82524 -80703 -82468 -80659
rect -82424 -80703 -82368 -80659
rect -82324 -80703 -82268 -80659
rect -82224 -80703 -82168 -80659
rect -82124 -80703 -82068 -80659
rect -82024 -80703 -81968 -80659
rect -81924 -80703 -81868 -80659
rect -81824 -80703 -81768 -80659
rect -81724 -80703 -81668 -80659
rect -81624 -80703 -81568 -80659
rect -81524 -80703 -81468 -80659
rect -81424 -80703 -80968 -80659
rect -80924 -80703 -80868 -80659
rect -80824 -80703 -80768 -80659
rect -80724 -80703 -80668 -80659
rect -80624 -80703 -80568 -80659
rect -80524 -80703 -80468 -80659
rect -80424 -80703 -80368 -80659
rect -80324 -80703 -80268 -80659
rect -80224 -80703 -80168 -80659
rect -80124 -80703 -80068 -80659
rect -80024 -80703 -79968 -80659
rect -79924 -80703 -79868 -80659
rect -79824 -80703 -79768 -80659
rect -79724 -80703 -79668 -80659
rect -79624 -80703 -79568 -80659
rect -79524 -80703 -79468 -80659
rect -79424 -80703 -78968 -80659
rect -78924 -80703 -78868 -80659
rect -78824 -80703 -78768 -80659
rect -78724 -80703 -78668 -80659
rect -78624 -80703 -78568 -80659
rect -78524 -80703 -78468 -80659
rect -78424 -80703 -78368 -80659
rect -78324 -80703 -78268 -80659
rect -78224 -80703 -78168 -80659
rect -78124 -80703 -78068 -80659
rect -78024 -80703 -77968 -80659
rect -77924 -80703 -77868 -80659
rect -77824 -80703 -77768 -80659
rect -77724 -80703 -77668 -80659
rect -77624 -80703 -77568 -80659
rect -77524 -80703 -77468 -80659
rect -77424 -80703 -76968 -80659
rect -76924 -80703 -76868 -80659
rect -76824 -80703 -76768 -80659
rect -76724 -80703 -76668 -80659
rect -76624 -80703 -76568 -80659
rect -76524 -80703 -76468 -80659
rect -76424 -80703 -76368 -80659
rect -76324 -80703 -76268 -80659
rect -76224 -80703 -76168 -80659
rect -76124 -80703 -76068 -80659
rect -76024 -80703 -75968 -80659
rect -75924 -80703 -75868 -80659
rect -75824 -80703 -75768 -80659
rect -75724 -80703 -75668 -80659
rect -75624 -80703 -75568 -80659
rect -75524 -80703 -75468 -80659
rect -75424 -80661 80737 -80659
rect -75424 -80703 -50017 -80661
rect -109116 -80705 -50017 -80703
rect -49973 -80705 -49917 -80661
rect -49873 -80705 -49817 -80661
rect -49773 -80705 -49717 -80661
rect -49673 -80705 -49617 -80661
rect -49573 -80705 -49517 -80661
rect -49473 -80705 -49417 -80661
rect -49373 -80705 -49317 -80661
rect -49273 -80705 -49217 -80661
rect -49173 -80705 -49117 -80661
rect -49073 -80705 -49017 -80661
rect -48973 -80705 -48917 -80661
rect -48873 -80705 -48817 -80661
rect -48773 -80705 -48717 -80661
rect -48673 -80705 -48617 -80661
rect -48573 -80705 -48517 -80661
rect -48473 -80705 -48017 -80661
rect -47973 -80705 -47917 -80661
rect -47873 -80705 -47817 -80661
rect -47773 -80705 -47717 -80661
rect -47673 -80705 -47617 -80661
rect -47573 -80705 -47517 -80661
rect -47473 -80705 -47417 -80661
rect -47373 -80705 -47317 -80661
rect -47273 -80705 -47217 -80661
rect -47173 -80705 -47117 -80661
rect -47073 -80705 -47017 -80661
rect -46973 -80705 -46917 -80661
rect -46873 -80705 -46817 -80661
rect -46773 -80705 -46717 -80661
rect -46673 -80705 -46617 -80661
rect -46573 -80705 -46517 -80661
rect -46473 -80705 -46017 -80661
rect -45973 -80705 -45917 -80661
rect -45873 -80705 -45817 -80661
rect -45773 -80705 -45717 -80661
rect -45673 -80705 -45617 -80661
rect -45573 -80705 -45517 -80661
rect -45473 -80705 -45417 -80661
rect -45373 -80705 -45317 -80661
rect -45273 -80705 -45217 -80661
rect -45173 -80705 -45117 -80661
rect -45073 -80705 -45017 -80661
rect -44973 -80705 -44917 -80661
rect -44873 -80705 -44817 -80661
rect -44773 -80705 -44717 -80661
rect -44673 -80705 -44617 -80661
rect -44573 -80705 -44517 -80661
rect -44473 -80705 -44017 -80661
rect -43973 -80705 -43917 -80661
rect -43873 -80705 -43817 -80661
rect -43773 -80705 -43717 -80661
rect -43673 -80705 -43617 -80661
rect -43573 -80705 -43517 -80661
rect -43473 -80705 -43417 -80661
rect -43373 -80705 -43317 -80661
rect -43273 -80705 -43217 -80661
rect -43173 -80705 -43117 -80661
rect -43073 -80705 -43017 -80661
rect -42973 -80705 -42917 -80661
rect -42873 -80705 -42817 -80661
rect -42773 -80705 -42717 -80661
rect -42673 -80705 -42617 -80661
rect -42573 -80705 -42517 -80661
rect -42473 -80699 80737 -80661
rect 80781 -80699 80837 -80655
rect 80881 -80699 80937 -80655
rect 80981 -80699 81037 -80655
rect 81081 -80699 81137 -80655
rect 81181 -80699 81237 -80655
rect 81281 -80699 81337 -80655
rect 81381 -80699 81437 -80655
rect 81481 -80699 81537 -80655
rect 81581 -80699 81637 -80655
rect 81681 -80699 81737 -80655
rect 81781 -80699 81837 -80655
rect 81881 -80699 81937 -80655
rect 81981 -80699 82037 -80655
rect 82081 -80699 82137 -80655
rect 82181 -80699 82237 -80655
rect 82281 -80699 82737 -80655
rect 82781 -80699 82837 -80655
rect 82881 -80699 82937 -80655
rect 82981 -80699 83037 -80655
rect 83081 -80699 83137 -80655
rect 83181 -80699 83237 -80655
rect 83281 -80699 83337 -80655
rect 83381 -80699 83437 -80655
rect 83481 -80699 83537 -80655
rect 83581 -80699 83637 -80655
rect 83681 -80699 83737 -80655
rect 83781 -80699 83837 -80655
rect 83881 -80699 83937 -80655
rect 83981 -80699 84037 -80655
rect 84081 -80699 84137 -80655
rect 84181 -80699 84237 -80655
rect 84281 -80699 84737 -80655
rect 84781 -80699 84837 -80655
rect 84881 -80699 84937 -80655
rect 84981 -80699 85037 -80655
rect 85081 -80699 85137 -80655
rect 85181 -80699 85237 -80655
rect 85281 -80699 85337 -80655
rect 85381 -80699 85437 -80655
rect 85481 -80699 85537 -80655
rect 85581 -80699 85637 -80655
rect 85681 -80699 85737 -80655
rect 85781 -80699 85837 -80655
rect 85881 -80699 85937 -80655
rect 85981 -80699 86037 -80655
rect 86081 -80699 86137 -80655
rect 86181 -80699 86237 -80655
rect 86281 -80699 86737 -80655
rect 86781 -80699 86837 -80655
rect 86881 -80699 86937 -80655
rect 86981 -80699 87037 -80655
rect 87081 -80699 87137 -80655
rect 87181 -80699 87237 -80655
rect 87281 -80699 87337 -80655
rect 87381 -80699 87437 -80655
rect 87481 -80699 87537 -80655
rect 87581 -80699 87637 -80655
rect 87681 -80699 87737 -80655
rect 87781 -80699 87837 -80655
rect 87881 -80699 87937 -80655
rect 87981 -80699 88037 -80655
rect 88081 -80699 88137 -80655
rect 88181 -80699 88237 -80655
rect 88281 -80699 177360 -80655
rect -42473 -80705 177360 -80699
rect -109116 -80755 177360 -80705
rect -109116 -80759 80737 -80755
rect -109116 -80803 -82968 -80759
rect -82924 -80803 -82868 -80759
rect -82824 -80803 -82768 -80759
rect -82724 -80803 -82668 -80759
rect -82624 -80803 -82568 -80759
rect -82524 -80803 -82468 -80759
rect -82424 -80803 -82368 -80759
rect -82324 -80803 -82268 -80759
rect -82224 -80803 -82168 -80759
rect -82124 -80803 -82068 -80759
rect -82024 -80803 -81968 -80759
rect -81924 -80803 -81868 -80759
rect -81824 -80803 -81768 -80759
rect -81724 -80803 -81668 -80759
rect -81624 -80803 -81568 -80759
rect -81524 -80803 -81468 -80759
rect -81424 -80803 -80968 -80759
rect -80924 -80803 -80868 -80759
rect -80824 -80803 -80768 -80759
rect -80724 -80803 -80668 -80759
rect -80624 -80803 -80568 -80759
rect -80524 -80803 -80468 -80759
rect -80424 -80803 -80368 -80759
rect -80324 -80803 -80268 -80759
rect -80224 -80803 -80168 -80759
rect -80124 -80803 -80068 -80759
rect -80024 -80803 -79968 -80759
rect -79924 -80803 -79868 -80759
rect -79824 -80803 -79768 -80759
rect -79724 -80803 -79668 -80759
rect -79624 -80803 -79568 -80759
rect -79524 -80803 -79468 -80759
rect -79424 -80803 -78968 -80759
rect -78924 -80803 -78868 -80759
rect -78824 -80803 -78768 -80759
rect -78724 -80803 -78668 -80759
rect -78624 -80803 -78568 -80759
rect -78524 -80803 -78468 -80759
rect -78424 -80803 -78368 -80759
rect -78324 -80803 -78268 -80759
rect -78224 -80803 -78168 -80759
rect -78124 -80803 -78068 -80759
rect -78024 -80803 -77968 -80759
rect -77924 -80803 -77868 -80759
rect -77824 -80803 -77768 -80759
rect -77724 -80803 -77668 -80759
rect -77624 -80803 -77568 -80759
rect -77524 -80803 -77468 -80759
rect -77424 -80803 -76968 -80759
rect -76924 -80803 -76868 -80759
rect -76824 -80803 -76768 -80759
rect -76724 -80803 -76668 -80759
rect -76624 -80803 -76568 -80759
rect -76524 -80803 -76468 -80759
rect -76424 -80803 -76368 -80759
rect -76324 -80803 -76268 -80759
rect -76224 -80803 -76168 -80759
rect -76124 -80803 -76068 -80759
rect -76024 -80803 -75968 -80759
rect -75924 -80803 -75868 -80759
rect -75824 -80803 -75768 -80759
rect -75724 -80803 -75668 -80759
rect -75624 -80803 -75568 -80759
rect -75524 -80803 -75468 -80759
rect -75424 -80761 80737 -80759
rect -75424 -80803 -50017 -80761
rect -109116 -80805 -50017 -80803
rect -49973 -80805 -49917 -80761
rect -49873 -80805 -49817 -80761
rect -49773 -80805 -49717 -80761
rect -49673 -80805 -49617 -80761
rect -49573 -80805 -49517 -80761
rect -49473 -80805 -49417 -80761
rect -49373 -80805 -49317 -80761
rect -49273 -80805 -49217 -80761
rect -49173 -80805 -49117 -80761
rect -49073 -80805 -49017 -80761
rect -48973 -80805 -48917 -80761
rect -48873 -80805 -48817 -80761
rect -48773 -80805 -48717 -80761
rect -48673 -80805 -48617 -80761
rect -48573 -80805 -48517 -80761
rect -48473 -80805 -48017 -80761
rect -47973 -80805 -47917 -80761
rect -47873 -80805 -47817 -80761
rect -47773 -80805 -47717 -80761
rect -47673 -80805 -47617 -80761
rect -47573 -80805 -47517 -80761
rect -47473 -80805 -47417 -80761
rect -47373 -80805 -47317 -80761
rect -47273 -80805 -47217 -80761
rect -47173 -80805 -47117 -80761
rect -47073 -80805 -47017 -80761
rect -46973 -80805 -46917 -80761
rect -46873 -80805 -46817 -80761
rect -46773 -80805 -46717 -80761
rect -46673 -80805 -46617 -80761
rect -46573 -80805 -46517 -80761
rect -46473 -80805 -46017 -80761
rect -45973 -80805 -45917 -80761
rect -45873 -80805 -45817 -80761
rect -45773 -80805 -45717 -80761
rect -45673 -80805 -45617 -80761
rect -45573 -80805 -45517 -80761
rect -45473 -80805 -45417 -80761
rect -45373 -80805 -45317 -80761
rect -45273 -80805 -45217 -80761
rect -45173 -80805 -45117 -80761
rect -45073 -80805 -45017 -80761
rect -44973 -80805 -44917 -80761
rect -44873 -80805 -44817 -80761
rect -44773 -80805 -44717 -80761
rect -44673 -80805 -44617 -80761
rect -44573 -80805 -44517 -80761
rect -44473 -80805 -44017 -80761
rect -43973 -80805 -43917 -80761
rect -43873 -80805 -43817 -80761
rect -43773 -80805 -43717 -80761
rect -43673 -80805 -43617 -80761
rect -43573 -80805 -43517 -80761
rect -43473 -80805 -43417 -80761
rect -43373 -80805 -43317 -80761
rect -43273 -80805 -43217 -80761
rect -43173 -80805 -43117 -80761
rect -43073 -80805 -43017 -80761
rect -42973 -80805 -42917 -80761
rect -42873 -80805 -42817 -80761
rect -42773 -80805 -42717 -80761
rect -42673 -80805 -42617 -80761
rect -42573 -80805 -42517 -80761
rect -42473 -80799 80737 -80761
rect 80781 -80799 80837 -80755
rect 80881 -80799 80937 -80755
rect 80981 -80799 81037 -80755
rect 81081 -80799 81137 -80755
rect 81181 -80799 81237 -80755
rect 81281 -80799 81337 -80755
rect 81381 -80799 81437 -80755
rect 81481 -80799 81537 -80755
rect 81581 -80799 81637 -80755
rect 81681 -80799 81737 -80755
rect 81781 -80799 81837 -80755
rect 81881 -80799 81937 -80755
rect 81981 -80799 82037 -80755
rect 82081 -80799 82137 -80755
rect 82181 -80799 82237 -80755
rect 82281 -80799 82737 -80755
rect 82781 -80799 82837 -80755
rect 82881 -80799 82937 -80755
rect 82981 -80799 83037 -80755
rect 83081 -80799 83137 -80755
rect 83181 -80799 83237 -80755
rect 83281 -80799 83337 -80755
rect 83381 -80799 83437 -80755
rect 83481 -80799 83537 -80755
rect 83581 -80799 83637 -80755
rect 83681 -80799 83737 -80755
rect 83781 -80799 83837 -80755
rect 83881 -80799 83937 -80755
rect 83981 -80799 84037 -80755
rect 84081 -80799 84137 -80755
rect 84181 -80799 84237 -80755
rect 84281 -80799 84737 -80755
rect 84781 -80799 84837 -80755
rect 84881 -80799 84937 -80755
rect 84981 -80799 85037 -80755
rect 85081 -80799 85137 -80755
rect 85181 -80799 85237 -80755
rect 85281 -80799 85337 -80755
rect 85381 -80799 85437 -80755
rect 85481 -80799 85537 -80755
rect 85581 -80799 85637 -80755
rect 85681 -80799 85737 -80755
rect 85781 -80799 85837 -80755
rect 85881 -80799 85937 -80755
rect 85981 -80799 86037 -80755
rect 86081 -80799 86137 -80755
rect 86181 -80799 86237 -80755
rect 86281 -80799 86737 -80755
rect 86781 -80799 86837 -80755
rect 86881 -80799 86937 -80755
rect 86981 -80799 87037 -80755
rect 87081 -80799 87137 -80755
rect 87181 -80799 87237 -80755
rect 87281 -80799 87337 -80755
rect 87381 -80799 87437 -80755
rect 87481 -80799 87537 -80755
rect 87581 -80799 87637 -80755
rect 87681 -80799 87737 -80755
rect 87781 -80799 87837 -80755
rect 87881 -80799 87937 -80755
rect 87981 -80799 88037 -80755
rect 88081 -80799 88137 -80755
rect 88181 -80799 88237 -80755
rect 88281 -80799 177360 -80755
rect -42473 -80805 177360 -80799
rect -109116 -80855 177360 -80805
rect -109116 -80859 80737 -80855
rect -109116 -80903 -82968 -80859
rect -82924 -80903 -82868 -80859
rect -82824 -80903 -82768 -80859
rect -82724 -80903 -82668 -80859
rect -82624 -80903 -82568 -80859
rect -82524 -80903 -82468 -80859
rect -82424 -80903 -82368 -80859
rect -82324 -80903 -82268 -80859
rect -82224 -80903 -82168 -80859
rect -82124 -80903 -82068 -80859
rect -82024 -80903 -81968 -80859
rect -81924 -80903 -81868 -80859
rect -81824 -80903 -81768 -80859
rect -81724 -80903 -81668 -80859
rect -81624 -80903 -81568 -80859
rect -81524 -80903 -81468 -80859
rect -81424 -80903 -80968 -80859
rect -80924 -80903 -80868 -80859
rect -80824 -80903 -80768 -80859
rect -80724 -80903 -80668 -80859
rect -80624 -80903 -80568 -80859
rect -80524 -80903 -80468 -80859
rect -80424 -80903 -80368 -80859
rect -80324 -80903 -80268 -80859
rect -80224 -80903 -80168 -80859
rect -80124 -80903 -80068 -80859
rect -80024 -80903 -79968 -80859
rect -79924 -80903 -79868 -80859
rect -79824 -80903 -79768 -80859
rect -79724 -80903 -79668 -80859
rect -79624 -80903 -79568 -80859
rect -79524 -80903 -79468 -80859
rect -79424 -80903 -78968 -80859
rect -78924 -80903 -78868 -80859
rect -78824 -80903 -78768 -80859
rect -78724 -80903 -78668 -80859
rect -78624 -80903 -78568 -80859
rect -78524 -80903 -78468 -80859
rect -78424 -80903 -78368 -80859
rect -78324 -80903 -78268 -80859
rect -78224 -80903 -78168 -80859
rect -78124 -80903 -78068 -80859
rect -78024 -80903 -77968 -80859
rect -77924 -80903 -77868 -80859
rect -77824 -80903 -77768 -80859
rect -77724 -80903 -77668 -80859
rect -77624 -80903 -77568 -80859
rect -77524 -80903 -77468 -80859
rect -77424 -80903 -76968 -80859
rect -76924 -80903 -76868 -80859
rect -76824 -80903 -76768 -80859
rect -76724 -80903 -76668 -80859
rect -76624 -80903 -76568 -80859
rect -76524 -80903 -76468 -80859
rect -76424 -80903 -76368 -80859
rect -76324 -80903 -76268 -80859
rect -76224 -80903 -76168 -80859
rect -76124 -80903 -76068 -80859
rect -76024 -80903 -75968 -80859
rect -75924 -80903 -75868 -80859
rect -75824 -80903 -75768 -80859
rect -75724 -80903 -75668 -80859
rect -75624 -80903 -75568 -80859
rect -75524 -80903 -75468 -80859
rect -75424 -80861 80737 -80859
rect -75424 -80903 -50017 -80861
rect -109116 -80905 -50017 -80903
rect -49973 -80905 -49917 -80861
rect -49873 -80905 -49817 -80861
rect -49773 -80905 -49717 -80861
rect -49673 -80905 -49617 -80861
rect -49573 -80905 -49517 -80861
rect -49473 -80905 -49417 -80861
rect -49373 -80905 -49317 -80861
rect -49273 -80905 -49217 -80861
rect -49173 -80905 -49117 -80861
rect -49073 -80905 -49017 -80861
rect -48973 -80905 -48917 -80861
rect -48873 -80905 -48817 -80861
rect -48773 -80905 -48717 -80861
rect -48673 -80905 -48617 -80861
rect -48573 -80905 -48517 -80861
rect -48473 -80905 -48017 -80861
rect -47973 -80905 -47917 -80861
rect -47873 -80905 -47817 -80861
rect -47773 -80905 -47717 -80861
rect -47673 -80905 -47617 -80861
rect -47573 -80905 -47517 -80861
rect -47473 -80905 -47417 -80861
rect -47373 -80905 -47317 -80861
rect -47273 -80905 -47217 -80861
rect -47173 -80905 -47117 -80861
rect -47073 -80905 -47017 -80861
rect -46973 -80905 -46917 -80861
rect -46873 -80905 -46817 -80861
rect -46773 -80905 -46717 -80861
rect -46673 -80905 -46617 -80861
rect -46573 -80905 -46517 -80861
rect -46473 -80905 -46017 -80861
rect -45973 -80905 -45917 -80861
rect -45873 -80905 -45817 -80861
rect -45773 -80905 -45717 -80861
rect -45673 -80905 -45617 -80861
rect -45573 -80905 -45517 -80861
rect -45473 -80905 -45417 -80861
rect -45373 -80905 -45317 -80861
rect -45273 -80905 -45217 -80861
rect -45173 -80905 -45117 -80861
rect -45073 -80905 -45017 -80861
rect -44973 -80905 -44917 -80861
rect -44873 -80905 -44817 -80861
rect -44773 -80905 -44717 -80861
rect -44673 -80905 -44617 -80861
rect -44573 -80905 -44517 -80861
rect -44473 -80905 -44017 -80861
rect -43973 -80905 -43917 -80861
rect -43873 -80905 -43817 -80861
rect -43773 -80905 -43717 -80861
rect -43673 -80905 -43617 -80861
rect -43573 -80905 -43517 -80861
rect -43473 -80905 -43417 -80861
rect -43373 -80905 -43317 -80861
rect -43273 -80905 -43217 -80861
rect -43173 -80905 -43117 -80861
rect -43073 -80905 -43017 -80861
rect -42973 -80905 -42917 -80861
rect -42873 -80905 -42817 -80861
rect -42773 -80905 -42717 -80861
rect -42673 -80905 -42617 -80861
rect -42573 -80905 -42517 -80861
rect -42473 -80899 80737 -80861
rect 80781 -80899 80837 -80855
rect 80881 -80899 80937 -80855
rect 80981 -80899 81037 -80855
rect 81081 -80899 81137 -80855
rect 81181 -80899 81237 -80855
rect 81281 -80899 81337 -80855
rect 81381 -80899 81437 -80855
rect 81481 -80899 81537 -80855
rect 81581 -80899 81637 -80855
rect 81681 -80899 81737 -80855
rect 81781 -80899 81837 -80855
rect 81881 -80899 81937 -80855
rect 81981 -80899 82037 -80855
rect 82081 -80899 82137 -80855
rect 82181 -80899 82237 -80855
rect 82281 -80899 82737 -80855
rect 82781 -80899 82837 -80855
rect 82881 -80899 82937 -80855
rect 82981 -80899 83037 -80855
rect 83081 -80899 83137 -80855
rect 83181 -80899 83237 -80855
rect 83281 -80899 83337 -80855
rect 83381 -80899 83437 -80855
rect 83481 -80899 83537 -80855
rect 83581 -80899 83637 -80855
rect 83681 -80899 83737 -80855
rect 83781 -80899 83837 -80855
rect 83881 -80899 83937 -80855
rect 83981 -80899 84037 -80855
rect 84081 -80899 84137 -80855
rect 84181 -80899 84237 -80855
rect 84281 -80899 84737 -80855
rect 84781 -80899 84837 -80855
rect 84881 -80899 84937 -80855
rect 84981 -80899 85037 -80855
rect 85081 -80899 85137 -80855
rect 85181 -80899 85237 -80855
rect 85281 -80899 85337 -80855
rect 85381 -80899 85437 -80855
rect 85481 -80899 85537 -80855
rect 85581 -80899 85637 -80855
rect 85681 -80899 85737 -80855
rect 85781 -80899 85837 -80855
rect 85881 -80899 85937 -80855
rect 85981 -80899 86037 -80855
rect 86081 -80899 86137 -80855
rect 86181 -80899 86237 -80855
rect 86281 -80899 86737 -80855
rect 86781 -80899 86837 -80855
rect 86881 -80899 86937 -80855
rect 86981 -80899 87037 -80855
rect 87081 -80899 87137 -80855
rect 87181 -80899 87237 -80855
rect 87281 -80899 87337 -80855
rect 87381 -80899 87437 -80855
rect 87481 -80899 87537 -80855
rect 87581 -80899 87637 -80855
rect 87681 -80899 87737 -80855
rect 87781 -80899 87837 -80855
rect 87881 -80899 87937 -80855
rect 87981 -80899 88037 -80855
rect 88081 -80899 88137 -80855
rect 88181 -80899 88237 -80855
rect 88281 -80899 177360 -80855
rect -42473 -80905 177360 -80899
rect -109116 -80955 177360 -80905
rect -109116 -80959 80737 -80955
rect -109116 -81003 -82968 -80959
rect -82924 -81003 -82868 -80959
rect -82824 -81003 -82768 -80959
rect -82724 -81003 -82668 -80959
rect -82624 -81003 -82568 -80959
rect -82524 -81003 -82468 -80959
rect -82424 -81003 -82368 -80959
rect -82324 -81003 -82268 -80959
rect -82224 -81003 -82168 -80959
rect -82124 -81003 -82068 -80959
rect -82024 -81003 -81968 -80959
rect -81924 -81003 -81868 -80959
rect -81824 -81003 -81768 -80959
rect -81724 -81003 -81668 -80959
rect -81624 -81003 -81568 -80959
rect -81524 -81003 -81468 -80959
rect -81424 -81003 -80968 -80959
rect -80924 -81003 -80868 -80959
rect -80824 -81003 -80768 -80959
rect -80724 -81003 -80668 -80959
rect -80624 -81003 -80568 -80959
rect -80524 -81003 -80468 -80959
rect -80424 -81003 -80368 -80959
rect -80324 -81003 -80268 -80959
rect -80224 -81003 -80168 -80959
rect -80124 -81003 -80068 -80959
rect -80024 -81003 -79968 -80959
rect -79924 -81003 -79868 -80959
rect -79824 -81003 -79768 -80959
rect -79724 -81003 -79668 -80959
rect -79624 -81003 -79568 -80959
rect -79524 -81003 -79468 -80959
rect -79424 -81003 -78968 -80959
rect -78924 -81003 -78868 -80959
rect -78824 -81003 -78768 -80959
rect -78724 -81003 -78668 -80959
rect -78624 -81003 -78568 -80959
rect -78524 -81003 -78468 -80959
rect -78424 -81003 -78368 -80959
rect -78324 -81003 -78268 -80959
rect -78224 -81003 -78168 -80959
rect -78124 -81003 -78068 -80959
rect -78024 -81003 -77968 -80959
rect -77924 -81003 -77868 -80959
rect -77824 -81003 -77768 -80959
rect -77724 -81003 -77668 -80959
rect -77624 -81003 -77568 -80959
rect -77524 -81003 -77468 -80959
rect -77424 -81003 -76968 -80959
rect -76924 -81003 -76868 -80959
rect -76824 -81003 -76768 -80959
rect -76724 -81003 -76668 -80959
rect -76624 -81003 -76568 -80959
rect -76524 -81003 -76468 -80959
rect -76424 -81003 -76368 -80959
rect -76324 -81003 -76268 -80959
rect -76224 -81003 -76168 -80959
rect -76124 -81003 -76068 -80959
rect -76024 -81003 -75968 -80959
rect -75924 -81003 -75868 -80959
rect -75824 -81003 -75768 -80959
rect -75724 -81003 -75668 -80959
rect -75624 -81003 -75568 -80959
rect -75524 -81003 -75468 -80959
rect -75424 -80961 80737 -80959
rect -75424 -81003 -50017 -80961
rect -109116 -81005 -50017 -81003
rect -49973 -81005 -49917 -80961
rect -49873 -81005 -49817 -80961
rect -49773 -81005 -49717 -80961
rect -49673 -81005 -49617 -80961
rect -49573 -81005 -49517 -80961
rect -49473 -81005 -49417 -80961
rect -49373 -81005 -49317 -80961
rect -49273 -81005 -49217 -80961
rect -49173 -81005 -49117 -80961
rect -49073 -81005 -49017 -80961
rect -48973 -81005 -48917 -80961
rect -48873 -81005 -48817 -80961
rect -48773 -81005 -48717 -80961
rect -48673 -81005 -48617 -80961
rect -48573 -81005 -48517 -80961
rect -48473 -81005 -48017 -80961
rect -47973 -81005 -47917 -80961
rect -47873 -81005 -47817 -80961
rect -47773 -81005 -47717 -80961
rect -47673 -81005 -47617 -80961
rect -47573 -81005 -47517 -80961
rect -47473 -81005 -47417 -80961
rect -47373 -81005 -47317 -80961
rect -47273 -81005 -47217 -80961
rect -47173 -81005 -47117 -80961
rect -47073 -81005 -47017 -80961
rect -46973 -81005 -46917 -80961
rect -46873 -81005 -46817 -80961
rect -46773 -81005 -46717 -80961
rect -46673 -81005 -46617 -80961
rect -46573 -81005 -46517 -80961
rect -46473 -81005 -46017 -80961
rect -45973 -81005 -45917 -80961
rect -45873 -81005 -45817 -80961
rect -45773 -81005 -45717 -80961
rect -45673 -81005 -45617 -80961
rect -45573 -81005 -45517 -80961
rect -45473 -81005 -45417 -80961
rect -45373 -81005 -45317 -80961
rect -45273 -81005 -45217 -80961
rect -45173 -81005 -45117 -80961
rect -45073 -81005 -45017 -80961
rect -44973 -81005 -44917 -80961
rect -44873 -81005 -44817 -80961
rect -44773 -81005 -44717 -80961
rect -44673 -81005 -44617 -80961
rect -44573 -81005 -44517 -80961
rect -44473 -81005 -44017 -80961
rect -43973 -81005 -43917 -80961
rect -43873 -81005 -43817 -80961
rect -43773 -81005 -43717 -80961
rect -43673 -81005 -43617 -80961
rect -43573 -81005 -43517 -80961
rect -43473 -81005 -43417 -80961
rect -43373 -81005 -43317 -80961
rect -43273 -81005 -43217 -80961
rect -43173 -81005 -43117 -80961
rect -43073 -81005 -43017 -80961
rect -42973 -81005 -42917 -80961
rect -42873 -81005 -42817 -80961
rect -42773 -81005 -42717 -80961
rect -42673 -81005 -42617 -80961
rect -42573 -81005 -42517 -80961
rect -42473 -80999 80737 -80961
rect 80781 -80999 80837 -80955
rect 80881 -80999 80937 -80955
rect 80981 -80999 81037 -80955
rect 81081 -80999 81137 -80955
rect 81181 -80999 81237 -80955
rect 81281 -80999 81337 -80955
rect 81381 -80999 81437 -80955
rect 81481 -80999 81537 -80955
rect 81581 -80999 81637 -80955
rect 81681 -80999 81737 -80955
rect 81781 -80999 81837 -80955
rect 81881 -80999 81937 -80955
rect 81981 -80999 82037 -80955
rect 82081 -80999 82137 -80955
rect 82181 -80999 82237 -80955
rect 82281 -80999 82737 -80955
rect 82781 -80999 82837 -80955
rect 82881 -80999 82937 -80955
rect 82981 -80999 83037 -80955
rect 83081 -80999 83137 -80955
rect 83181 -80999 83237 -80955
rect 83281 -80999 83337 -80955
rect 83381 -80999 83437 -80955
rect 83481 -80999 83537 -80955
rect 83581 -80999 83637 -80955
rect 83681 -80999 83737 -80955
rect 83781 -80999 83837 -80955
rect 83881 -80999 83937 -80955
rect 83981 -80999 84037 -80955
rect 84081 -80999 84137 -80955
rect 84181 -80999 84237 -80955
rect 84281 -80999 84737 -80955
rect 84781 -80999 84837 -80955
rect 84881 -80999 84937 -80955
rect 84981 -80999 85037 -80955
rect 85081 -80999 85137 -80955
rect 85181 -80999 85237 -80955
rect 85281 -80999 85337 -80955
rect 85381 -80999 85437 -80955
rect 85481 -80999 85537 -80955
rect 85581 -80999 85637 -80955
rect 85681 -80999 85737 -80955
rect 85781 -80999 85837 -80955
rect 85881 -80999 85937 -80955
rect 85981 -80999 86037 -80955
rect 86081 -80999 86137 -80955
rect 86181 -80999 86237 -80955
rect 86281 -80999 86737 -80955
rect 86781 -80999 86837 -80955
rect 86881 -80999 86937 -80955
rect 86981 -80999 87037 -80955
rect 87081 -80999 87137 -80955
rect 87181 -80999 87237 -80955
rect 87281 -80999 87337 -80955
rect 87381 -80999 87437 -80955
rect 87481 -80999 87537 -80955
rect 87581 -80999 87637 -80955
rect 87681 -80999 87737 -80955
rect 87781 -80999 87837 -80955
rect 87881 -80999 87937 -80955
rect 87981 -80999 88037 -80955
rect 88081 -80999 88137 -80955
rect 88181 -80999 88237 -80955
rect 88281 -80999 177360 -80955
rect -42473 -81005 177360 -80999
rect -109116 -81055 177360 -81005
rect -109116 -81059 80737 -81055
rect -109116 -81103 -82968 -81059
rect -82924 -81103 -82868 -81059
rect -82824 -81103 -82768 -81059
rect -82724 -81103 -82668 -81059
rect -82624 -81103 -82568 -81059
rect -82524 -81103 -82468 -81059
rect -82424 -81103 -82368 -81059
rect -82324 -81103 -82268 -81059
rect -82224 -81103 -82168 -81059
rect -82124 -81103 -82068 -81059
rect -82024 -81103 -81968 -81059
rect -81924 -81103 -81868 -81059
rect -81824 -81103 -81768 -81059
rect -81724 -81103 -81668 -81059
rect -81624 -81103 -81568 -81059
rect -81524 -81103 -81468 -81059
rect -81424 -81103 -80968 -81059
rect -80924 -81103 -80868 -81059
rect -80824 -81103 -80768 -81059
rect -80724 -81103 -80668 -81059
rect -80624 -81103 -80568 -81059
rect -80524 -81103 -80468 -81059
rect -80424 -81103 -80368 -81059
rect -80324 -81103 -80268 -81059
rect -80224 -81103 -80168 -81059
rect -80124 -81103 -80068 -81059
rect -80024 -81103 -79968 -81059
rect -79924 -81103 -79868 -81059
rect -79824 -81103 -79768 -81059
rect -79724 -81103 -79668 -81059
rect -79624 -81103 -79568 -81059
rect -79524 -81103 -79468 -81059
rect -79424 -81103 -78968 -81059
rect -78924 -81103 -78868 -81059
rect -78824 -81103 -78768 -81059
rect -78724 -81103 -78668 -81059
rect -78624 -81103 -78568 -81059
rect -78524 -81103 -78468 -81059
rect -78424 -81103 -78368 -81059
rect -78324 -81103 -78268 -81059
rect -78224 -81103 -78168 -81059
rect -78124 -81103 -78068 -81059
rect -78024 -81103 -77968 -81059
rect -77924 -81103 -77868 -81059
rect -77824 -81103 -77768 -81059
rect -77724 -81103 -77668 -81059
rect -77624 -81103 -77568 -81059
rect -77524 -81103 -77468 -81059
rect -77424 -81103 -76968 -81059
rect -76924 -81103 -76868 -81059
rect -76824 -81103 -76768 -81059
rect -76724 -81103 -76668 -81059
rect -76624 -81103 -76568 -81059
rect -76524 -81103 -76468 -81059
rect -76424 -81103 -76368 -81059
rect -76324 -81103 -76268 -81059
rect -76224 -81103 -76168 -81059
rect -76124 -81103 -76068 -81059
rect -76024 -81103 -75968 -81059
rect -75924 -81103 -75868 -81059
rect -75824 -81103 -75768 -81059
rect -75724 -81103 -75668 -81059
rect -75624 -81103 -75568 -81059
rect -75524 -81103 -75468 -81059
rect -75424 -81061 80737 -81059
rect -75424 -81103 -50017 -81061
rect -109116 -81105 -50017 -81103
rect -49973 -81105 -49917 -81061
rect -49873 -81105 -49817 -81061
rect -49773 -81105 -49717 -81061
rect -49673 -81105 -49617 -81061
rect -49573 -81105 -49517 -81061
rect -49473 -81105 -49417 -81061
rect -49373 -81105 -49317 -81061
rect -49273 -81105 -49217 -81061
rect -49173 -81105 -49117 -81061
rect -49073 -81105 -49017 -81061
rect -48973 -81105 -48917 -81061
rect -48873 -81105 -48817 -81061
rect -48773 -81105 -48717 -81061
rect -48673 -81105 -48617 -81061
rect -48573 -81105 -48517 -81061
rect -48473 -81105 -48017 -81061
rect -47973 -81105 -47917 -81061
rect -47873 -81105 -47817 -81061
rect -47773 -81105 -47717 -81061
rect -47673 -81105 -47617 -81061
rect -47573 -81105 -47517 -81061
rect -47473 -81105 -47417 -81061
rect -47373 -81105 -47317 -81061
rect -47273 -81105 -47217 -81061
rect -47173 -81105 -47117 -81061
rect -47073 -81105 -47017 -81061
rect -46973 -81105 -46917 -81061
rect -46873 -81105 -46817 -81061
rect -46773 -81105 -46717 -81061
rect -46673 -81105 -46617 -81061
rect -46573 -81105 -46517 -81061
rect -46473 -81105 -46017 -81061
rect -45973 -81105 -45917 -81061
rect -45873 -81105 -45817 -81061
rect -45773 -81105 -45717 -81061
rect -45673 -81105 -45617 -81061
rect -45573 -81105 -45517 -81061
rect -45473 -81105 -45417 -81061
rect -45373 -81105 -45317 -81061
rect -45273 -81105 -45217 -81061
rect -45173 -81105 -45117 -81061
rect -45073 -81105 -45017 -81061
rect -44973 -81105 -44917 -81061
rect -44873 -81105 -44817 -81061
rect -44773 -81105 -44717 -81061
rect -44673 -81105 -44617 -81061
rect -44573 -81105 -44517 -81061
rect -44473 -81105 -44017 -81061
rect -43973 -81105 -43917 -81061
rect -43873 -81105 -43817 -81061
rect -43773 -81105 -43717 -81061
rect -43673 -81105 -43617 -81061
rect -43573 -81105 -43517 -81061
rect -43473 -81105 -43417 -81061
rect -43373 -81105 -43317 -81061
rect -43273 -81105 -43217 -81061
rect -43173 -81105 -43117 -81061
rect -43073 -81105 -43017 -81061
rect -42973 -81105 -42917 -81061
rect -42873 -81105 -42817 -81061
rect -42773 -81105 -42717 -81061
rect -42673 -81105 -42617 -81061
rect -42573 -81105 -42517 -81061
rect -42473 -81099 80737 -81061
rect 80781 -81099 80837 -81055
rect 80881 -81099 80937 -81055
rect 80981 -81099 81037 -81055
rect 81081 -81099 81137 -81055
rect 81181 -81099 81237 -81055
rect 81281 -81099 81337 -81055
rect 81381 -81099 81437 -81055
rect 81481 -81099 81537 -81055
rect 81581 -81099 81637 -81055
rect 81681 -81099 81737 -81055
rect 81781 -81099 81837 -81055
rect 81881 -81099 81937 -81055
rect 81981 -81099 82037 -81055
rect 82081 -81099 82137 -81055
rect 82181 -81099 82237 -81055
rect 82281 -81099 82737 -81055
rect 82781 -81099 82837 -81055
rect 82881 -81099 82937 -81055
rect 82981 -81099 83037 -81055
rect 83081 -81099 83137 -81055
rect 83181 -81099 83237 -81055
rect 83281 -81099 83337 -81055
rect 83381 -81099 83437 -81055
rect 83481 -81099 83537 -81055
rect 83581 -81099 83637 -81055
rect 83681 -81099 83737 -81055
rect 83781 -81099 83837 -81055
rect 83881 -81099 83937 -81055
rect 83981 -81099 84037 -81055
rect 84081 -81099 84137 -81055
rect 84181 -81099 84237 -81055
rect 84281 -81099 84737 -81055
rect 84781 -81099 84837 -81055
rect 84881 -81099 84937 -81055
rect 84981 -81099 85037 -81055
rect 85081 -81099 85137 -81055
rect 85181 -81099 85237 -81055
rect 85281 -81099 85337 -81055
rect 85381 -81099 85437 -81055
rect 85481 -81099 85537 -81055
rect 85581 -81099 85637 -81055
rect 85681 -81099 85737 -81055
rect 85781 -81099 85837 -81055
rect 85881 -81099 85937 -81055
rect 85981 -81099 86037 -81055
rect 86081 -81099 86137 -81055
rect 86181 -81099 86237 -81055
rect 86281 -81099 86737 -81055
rect 86781 -81099 86837 -81055
rect 86881 -81099 86937 -81055
rect 86981 -81099 87037 -81055
rect 87081 -81099 87137 -81055
rect 87181 -81099 87237 -81055
rect 87281 -81099 87337 -81055
rect 87381 -81099 87437 -81055
rect 87481 -81099 87537 -81055
rect 87581 -81099 87637 -81055
rect 87681 -81099 87737 -81055
rect 87781 -81099 87837 -81055
rect 87881 -81099 87937 -81055
rect 87981 -81099 88037 -81055
rect 88081 -81099 88137 -81055
rect 88181 -81099 88237 -81055
rect 88281 -81099 177360 -81055
rect -42473 -81105 177360 -81099
rect -109116 -81155 177360 -81105
rect -109116 -81159 80737 -81155
rect -109116 -81203 -82968 -81159
rect -82924 -81203 -82868 -81159
rect -82824 -81203 -82768 -81159
rect -82724 -81203 -82668 -81159
rect -82624 -81203 -82568 -81159
rect -82524 -81203 -82468 -81159
rect -82424 -81203 -82368 -81159
rect -82324 -81203 -82268 -81159
rect -82224 -81203 -82168 -81159
rect -82124 -81203 -82068 -81159
rect -82024 -81203 -81968 -81159
rect -81924 -81203 -81868 -81159
rect -81824 -81203 -81768 -81159
rect -81724 -81203 -81668 -81159
rect -81624 -81203 -81568 -81159
rect -81524 -81203 -81468 -81159
rect -81424 -81203 -80968 -81159
rect -80924 -81203 -80868 -81159
rect -80824 -81203 -80768 -81159
rect -80724 -81203 -80668 -81159
rect -80624 -81203 -80568 -81159
rect -80524 -81203 -80468 -81159
rect -80424 -81203 -80368 -81159
rect -80324 -81203 -80268 -81159
rect -80224 -81203 -80168 -81159
rect -80124 -81203 -80068 -81159
rect -80024 -81203 -79968 -81159
rect -79924 -81203 -79868 -81159
rect -79824 -81203 -79768 -81159
rect -79724 -81203 -79668 -81159
rect -79624 -81203 -79568 -81159
rect -79524 -81203 -79468 -81159
rect -79424 -81203 -78968 -81159
rect -78924 -81203 -78868 -81159
rect -78824 -81203 -78768 -81159
rect -78724 -81203 -78668 -81159
rect -78624 -81203 -78568 -81159
rect -78524 -81203 -78468 -81159
rect -78424 -81203 -78368 -81159
rect -78324 -81203 -78268 -81159
rect -78224 -81203 -78168 -81159
rect -78124 -81203 -78068 -81159
rect -78024 -81203 -77968 -81159
rect -77924 -81203 -77868 -81159
rect -77824 -81203 -77768 -81159
rect -77724 -81203 -77668 -81159
rect -77624 -81203 -77568 -81159
rect -77524 -81203 -77468 -81159
rect -77424 -81203 -76968 -81159
rect -76924 -81203 -76868 -81159
rect -76824 -81203 -76768 -81159
rect -76724 -81203 -76668 -81159
rect -76624 -81203 -76568 -81159
rect -76524 -81203 -76468 -81159
rect -76424 -81203 -76368 -81159
rect -76324 -81203 -76268 -81159
rect -76224 -81203 -76168 -81159
rect -76124 -81203 -76068 -81159
rect -76024 -81203 -75968 -81159
rect -75924 -81203 -75868 -81159
rect -75824 -81203 -75768 -81159
rect -75724 -81203 -75668 -81159
rect -75624 -81203 -75568 -81159
rect -75524 -81203 -75468 -81159
rect -75424 -81161 80737 -81159
rect -75424 -81203 -50017 -81161
rect -109116 -81205 -50017 -81203
rect -49973 -81205 -49917 -81161
rect -49873 -81205 -49817 -81161
rect -49773 -81205 -49717 -81161
rect -49673 -81205 -49617 -81161
rect -49573 -81205 -49517 -81161
rect -49473 -81205 -49417 -81161
rect -49373 -81205 -49317 -81161
rect -49273 -81205 -49217 -81161
rect -49173 -81205 -49117 -81161
rect -49073 -81205 -49017 -81161
rect -48973 -81205 -48917 -81161
rect -48873 -81205 -48817 -81161
rect -48773 -81205 -48717 -81161
rect -48673 -81205 -48617 -81161
rect -48573 -81205 -48517 -81161
rect -48473 -81205 -48017 -81161
rect -47973 -81205 -47917 -81161
rect -47873 -81205 -47817 -81161
rect -47773 -81205 -47717 -81161
rect -47673 -81205 -47617 -81161
rect -47573 -81205 -47517 -81161
rect -47473 -81205 -47417 -81161
rect -47373 -81205 -47317 -81161
rect -47273 -81205 -47217 -81161
rect -47173 -81205 -47117 -81161
rect -47073 -81205 -47017 -81161
rect -46973 -81205 -46917 -81161
rect -46873 -81205 -46817 -81161
rect -46773 -81205 -46717 -81161
rect -46673 -81205 -46617 -81161
rect -46573 -81205 -46517 -81161
rect -46473 -81205 -46017 -81161
rect -45973 -81205 -45917 -81161
rect -45873 -81205 -45817 -81161
rect -45773 -81205 -45717 -81161
rect -45673 -81205 -45617 -81161
rect -45573 -81205 -45517 -81161
rect -45473 -81205 -45417 -81161
rect -45373 -81205 -45317 -81161
rect -45273 -81205 -45217 -81161
rect -45173 -81205 -45117 -81161
rect -45073 -81205 -45017 -81161
rect -44973 -81205 -44917 -81161
rect -44873 -81205 -44817 -81161
rect -44773 -81205 -44717 -81161
rect -44673 -81205 -44617 -81161
rect -44573 -81205 -44517 -81161
rect -44473 -81205 -44017 -81161
rect -43973 -81205 -43917 -81161
rect -43873 -81205 -43817 -81161
rect -43773 -81205 -43717 -81161
rect -43673 -81205 -43617 -81161
rect -43573 -81205 -43517 -81161
rect -43473 -81205 -43417 -81161
rect -43373 -81205 -43317 -81161
rect -43273 -81205 -43217 -81161
rect -43173 -81205 -43117 -81161
rect -43073 -81205 -43017 -81161
rect -42973 -81205 -42917 -81161
rect -42873 -81205 -42817 -81161
rect -42773 -81205 -42717 -81161
rect -42673 -81205 -42617 -81161
rect -42573 -81205 -42517 -81161
rect -42473 -81199 80737 -81161
rect 80781 -81199 80837 -81155
rect 80881 -81199 80937 -81155
rect 80981 -81199 81037 -81155
rect 81081 -81199 81137 -81155
rect 81181 -81199 81237 -81155
rect 81281 -81199 81337 -81155
rect 81381 -81199 81437 -81155
rect 81481 -81199 81537 -81155
rect 81581 -81199 81637 -81155
rect 81681 -81199 81737 -81155
rect 81781 -81199 81837 -81155
rect 81881 -81199 81937 -81155
rect 81981 -81199 82037 -81155
rect 82081 -81199 82137 -81155
rect 82181 -81199 82237 -81155
rect 82281 -81199 82737 -81155
rect 82781 -81199 82837 -81155
rect 82881 -81199 82937 -81155
rect 82981 -81199 83037 -81155
rect 83081 -81199 83137 -81155
rect 83181 -81199 83237 -81155
rect 83281 -81199 83337 -81155
rect 83381 -81199 83437 -81155
rect 83481 -81199 83537 -81155
rect 83581 -81199 83637 -81155
rect 83681 -81199 83737 -81155
rect 83781 -81199 83837 -81155
rect 83881 -81199 83937 -81155
rect 83981 -81199 84037 -81155
rect 84081 -81199 84137 -81155
rect 84181 -81199 84237 -81155
rect 84281 -81199 84737 -81155
rect 84781 -81199 84837 -81155
rect 84881 -81199 84937 -81155
rect 84981 -81199 85037 -81155
rect 85081 -81199 85137 -81155
rect 85181 -81199 85237 -81155
rect 85281 -81199 85337 -81155
rect 85381 -81199 85437 -81155
rect 85481 -81199 85537 -81155
rect 85581 -81199 85637 -81155
rect 85681 -81199 85737 -81155
rect 85781 -81199 85837 -81155
rect 85881 -81199 85937 -81155
rect 85981 -81199 86037 -81155
rect 86081 -81199 86137 -81155
rect 86181 -81199 86237 -81155
rect 86281 -81199 86737 -81155
rect 86781 -81199 86837 -81155
rect 86881 -81199 86937 -81155
rect 86981 -81199 87037 -81155
rect 87081 -81199 87137 -81155
rect 87181 -81199 87237 -81155
rect 87281 -81199 87337 -81155
rect 87381 -81199 87437 -81155
rect 87481 -81199 87537 -81155
rect 87581 -81199 87637 -81155
rect 87681 -81199 87737 -81155
rect 87781 -81199 87837 -81155
rect 87881 -81199 87937 -81155
rect 87981 -81199 88037 -81155
rect 88081 -81199 88137 -81155
rect 88181 -81199 88237 -81155
rect 88281 -81199 177360 -81155
rect -42473 -81205 177360 -81199
rect -109116 -81255 177360 -81205
rect -109116 -81259 80737 -81255
rect -109116 -81303 -82968 -81259
rect -82924 -81303 -82868 -81259
rect -82824 -81303 -82768 -81259
rect -82724 -81303 -82668 -81259
rect -82624 -81303 -82568 -81259
rect -82524 -81303 -82468 -81259
rect -82424 -81303 -82368 -81259
rect -82324 -81303 -82268 -81259
rect -82224 -81303 -82168 -81259
rect -82124 -81303 -82068 -81259
rect -82024 -81303 -81968 -81259
rect -81924 -81303 -81868 -81259
rect -81824 -81303 -81768 -81259
rect -81724 -81303 -81668 -81259
rect -81624 -81303 -81568 -81259
rect -81524 -81303 -81468 -81259
rect -81424 -81303 -80968 -81259
rect -80924 -81303 -80868 -81259
rect -80824 -81303 -80768 -81259
rect -80724 -81303 -80668 -81259
rect -80624 -81303 -80568 -81259
rect -80524 -81303 -80468 -81259
rect -80424 -81303 -80368 -81259
rect -80324 -81303 -80268 -81259
rect -80224 -81303 -80168 -81259
rect -80124 -81303 -80068 -81259
rect -80024 -81303 -79968 -81259
rect -79924 -81303 -79868 -81259
rect -79824 -81303 -79768 -81259
rect -79724 -81303 -79668 -81259
rect -79624 -81303 -79568 -81259
rect -79524 -81303 -79468 -81259
rect -79424 -81303 -78968 -81259
rect -78924 -81303 -78868 -81259
rect -78824 -81303 -78768 -81259
rect -78724 -81303 -78668 -81259
rect -78624 -81303 -78568 -81259
rect -78524 -81303 -78468 -81259
rect -78424 -81303 -78368 -81259
rect -78324 -81303 -78268 -81259
rect -78224 -81303 -78168 -81259
rect -78124 -81303 -78068 -81259
rect -78024 -81303 -77968 -81259
rect -77924 -81303 -77868 -81259
rect -77824 -81303 -77768 -81259
rect -77724 -81303 -77668 -81259
rect -77624 -81303 -77568 -81259
rect -77524 -81303 -77468 -81259
rect -77424 -81303 -76968 -81259
rect -76924 -81303 -76868 -81259
rect -76824 -81303 -76768 -81259
rect -76724 -81303 -76668 -81259
rect -76624 -81303 -76568 -81259
rect -76524 -81303 -76468 -81259
rect -76424 -81303 -76368 -81259
rect -76324 -81303 -76268 -81259
rect -76224 -81303 -76168 -81259
rect -76124 -81303 -76068 -81259
rect -76024 -81303 -75968 -81259
rect -75924 -81303 -75868 -81259
rect -75824 -81303 -75768 -81259
rect -75724 -81303 -75668 -81259
rect -75624 -81303 -75568 -81259
rect -75524 -81303 -75468 -81259
rect -75424 -81261 80737 -81259
rect -75424 -81303 -50017 -81261
rect -109116 -81305 -50017 -81303
rect -49973 -81305 -49917 -81261
rect -49873 -81305 -49817 -81261
rect -49773 -81305 -49717 -81261
rect -49673 -81305 -49617 -81261
rect -49573 -81305 -49517 -81261
rect -49473 -81305 -49417 -81261
rect -49373 -81305 -49317 -81261
rect -49273 -81305 -49217 -81261
rect -49173 -81305 -49117 -81261
rect -49073 -81305 -49017 -81261
rect -48973 -81305 -48917 -81261
rect -48873 -81305 -48817 -81261
rect -48773 -81305 -48717 -81261
rect -48673 -81305 -48617 -81261
rect -48573 -81305 -48517 -81261
rect -48473 -81305 -48017 -81261
rect -47973 -81305 -47917 -81261
rect -47873 -81305 -47817 -81261
rect -47773 -81305 -47717 -81261
rect -47673 -81305 -47617 -81261
rect -47573 -81305 -47517 -81261
rect -47473 -81305 -47417 -81261
rect -47373 -81305 -47317 -81261
rect -47273 -81305 -47217 -81261
rect -47173 -81305 -47117 -81261
rect -47073 -81305 -47017 -81261
rect -46973 -81305 -46917 -81261
rect -46873 -81305 -46817 -81261
rect -46773 -81305 -46717 -81261
rect -46673 -81305 -46617 -81261
rect -46573 -81305 -46517 -81261
rect -46473 -81305 -46017 -81261
rect -45973 -81305 -45917 -81261
rect -45873 -81305 -45817 -81261
rect -45773 -81305 -45717 -81261
rect -45673 -81305 -45617 -81261
rect -45573 -81305 -45517 -81261
rect -45473 -81305 -45417 -81261
rect -45373 -81305 -45317 -81261
rect -45273 -81305 -45217 -81261
rect -45173 -81305 -45117 -81261
rect -45073 -81305 -45017 -81261
rect -44973 -81305 -44917 -81261
rect -44873 -81305 -44817 -81261
rect -44773 -81305 -44717 -81261
rect -44673 -81305 -44617 -81261
rect -44573 -81305 -44517 -81261
rect -44473 -81305 -44017 -81261
rect -43973 -81305 -43917 -81261
rect -43873 -81305 -43817 -81261
rect -43773 -81305 -43717 -81261
rect -43673 -81305 -43617 -81261
rect -43573 -81305 -43517 -81261
rect -43473 -81305 -43417 -81261
rect -43373 -81305 -43317 -81261
rect -43273 -81305 -43217 -81261
rect -43173 -81305 -43117 -81261
rect -43073 -81305 -43017 -81261
rect -42973 -81305 -42917 -81261
rect -42873 -81305 -42817 -81261
rect -42773 -81305 -42717 -81261
rect -42673 -81305 -42617 -81261
rect -42573 -81305 -42517 -81261
rect -42473 -81299 80737 -81261
rect 80781 -81299 80837 -81255
rect 80881 -81299 80937 -81255
rect 80981 -81299 81037 -81255
rect 81081 -81299 81137 -81255
rect 81181 -81299 81237 -81255
rect 81281 -81299 81337 -81255
rect 81381 -81299 81437 -81255
rect 81481 -81299 81537 -81255
rect 81581 -81299 81637 -81255
rect 81681 -81299 81737 -81255
rect 81781 -81299 81837 -81255
rect 81881 -81299 81937 -81255
rect 81981 -81299 82037 -81255
rect 82081 -81299 82137 -81255
rect 82181 -81299 82237 -81255
rect 82281 -81299 82737 -81255
rect 82781 -81299 82837 -81255
rect 82881 -81299 82937 -81255
rect 82981 -81299 83037 -81255
rect 83081 -81299 83137 -81255
rect 83181 -81299 83237 -81255
rect 83281 -81299 83337 -81255
rect 83381 -81299 83437 -81255
rect 83481 -81299 83537 -81255
rect 83581 -81299 83637 -81255
rect 83681 -81299 83737 -81255
rect 83781 -81299 83837 -81255
rect 83881 -81299 83937 -81255
rect 83981 -81299 84037 -81255
rect 84081 -81299 84137 -81255
rect 84181 -81299 84237 -81255
rect 84281 -81299 84737 -81255
rect 84781 -81299 84837 -81255
rect 84881 -81299 84937 -81255
rect 84981 -81299 85037 -81255
rect 85081 -81299 85137 -81255
rect 85181 -81299 85237 -81255
rect 85281 -81299 85337 -81255
rect 85381 -81299 85437 -81255
rect 85481 -81299 85537 -81255
rect 85581 -81299 85637 -81255
rect 85681 -81299 85737 -81255
rect 85781 -81299 85837 -81255
rect 85881 -81299 85937 -81255
rect 85981 -81299 86037 -81255
rect 86081 -81299 86137 -81255
rect 86181 -81299 86237 -81255
rect 86281 -81299 86737 -81255
rect 86781 -81299 86837 -81255
rect 86881 -81299 86937 -81255
rect 86981 -81299 87037 -81255
rect 87081 -81299 87137 -81255
rect 87181 -81299 87237 -81255
rect 87281 -81299 87337 -81255
rect 87381 -81299 87437 -81255
rect 87481 -81299 87537 -81255
rect 87581 -81299 87637 -81255
rect 87681 -81299 87737 -81255
rect 87781 -81299 87837 -81255
rect 87881 -81299 87937 -81255
rect 87981 -81299 88037 -81255
rect 88081 -81299 88137 -81255
rect 88181 -81299 88237 -81255
rect 88281 -81299 177360 -81255
rect -42473 -81305 177360 -81299
rect -109116 -81355 177360 -81305
rect -109116 -81359 80737 -81355
rect -109116 -81403 -82968 -81359
rect -82924 -81403 -82868 -81359
rect -82824 -81403 -82768 -81359
rect -82724 -81403 -82668 -81359
rect -82624 -81403 -82568 -81359
rect -82524 -81403 -82468 -81359
rect -82424 -81403 -82368 -81359
rect -82324 -81403 -82268 -81359
rect -82224 -81403 -82168 -81359
rect -82124 -81403 -82068 -81359
rect -82024 -81403 -81968 -81359
rect -81924 -81403 -81868 -81359
rect -81824 -81403 -81768 -81359
rect -81724 -81403 -81668 -81359
rect -81624 -81403 -81568 -81359
rect -81524 -81403 -81468 -81359
rect -81424 -81403 -80968 -81359
rect -80924 -81403 -80868 -81359
rect -80824 -81403 -80768 -81359
rect -80724 -81403 -80668 -81359
rect -80624 -81403 -80568 -81359
rect -80524 -81403 -80468 -81359
rect -80424 -81403 -80368 -81359
rect -80324 -81403 -80268 -81359
rect -80224 -81403 -80168 -81359
rect -80124 -81403 -80068 -81359
rect -80024 -81403 -79968 -81359
rect -79924 -81403 -79868 -81359
rect -79824 -81403 -79768 -81359
rect -79724 -81403 -79668 -81359
rect -79624 -81403 -79568 -81359
rect -79524 -81403 -79468 -81359
rect -79424 -81403 -78968 -81359
rect -78924 -81403 -78868 -81359
rect -78824 -81403 -78768 -81359
rect -78724 -81403 -78668 -81359
rect -78624 -81403 -78568 -81359
rect -78524 -81403 -78468 -81359
rect -78424 -81403 -78368 -81359
rect -78324 -81403 -78268 -81359
rect -78224 -81403 -78168 -81359
rect -78124 -81403 -78068 -81359
rect -78024 -81403 -77968 -81359
rect -77924 -81403 -77868 -81359
rect -77824 -81403 -77768 -81359
rect -77724 -81403 -77668 -81359
rect -77624 -81403 -77568 -81359
rect -77524 -81403 -77468 -81359
rect -77424 -81403 -76968 -81359
rect -76924 -81403 -76868 -81359
rect -76824 -81403 -76768 -81359
rect -76724 -81403 -76668 -81359
rect -76624 -81403 -76568 -81359
rect -76524 -81403 -76468 -81359
rect -76424 -81403 -76368 -81359
rect -76324 -81403 -76268 -81359
rect -76224 -81403 -76168 -81359
rect -76124 -81403 -76068 -81359
rect -76024 -81403 -75968 -81359
rect -75924 -81403 -75868 -81359
rect -75824 -81403 -75768 -81359
rect -75724 -81403 -75668 -81359
rect -75624 -81403 -75568 -81359
rect -75524 -81403 -75468 -81359
rect -75424 -81361 80737 -81359
rect -75424 -81403 -50017 -81361
rect -109116 -81405 -50017 -81403
rect -49973 -81405 -49917 -81361
rect -49873 -81405 -49817 -81361
rect -49773 -81405 -49717 -81361
rect -49673 -81405 -49617 -81361
rect -49573 -81405 -49517 -81361
rect -49473 -81405 -49417 -81361
rect -49373 -81405 -49317 -81361
rect -49273 -81405 -49217 -81361
rect -49173 -81405 -49117 -81361
rect -49073 -81405 -49017 -81361
rect -48973 -81405 -48917 -81361
rect -48873 -81405 -48817 -81361
rect -48773 -81405 -48717 -81361
rect -48673 -81405 -48617 -81361
rect -48573 -81405 -48517 -81361
rect -48473 -81405 -48017 -81361
rect -47973 -81405 -47917 -81361
rect -47873 -81405 -47817 -81361
rect -47773 -81405 -47717 -81361
rect -47673 -81405 -47617 -81361
rect -47573 -81405 -47517 -81361
rect -47473 -81405 -47417 -81361
rect -47373 -81405 -47317 -81361
rect -47273 -81405 -47217 -81361
rect -47173 -81405 -47117 -81361
rect -47073 -81405 -47017 -81361
rect -46973 -81405 -46917 -81361
rect -46873 -81405 -46817 -81361
rect -46773 -81405 -46717 -81361
rect -46673 -81405 -46617 -81361
rect -46573 -81405 -46517 -81361
rect -46473 -81405 -46017 -81361
rect -45973 -81405 -45917 -81361
rect -45873 -81405 -45817 -81361
rect -45773 -81405 -45717 -81361
rect -45673 -81405 -45617 -81361
rect -45573 -81405 -45517 -81361
rect -45473 -81405 -45417 -81361
rect -45373 -81405 -45317 -81361
rect -45273 -81405 -45217 -81361
rect -45173 -81405 -45117 -81361
rect -45073 -81405 -45017 -81361
rect -44973 -81405 -44917 -81361
rect -44873 -81405 -44817 -81361
rect -44773 -81405 -44717 -81361
rect -44673 -81405 -44617 -81361
rect -44573 -81405 -44517 -81361
rect -44473 -81405 -44017 -81361
rect -43973 -81405 -43917 -81361
rect -43873 -81405 -43817 -81361
rect -43773 -81405 -43717 -81361
rect -43673 -81405 -43617 -81361
rect -43573 -81405 -43517 -81361
rect -43473 -81405 -43417 -81361
rect -43373 -81405 -43317 -81361
rect -43273 -81405 -43217 -81361
rect -43173 -81405 -43117 -81361
rect -43073 -81405 -43017 -81361
rect -42973 -81405 -42917 -81361
rect -42873 -81405 -42817 -81361
rect -42773 -81405 -42717 -81361
rect -42673 -81405 -42617 -81361
rect -42573 -81405 -42517 -81361
rect -42473 -81399 80737 -81361
rect 80781 -81399 80837 -81355
rect 80881 -81399 80937 -81355
rect 80981 -81399 81037 -81355
rect 81081 -81399 81137 -81355
rect 81181 -81399 81237 -81355
rect 81281 -81399 81337 -81355
rect 81381 -81399 81437 -81355
rect 81481 -81399 81537 -81355
rect 81581 -81399 81637 -81355
rect 81681 -81399 81737 -81355
rect 81781 -81399 81837 -81355
rect 81881 -81399 81937 -81355
rect 81981 -81399 82037 -81355
rect 82081 -81399 82137 -81355
rect 82181 -81399 82237 -81355
rect 82281 -81399 82737 -81355
rect 82781 -81399 82837 -81355
rect 82881 -81399 82937 -81355
rect 82981 -81399 83037 -81355
rect 83081 -81399 83137 -81355
rect 83181 -81399 83237 -81355
rect 83281 -81399 83337 -81355
rect 83381 -81399 83437 -81355
rect 83481 -81399 83537 -81355
rect 83581 -81399 83637 -81355
rect 83681 -81399 83737 -81355
rect 83781 -81399 83837 -81355
rect 83881 -81399 83937 -81355
rect 83981 -81399 84037 -81355
rect 84081 -81399 84137 -81355
rect 84181 -81399 84237 -81355
rect 84281 -81399 84737 -81355
rect 84781 -81399 84837 -81355
rect 84881 -81399 84937 -81355
rect 84981 -81399 85037 -81355
rect 85081 -81399 85137 -81355
rect 85181 -81399 85237 -81355
rect 85281 -81399 85337 -81355
rect 85381 -81399 85437 -81355
rect 85481 -81399 85537 -81355
rect 85581 -81399 85637 -81355
rect 85681 -81399 85737 -81355
rect 85781 -81399 85837 -81355
rect 85881 -81399 85937 -81355
rect 85981 -81399 86037 -81355
rect 86081 -81399 86137 -81355
rect 86181 -81399 86237 -81355
rect 86281 -81399 86737 -81355
rect 86781 -81399 86837 -81355
rect 86881 -81399 86937 -81355
rect 86981 -81399 87037 -81355
rect 87081 -81399 87137 -81355
rect 87181 -81399 87237 -81355
rect 87281 -81399 87337 -81355
rect 87381 -81399 87437 -81355
rect 87481 -81399 87537 -81355
rect 87581 -81399 87637 -81355
rect 87681 -81399 87737 -81355
rect 87781 -81399 87837 -81355
rect 87881 -81399 87937 -81355
rect 87981 -81399 88037 -81355
rect 88081 -81399 88137 -81355
rect 88181 -81399 88237 -81355
rect 88281 -81399 177360 -81355
rect -42473 -81405 177360 -81399
rect -109116 -81455 177360 -81405
rect -109116 -81459 80737 -81455
rect -109116 -81503 -82968 -81459
rect -82924 -81503 -82868 -81459
rect -82824 -81503 -82768 -81459
rect -82724 -81503 -82668 -81459
rect -82624 -81503 -82568 -81459
rect -82524 -81503 -82468 -81459
rect -82424 -81503 -82368 -81459
rect -82324 -81503 -82268 -81459
rect -82224 -81503 -82168 -81459
rect -82124 -81503 -82068 -81459
rect -82024 -81503 -81968 -81459
rect -81924 -81503 -81868 -81459
rect -81824 -81503 -81768 -81459
rect -81724 -81503 -81668 -81459
rect -81624 -81503 -81568 -81459
rect -81524 -81503 -81468 -81459
rect -81424 -81503 -80968 -81459
rect -80924 -81503 -80868 -81459
rect -80824 -81503 -80768 -81459
rect -80724 -81503 -80668 -81459
rect -80624 -81503 -80568 -81459
rect -80524 -81503 -80468 -81459
rect -80424 -81503 -80368 -81459
rect -80324 -81503 -80268 -81459
rect -80224 -81503 -80168 -81459
rect -80124 -81503 -80068 -81459
rect -80024 -81503 -79968 -81459
rect -79924 -81503 -79868 -81459
rect -79824 -81503 -79768 -81459
rect -79724 -81503 -79668 -81459
rect -79624 -81503 -79568 -81459
rect -79524 -81503 -79468 -81459
rect -79424 -81503 -78968 -81459
rect -78924 -81503 -78868 -81459
rect -78824 -81503 -78768 -81459
rect -78724 -81503 -78668 -81459
rect -78624 -81503 -78568 -81459
rect -78524 -81503 -78468 -81459
rect -78424 -81503 -78368 -81459
rect -78324 -81503 -78268 -81459
rect -78224 -81503 -78168 -81459
rect -78124 -81503 -78068 -81459
rect -78024 -81503 -77968 -81459
rect -77924 -81503 -77868 -81459
rect -77824 -81503 -77768 -81459
rect -77724 -81503 -77668 -81459
rect -77624 -81503 -77568 -81459
rect -77524 -81503 -77468 -81459
rect -77424 -81503 -76968 -81459
rect -76924 -81503 -76868 -81459
rect -76824 -81503 -76768 -81459
rect -76724 -81503 -76668 -81459
rect -76624 -81503 -76568 -81459
rect -76524 -81503 -76468 -81459
rect -76424 -81503 -76368 -81459
rect -76324 -81503 -76268 -81459
rect -76224 -81503 -76168 -81459
rect -76124 -81503 -76068 -81459
rect -76024 -81503 -75968 -81459
rect -75924 -81503 -75868 -81459
rect -75824 -81503 -75768 -81459
rect -75724 -81503 -75668 -81459
rect -75624 -81503 -75568 -81459
rect -75524 -81503 -75468 -81459
rect -75424 -81461 80737 -81459
rect -75424 -81503 -50017 -81461
rect -109116 -81505 -50017 -81503
rect -49973 -81505 -49917 -81461
rect -49873 -81505 -49817 -81461
rect -49773 -81505 -49717 -81461
rect -49673 -81505 -49617 -81461
rect -49573 -81505 -49517 -81461
rect -49473 -81505 -49417 -81461
rect -49373 -81505 -49317 -81461
rect -49273 -81505 -49217 -81461
rect -49173 -81505 -49117 -81461
rect -49073 -81505 -49017 -81461
rect -48973 -81505 -48917 -81461
rect -48873 -81505 -48817 -81461
rect -48773 -81505 -48717 -81461
rect -48673 -81505 -48617 -81461
rect -48573 -81505 -48517 -81461
rect -48473 -81505 -48017 -81461
rect -47973 -81505 -47917 -81461
rect -47873 -81505 -47817 -81461
rect -47773 -81505 -47717 -81461
rect -47673 -81505 -47617 -81461
rect -47573 -81505 -47517 -81461
rect -47473 -81505 -47417 -81461
rect -47373 -81505 -47317 -81461
rect -47273 -81505 -47217 -81461
rect -47173 -81505 -47117 -81461
rect -47073 -81505 -47017 -81461
rect -46973 -81505 -46917 -81461
rect -46873 -81505 -46817 -81461
rect -46773 -81505 -46717 -81461
rect -46673 -81505 -46617 -81461
rect -46573 -81505 -46517 -81461
rect -46473 -81505 -46017 -81461
rect -45973 -81505 -45917 -81461
rect -45873 -81505 -45817 -81461
rect -45773 -81505 -45717 -81461
rect -45673 -81505 -45617 -81461
rect -45573 -81505 -45517 -81461
rect -45473 -81505 -45417 -81461
rect -45373 -81505 -45317 -81461
rect -45273 -81505 -45217 -81461
rect -45173 -81505 -45117 -81461
rect -45073 -81505 -45017 -81461
rect -44973 -81505 -44917 -81461
rect -44873 -81505 -44817 -81461
rect -44773 -81505 -44717 -81461
rect -44673 -81505 -44617 -81461
rect -44573 -81505 -44517 -81461
rect -44473 -81505 -44017 -81461
rect -43973 -81505 -43917 -81461
rect -43873 -81505 -43817 -81461
rect -43773 -81505 -43717 -81461
rect -43673 -81505 -43617 -81461
rect -43573 -81505 -43517 -81461
rect -43473 -81505 -43417 -81461
rect -43373 -81505 -43317 -81461
rect -43273 -81505 -43217 -81461
rect -43173 -81505 -43117 -81461
rect -43073 -81505 -43017 -81461
rect -42973 -81505 -42917 -81461
rect -42873 -81505 -42817 -81461
rect -42773 -81505 -42717 -81461
rect -42673 -81505 -42617 -81461
rect -42573 -81505 -42517 -81461
rect -42473 -81499 80737 -81461
rect 80781 -81499 80837 -81455
rect 80881 -81499 80937 -81455
rect 80981 -81499 81037 -81455
rect 81081 -81499 81137 -81455
rect 81181 -81499 81237 -81455
rect 81281 -81499 81337 -81455
rect 81381 -81499 81437 -81455
rect 81481 -81499 81537 -81455
rect 81581 -81499 81637 -81455
rect 81681 -81499 81737 -81455
rect 81781 -81499 81837 -81455
rect 81881 -81499 81937 -81455
rect 81981 -81499 82037 -81455
rect 82081 -81499 82137 -81455
rect 82181 -81499 82237 -81455
rect 82281 -81499 82737 -81455
rect 82781 -81499 82837 -81455
rect 82881 -81499 82937 -81455
rect 82981 -81499 83037 -81455
rect 83081 -81499 83137 -81455
rect 83181 -81499 83237 -81455
rect 83281 -81499 83337 -81455
rect 83381 -81499 83437 -81455
rect 83481 -81499 83537 -81455
rect 83581 -81499 83637 -81455
rect 83681 -81499 83737 -81455
rect 83781 -81499 83837 -81455
rect 83881 -81499 83937 -81455
rect 83981 -81499 84037 -81455
rect 84081 -81499 84137 -81455
rect 84181 -81499 84237 -81455
rect 84281 -81499 84737 -81455
rect 84781 -81499 84837 -81455
rect 84881 -81499 84937 -81455
rect 84981 -81499 85037 -81455
rect 85081 -81499 85137 -81455
rect 85181 -81499 85237 -81455
rect 85281 -81499 85337 -81455
rect 85381 -81499 85437 -81455
rect 85481 -81499 85537 -81455
rect 85581 -81499 85637 -81455
rect 85681 -81499 85737 -81455
rect 85781 -81499 85837 -81455
rect 85881 -81499 85937 -81455
rect 85981 -81499 86037 -81455
rect 86081 -81499 86137 -81455
rect 86181 -81499 86237 -81455
rect 86281 -81499 86737 -81455
rect 86781 -81499 86837 -81455
rect 86881 -81499 86937 -81455
rect 86981 -81499 87037 -81455
rect 87081 -81499 87137 -81455
rect 87181 -81499 87237 -81455
rect 87281 -81499 87337 -81455
rect 87381 -81499 87437 -81455
rect 87481 -81499 87537 -81455
rect 87581 -81499 87637 -81455
rect 87681 -81499 87737 -81455
rect 87781 -81499 87837 -81455
rect 87881 -81499 87937 -81455
rect 87981 -81499 88037 -81455
rect 88081 -81499 88137 -81455
rect 88181 -81499 88237 -81455
rect 88281 -81499 177360 -81455
rect -42473 -81505 177360 -81499
rect -109116 -81555 177360 -81505
rect -109116 -81559 80737 -81555
rect -109116 -81603 -82968 -81559
rect -82924 -81603 -82868 -81559
rect -82824 -81603 -82768 -81559
rect -82724 -81603 -82668 -81559
rect -82624 -81603 -82568 -81559
rect -82524 -81603 -82468 -81559
rect -82424 -81603 -82368 -81559
rect -82324 -81603 -82268 -81559
rect -82224 -81603 -82168 -81559
rect -82124 -81603 -82068 -81559
rect -82024 -81603 -81968 -81559
rect -81924 -81603 -81868 -81559
rect -81824 -81603 -81768 -81559
rect -81724 -81603 -81668 -81559
rect -81624 -81603 -81568 -81559
rect -81524 -81603 -81468 -81559
rect -81424 -81603 -80968 -81559
rect -80924 -81603 -80868 -81559
rect -80824 -81603 -80768 -81559
rect -80724 -81603 -80668 -81559
rect -80624 -81603 -80568 -81559
rect -80524 -81603 -80468 -81559
rect -80424 -81603 -80368 -81559
rect -80324 -81603 -80268 -81559
rect -80224 -81603 -80168 -81559
rect -80124 -81603 -80068 -81559
rect -80024 -81603 -79968 -81559
rect -79924 -81603 -79868 -81559
rect -79824 -81603 -79768 -81559
rect -79724 -81603 -79668 -81559
rect -79624 -81603 -79568 -81559
rect -79524 -81603 -79468 -81559
rect -79424 -81603 -78968 -81559
rect -78924 -81603 -78868 -81559
rect -78824 -81603 -78768 -81559
rect -78724 -81603 -78668 -81559
rect -78624 -81603 -78568 -81559
rect -78524 -81603 -78468 -81559
rect -78424 -81603 -78368 -81559
rect -78324 -81603 -78268 -81559
rect -78224 -81603 -78168 -81559
rect -78124 -81603 -78068 -81559
rect -78024 -81603 -77968 -81559
rect -77924 -81603 -77868 -81559
rect -77824 -81603 -77768 -81559
rect -77724 -81603 -77668 -81559
rect -77624 -81603 -77568 -81559
rect -77524 -81603 -77468 -81559
rect -77424 -81603 -76968 -81559
rect -76924 -81603 -76868 -81559
rect -76824 -81603 -76768 -81559
rect -76724 -81603 -76668 -81559
rect -76624 -81603 -76568 -81559
rect -76524 -81603 -76468 -81559
rect -76424 -81603 -76368 -81559
rect -76324 -81603 -76268 -81559
rect -76224 -81603 -76168 -81559
rect -76124 -81603 -76068 -81559
rect -76024 -81603 -75968 -81559
rect -75924 -81603 -75868 -81559
rect -75824 -81603 -75768 -81559
rect -75724 -81603 -75668 -81559
rect -75624 -81603 -75568 -81559
rect -75524 -81603 -75468 -81559
rect -75424 -81561 80737 -81559
rect -75424 -81603 -50017 -81561
rect -109116 -81605 -50017 -81603
rect -49973 -81605 -49917 -81561
rect -49873 -81605 -49817 -81561
rect -49773 -81605 -49717 -81561
rect -49673 -81605 -49617 -81561
rect -49573 -81605 -49517 -81561
rect -49473 -81605 -49417 -81561
rect -49373 -81605 -49317 -81561
rect -49273 -81605 -49217 -81561
rect -49173 -81605 -49117 -81561
rect -49073 -81605 -49017 -81561
rect -48973 -81605 -48917 -81561
rect -48873 -81605 -48817 -81561
rect -48773 -81605 -48717 -81561
rect -48673 -81605 -48617 -81561
rect -48573 -81605 -48517 -81561
rect -48473 -81605 -48017 -81561
rect -47973 -81605 -47917 -81561
rect -47873 -81605 -47817 -81561
rect -47773 -81605 -47717 -81561
rect -47673 -81605 -47617 -81561
rect -47573 -81605 -47517 -81561
rect -47473 -81605 -47417 -81561
rect -47373 -81605 -47317 -81561
rect -47273 -81605 -47217 -81561
rect -47173 -81605 -47117 -81561
rect -47073 -81605 -47017 -81561
rect -46973 -81605 -46917 -81561
rect -46873 -81605 -46817 -81561
rect -46773 -81605 -46717 -81561
rect -46673 -81605 -46617 -81561
rect -46573 -81605 -46517 -81561
rect -46473 -81605 -46017 -81561
rect -45973 -81605 -45917 -81561
rect -45873 -81605 -45817 -81561
rect -45773 -81605 -45717 -81561
rect -45673 -81605 -45617 -81561
rect -45573 -81605 -45517 -81561
rect -45473 -81605 -45417 -81561
rect -45373 -81605 -45317 -81561
rect -45273 -81605 -45217 -81561
rect -45173 -81605 -45117 -81561
rect -45073 -81605 -45017 -81561
rect -44973 -81605 -44917 -81561
rect -44873 -81605 -44817 -81561
rect -44773 -81605 -44717 -81561
rect -44673 -81605 -44617 -81561
rect -44573 -81605 -44517 -81561
rect -44473 -81605 -44017 -81561
rect -43973 -81605 -43917 -81561
rect -43873 -81605 -43817 -81561
rect -43773 -81605 -43717 -81561
rect -43673 -81605 -43617 -81561
rect -43573 -81605 -43517 -81561
rect -43473 -81605 -43417 -81561
rect -43373 -81605 -43317 -81561
rect -43273 -81605 -43217 -81561
rect -43173 -81605 -43117 -81561
rect -43073 -81605 -43017 -81561
rect -42973 -81605 -42917 -81561
rect -42873 -81605 -42817 -81561
rect -42773 -81605 -42717 -81561
rect -42673 -81605 -42617 -81561
rect -42573 -81605 -42517 -81561
rect -42473 -81599 80737 -81561
rect 80781 -81599 80837 -81555
rect 80881 -81599 80937 -81555
rect 80981 -81599 81037 -81555
rect 81081 -81599 81137 -81555
rect 81181 -81599 81237 -81555
rect 81281 -81599 81337 -81555
rect 81381 -81599 81437 -81555
rect 81481 -81599 81537 -81555
rect 81581 -81599 81637 -81555
rect 81681 -81599 81737 -81555
rect 81781 -81599 81837 -81555
rect 81881 -81599 81937 -81555
rect 81981 -81599 82037 -81555
rect 82081 -81599 82137 -81555
rect 82181 -81599 82237 -81555
rect 82281 -81599 82737 -81555
rect 82781 -81599 82837 -81555
rect 82881 -81599 82937 -81555
rect 82981 -81599 83037 -81555
rect 83081 -81599 83137 -81555
rect 83181 -81599 83237 -81555
rect 83281 -81599 83337 -81555
rect 83381 -81599 83437 -81555
rect 83481 -81599 83537 -81555
rect 83581 -81599 83637 -81555
rect 83681 -81599 83737 -81555
rect 83781 -81599 83837 -81555
rect 83881 -81599 83937 -81555
rect 83981 -81599 84037 -81555
rect 84081 -81599 84137 -81555
rect 84181 -81599 84237 -81555
rect 84281 -81599 84737 -81555
rect 84781 -81599 84837 -81555
rect 84881 -81599 84937 -81555
rect 84981 -81599 85037 -81555
rect 85081 -81599 85137 -81555
rect 85181 -81599 85237 -81555
rect 85281 -81599 85337 -81555
rect 85381 -81599 85437 -81555
rect 85481 -81599 85537 -81555
rect 85581 -81599 85637 -81555
rect 85681 -81599 85737 -81555
rect 85781 -81599 85837 -81555
rect 85881 -81599 85937 -81555
rect 85981 -81599 86037 -81555
rect 86081 -81599 86137 -81555
rect 86181 -81599 86237 -81555
rect 86281 -81599 86737 -81555
rect 86781 -81599 86837 -81555
rect 86881 -81599 86937 -81555
rect 86981 -81599 87037 -81555
rect 87081 -81599 87137 -81555
rect 87181 -81599 87237 -81555
rect 87281 -81599 87337 -81555
rect 87381 -81599 87437 -81555
rect 87481 -81599 87537 -81555
rect 87581 -81599 87637 -81555
rect 87681 -81599 87737 -81555
rect 87781 -81599 87837 -81555
rect 87881 -81599 87937 -81555
rect 87981 -81599 88037 -81555
rect 88081 -81599 88137 -81555
rect 88181 -81599 88237 -81555
rect 88281 -81599 177360 -81555
rect -42473 -81605 177360 -81599
rect -109116 -81655 177360 -81605
rect -109116 -81659 80737 -81655
rect -109116 -81703 -82968 -81659
rect -82924 -81703 -82868 -81659
rect -82824 -81703 -82768 -81659
rect -82724 -81703 -82668 -81659
rect -82624 -81703 -82568 -81659
rect -82524 -81703 -82468 -81659
rect -82424 -81703 -82368 -81659
rect -82324 -81703 -82268 -81659
rect -82224 -81703 -82168 -81659
rect -82124 -81703 -82068 -81659
rect -82024 -81703 -81968 -81659
rect -81924 -81703 -81868 -81659
rect -81824 -81703 -81768 -81659
rect -81724 -81703 -81668 -81659
rect -81624 -81703 -81568 -81659
rect -81524 -81703 -81468 -81659
rect -81424 -81703 -80968 -81659
rect -80924 -81703 -80868 -81659
rect -80824 -81703 -80768 -81659
rect -80724 -81703 -80668 -81659
rect -80624 -81703 -80568 -81659
rect -80524 -81703 -80468 -81659
rect -80424 -81703 -80368 -81659
rect -80324 -81703 -80268 -81659
rect -80224 -81703 -80168 -81659
rect -80124 -81703 -80068 -81659
rect -80024 -81703 -79968 -81659
rect -79924 -81703 -79868 -81659
rect -79824 -81703 -79768 -81659
rect -79724 -81703 -79668 -81659
rect -79624 -81703 -79568 -81659
rect -79524 -81703 -79468 -81659
rect -79424 -81703 -78968 -81659
rect -78924 -81703 -78868 -81659
rect -78824 -81703 -78768 -81659
rect -78724 -81703 -78668 -81659
rect -78624 -81703 -78568 -81659
rect -78524 -81703 -78468 -81659
rect -78424 -81703 -78368 -81659
rect -78324 -81703 -78268 -81659
rect -78224 -81703 -78168 -81659
rect -78124 -81703 -78068 -81659
rect -78024 -81703 -77968 -81659
rect -77924 -81703 -77868 -81659
rect -77824 -81703 -77768 -81659
rect -77724 -81703 -77668 -81659
rect -77624 -81703 -77568 -81659
rect -77524 -81703 -77468 -81659
rect -77424 -81703 -76968 -81659
rect -76924 -81703 -76868 -81659
rect -76824 -81703 -76768 -81659
rect -76724 -81703 -76668 -81659
rect -76624 -81703 -76568 -81659
rect -76524 -81703 -76468 -81659
rect -76424 -81703 -76368 -81659
rect -76324 -81703 -76268 -81659
rect -76224 -81703 -76168 -81659
rect -76124 -81703 -76068 -81659
rect -76024 -81703 -75968 -81659
rect -75924 -81703 -75868 -81659
rect -75824 -81703 -75768 -81659
rect -75724 -81703 -75668 -81659
rect -75624 -81703 -75568 -81659
rect -75524 -81703 -75468 -81659
rect -75424 -81661 80737 -81659
rect -75424 -81703 -50017 -81661
rect -109116 -81705 -50017 -81703
rect -49973 -81705 -49917 -81661
rect -49873 -81705 -49817 -81661
rect -49773 -81705 -49717 -81661
rect -49673 -81705 -49617 -81661
rect -49573 -81705 -49517 -81661
rect -49473 -81705 -49417 -81661
rect -49373 -81705 -49317 -81661
rect -49273 -81705 -49217 -81661
rect -49173 -81705 -49117 -81661
rect -49073 -81705 -49017 -81661
rect -48973 -81705 -48917 -81661
rect -48873 -81705 -48817 -81661
rect -48773 -81705 -48717 -81661
rect -48673 -81705 -48617 -81661
rect -48573 -81705 -48517 -81661
rect -48473 -81705 -48017 -81661
rect -47973 -81705 -47917 -81661
rect -47873 -81705 -47817 -81661
rect -47773 -81705 -47717 -81661
rect -47673 -81705 -47617 -81661
rect -47573 -81705 -47517 -81661
rect -47473 -81705 -47417 -81661
rect -47373 -81705 -47317 -81661
rect -47273 -81705 -47217 -81661
rect -47173 -81705 -47117 -81661
rect -47073 -81705 -47017 -81661
rect -46973 -81705 -46917 -81661
rect -46873 -81705 -46817 -81661
rect -46773 -81705 -46717 -81661
rect -46673 -81705 -46617 -81661
rect -46573 -81705 -46517 -81661
rect -46473 -81705 -46017 -81661
rect -45973 -81705 -45917 -81661
rect -45873 -81705 -45817 -81661
rect -45773 -81705 -45717 -81661
rect -45673 -81705 -45617 -81661
rect -45573 -81705 -45517 -81661
rect -45473 -81705 -45417 -81661
rect -45373 -81705 -45317 -81661
rect -45273 -81705 -45217 -81661
rect -45173 -81705 -45117 -81661
rect -45073 -81705 -45017 -81661
rect -44973 -81705 -44917 -81661
rect -44873 -81705 -44817 -81661
rect -44773 -81705 -44717 -81661
rect -44673 -81705 -44617 -81661
rect -44573 -81705 -44517 -81661
rect -44473 -81705 -44017 -81661
rect -43973 -81705 -43917 -81661
rect -43873 -81705 -43817 -81661
rect -43773 -81705 -43717 -81661
rect -43673 -81705 -43617 -81661
rect -43573 -81705 -43517 -81661
rect -43473 -81705 -43417 -81661
rect -43373 -81705 -43317 -81661
rect -43273 -81705 -43217 -81661
rect -43173 -81705 -43117 -81661
rect -43073 -81705 -43017 -81661
rect -42973 -81705 -42917 -81661
rect -42873 -81705 -42817 -81661
rect -42773 -81705 -42717 -81661
rect -42673 -81705 -42617 -81661
rect -42573 -81705 -42517 -81661
rect -42473 -81699 80737 -81661
rect 80781 -81699 80837 -81655
rect 80881 -81699 80937 -81655
rect 80981 -81699 81037 -81655
rect 81081 -81699 81137 -81655
rect 81181 -81699 81237 -81655
rect 81281 -81699 81337 -81655
rect 81381 -81699 81437 -81655
rect 81481 -81699 81537 -81655
rect 81581 -81699 81637 -81655
rect 81681 -81699 81737 -81655
rect 81781 -81699 81837 -81655
rect 81881 -81699 81937 -81655
rect 81981 -81699 82037 -81655
rect 82081 -81699 82137 -81655
rect 82181 -81699 82237 -81655
rect 82281 -81699 82737 -81655
rect 82781 -81699 82837 -81655
rect 82881 -81699 82937 -81655
rect 82981 -81699 83037 -81655
rect 83081 -81699 83137 -81655
rect 83181 -81699 83237 -81655
rect 83281 -81699 83337 -81655
rect 83381 -81699 83437 -81655
rect 83481 -81699 83537 -81655
rect 83581 -81699 83637 -81655
rect 83681 -81699 83737 -81655
rect 83781 -81699 83837 -81655
rect 83881 -81699 83937 -81655
rect 83981 -81699 84037 -81655
rect 84081 -81699 84137 -81655
rect 84181 -81699 84237 -81655
rect 84281 -81699 84737 -81655
rect 84781 -81699 84837 -81655
rect 84881 -81699 84937 -81655
rect 84981 -81699 85037 -81655
rect 85081 -81699 85137 -81655
rect 85181 -81699 85237 -81655
rect 85281 -81699 85337 -81655
rect 85381 -81699 85437 -81655
rect 85481 -81699 85537 -81655
rect 85581 -81699 85637 -81655
rect 85681 -81699 85737 -81655
rect 85781 -81699 85837 -81655
rect 85881 -81699 85937 -81655
rect 85981 -81699 86037 -81655
rect 86081 -81699 86137 -81655
rect 86181 -81699 86237 -81655
rect 86281 -81699 86737 -81655
rect 86781 -81699 86837 -81655
rect 86881 -81699 86937 -81655
rect 86981 -81699 87037 -81655
rect 87081 -81699 87137 -81655
rect 87181 -81699 87237 -81655
rect 87281 -81699 87337 -81655
rect 87381 -81699 87437 -81655
rect 87481 -81699 87537 -81655
rect 87581 -81699 87637 -81655
rect 87681 -81699 87737 -81655
rect 87781 -81699 87837 -81655
rect 87881 -81699 87937 -81655
rect 87981 -81699 88037 -81655
rect 88081 -81699 88137 -81655
rect 88181 -81699 88237 -81655
rect 88281 -81699 177360 -81655
rect -42473 -81705 177360 -81699
rect -109116 -81755 177360 -81705
rect -109116 -81759 80737 -81755
rect -109116 -81803 -82968 -81759
rect -82924 -81803 -82868 -81759
rect -82824 -81803 -82768 -81759
rect -82724 -81803 -82668 -81759
rect -82624 -81803 -82568 -81759
rect -82524 -81803 -82468 -81759
rect -82424 -81803 -82368 -81759
rect -82324 -81803 -82268 -81759
rect -82224 -81803 -82168 -81759
rect -82124 -81803 -82068 -81759
rect -82024 -81803 -81968 -81759
rect -81924 -81803 -81868 -81759
rect -81824 -81803 -81768 -81759
rect -81724 -81803 -81668 -81759
rect -81624 -81803 -81568 -81759
rect -81524 -81803 -81468 -81759
rect -81424 -81803 -80968 -81759
rect -80924 -81803 -80868 -81759
rect -80824 -81803 -80768 -81759
rect -80724 -81803 -80668 -81759
rect -80624 -81803 -80568 -81759
rect -80524 -81803 -80468 -81759
rect -80424 -81803 -80368 -81759
rect -80324 -81803 -80268 -81759
rect -80224 -81803 -80168 -81759
rect -80124 -81803 -80068 -81759
rect -80024 -81803 -79968 -81759
rect -79924 -81803 -79868 -81759
rect -79824 -81803 -79768 -81759
rect -79724 -81803 -79668 -81759
rect -79624 -81803 -79568 -81759
rect -79524 -81803 -79468 -81759
rect -79424 -81803 -78968 -81759
rect -78924 -81803 -78868 -81759
rect -78824 -81803 -78768 -81759
rect -78724 -81803 -78668 -81759
rect -78624 -81803 -78568 -81759
rect -78524 -81803 -78468 -81759
rect -78424 -81803 -78368 -81759
rect -78324 -81803 -78268 -81759
rect -78224 -81803 -78168 -81759
rect -78124 -81803 -78068 -81759
rect -78024 -81803 -77968 -81759
rect -77924 -81803 -77868 -81759
rect -77824 -81803 -77768 -81759
rect -77724 -81803 -77668 -81759
rect -77624 -81803 -77568 -81759
rect -77524 -81803 -77468 -81759
rect -77424 -81803 -76968 -81759
rect -76924 -81803 -76868 -81759
rect -76824 -81803 -76768 -81759
rect -76724 -81803 -76668 -81759
rect -76624 -81803 -76568 -81759
rect -76524 -81803 -76468 -81759
rect -76424 -81803 -76368 -81759
rect -76324 -81803 -76268 -81759
rect -76224 -81803 -76168 -81759
rect -76124 -81803 -76068 -81759
rect -76024 -81803 -75968 -81759
rect -75924 -81803 -75868 -81759
rect -75824 -81803 -75768 -81759
rect -75724 -81803 -75668 -81759
rect -75624 -81803 -75568 -81759
rect -75524 -81803 -75468 -81759
rect -75424 -81761 80737 -81759
rect -75424 -81803 -50017 -81761
rect -109116 -81805 -50017 -81803
rect -49973 -81805 -49917 -81761
rect -49873 -81805 -49817 -81761
rect -49773 -81805 -49717 -81761
rect -49673 -81805 -49617 -81761
rect -49573 -81805 -49517 -81761
rect -49473 -81805 -49417 -81761
rect -49373 -81805 -49317 -81761
rect -49273 -81805 -49217 -81761
rect -49173 -81805 -49117 -81761
rect -49073 -81805 -49017 -81761
rect -48973 -81805 -48917 -81761
rect -48873 -81805 -48817 -81761
rect -48773 -81805 -48717 -81761
rect -48673 -81805 -48617 -81761
rect -48573 -81805 -48517 -81761
rect -48473 -81805 -48017 -81761
rect -47973 -81805 -47917 -81761
rect -47873 -81805 -47817 -81761
rect -47773 -81805 -47717 -81761
rect -47673 -81805 -47617 -81761
rect -47573 -81805 -47517 -81761
rect -47473 -81805 -47417 -81761
rect -47373 -81805 -47317 -81761
rect -47273 -81805 -47217 -81761
rect -47173 -81805 -47117 -81761
rect -47073 -81805 -47017 -81761
rect -46973 -81805 -46917 -81761
rect -46873 -81805 -46817 -81761
rect -46773 -81805 -46717 -81761
rect -46673 -81805 -46617 -81761
rect -46573 -81805 -46517 -81761
rect -46473 -81805 -46017 -81761
rect -45973 -81805 -45917 -81761
rect -45873 -81805 -45817 -81761
rect -45773 -81805 -45717 -81761
rect -45673 -81805 -45617 -81761
rect -45573 -81805 -45517 -81761
rect -45473 -81805 -45417 -81761
rect -45373 -81805 -45317 -81761
rect -45273 -81805 -45217 -81761
rect -45173 -81805 -45117 -81761
rect -45073 -81805 -45017 -81761
rect -44973 -81805 -44917 -81761
rect -44873 -81805 -44817 -81761
rect -44773 -81805 -44717 -81761
rect -44673 -81805 -44617 -81761
rect -44573 -81805 -44517 -81761
rect -44473 -81805 -44017 -81761
rect -43973 -81805 -43917 -81761
rect -43873 -81805 -43817 -81761
rect -43773 -81805 -43717 -81761
rect -43673 -81805 -43617 -81761
rect -43573 -81805 -43517 -81761
rect -43473 -81805 -43417 -81761
rect -43373 -81805 -43317 -81761
rect -43273 -81805 -43217 -81761
rect -43173 -81805 -43117 -81761
rect -43073 -81805 -43017 -81761
rect -42973 -81805 -42917 -81761
rect -42873 -81805 -42817 -81761
rect -42773 -81805 -42717 -81761
rect -42673 -81805 -42617 -81761
rect -42573 -81805 -42517 -81761
rect -42473 -81799 80737 -81761
rect 80781 -81799 80837 -81755
rect 80881 -81799 80937 -81755
rect 80981 -81799 81037 -81755
rect 81081 -81799 81137 -81755
rect 81181 -81799 81237 -81755
rect 81281 -81799 81337 -81755
rect 81381 -81799 81437 -81755
rect 81481 -81799 81537 -81755
rect 81581 -81799 81637 -81755
rect 81681 -81799 81737 -81755
rect 81781 -81799 81837 -81755
rect 81881 -81799 81937 -81755
rect 81981 -81799 82037 -81755
rect 82081 -81799 82137 -81755
rect 82181 -81799 82237 -81755
rect 82281 -81799 82737 -81755
rect 82781 -81799 82837 -81755
rect 82881 -81799 82937 -81755
rect 82981 -81799 83037 -81755
rect 83081 -81799 83137 -81755
rect 83181 -81799 83237 -81755
rect 83281 -81799 83337 -81755
rect 83381 -81799 83437 -81755
rect 83481 -81799 83537 -81755
rect 83581 -81799 83637 -81755
rect 83681 -81799 83737 -81755
rect 83781 -81799 83837 -81755
rect 83881 -81799 83937 -81755
rect 83981 -81799 84037 -81755
rect 84081 -81799 84137 -81755
rect 84181 -81799 84237 -81755
rect 84281 -81799 84737 -81755
rect 84781 -81799 84837 -81755
rect 84881 -81799 84937 -81755
rect 84981 -81799 85037 -81755
rect 85081 -81799 85137 -81755
rect 85181 -81799 85237 -81755
rect 85281 -81799 85337 -81755
rect 85381 -81799 85437 -81755
rect 85481 -81799 85537 -81755
rect 85581 -81799 85637 -81755
rect 85681 -81799 85737 -81755
rect 85781 -81799 85837 -81755
rect 85881 -81799 85937 -81755
rect 85981 -81799 86037 -81755
rect 86081 -81799 86137 -81755
rect 86181 -81799 86237 -81755
rect 86281 -81799 86737 -81755
rect 86781 -81799 86837 -81755
rect 86881 -81799 86937 -81755
rect 86981 -81799 87037 -81755
rect 87081 -81799 87137 -81755
rect 87181 -81799 87237 -81755
rect 87281 -81799 87337 -81755
rect 87381 -81799 87437 -81755
rect 87481 -81799 87537 -81755
rect 87581 -81799 87637 -81755
rect 87681 -81799 87737 -81755
rect 87781 -81799 87837 -81755
rect 87881 -81799 87937 -81755
rect 87981 -81799 88037 -81755
rect 88081 -81799 88137 -81755
rect 88181 -81799 88237 -81755
rect 88281 -81799 177360 -81755
rect -42473 -81805 177360 -81799
rect -109116 -81855 177360 -81805
rect -109116 -81859 80737 -81855
rect -109116 -81903 -82968 -81859
rect -82924 -81903 -82868 -81859
rect -82824 -81903 -82768 -81859
rect -82724 -81903 -82668 -81859
rect -82624 -81903 -82568 -81859
rect -82524 -81903 -82468 -81859
rect -82424 -81903 -82368 -81859
rect -82324 -81903 -82268 -81859
rect -82224 -81903 -82168 -81859
rect -82124 -81903 -82068 -81859
rect -82024 -81903 -81968 -81859
rect -81924 -81903 -81868 -81859
rect -81824 -81903 -81768 -81859
rect -81724 -81903 -81668 -81859
rect -81624 -81903 -81568 -81859
rect -81524 -81903 -81468 -81859
rect -81424 -81903 -80968 -81859
rect -80924 -81903 -80868 -81859
rect -80824 -81903 -80768 -81859
rect -80724 -81903 -80668 -81859
rect -80624 -81903 -80568 -81859
rect -80524 -81903 -80468 -81859
rect -80424 -81903 -80368 -81859
rect -80324 -81903 -80268 -81859
rect -80224 -81903 -80168 -81859
rect -80124 -81903 -80068 -81859
rect -80024 -81903 -79968 -81859
rect -79924 -81903 -79868 -81859
rect -79824 -81903 -79768 -81859
rect -79724 -81903 -79668 -81859
rect -79624 -81903 -79568 -81859
rect -79524 -81903 -79468 -81859
rect -79424 -81903 -78968 -81859
rect -78924 -81903 -78868 -81859
rect -78824 -81903 -78768 -81859
rect -78724 -81903 -78668 -81859
rect -78624 -81903 -78568 -81859
rect -78524 -81903 -78468 -81859
rect -78424 -81903 -78368 -81859
rect -78324 -81903 -78268 -81859
rect -78224 -81903 -78168 -81859
rect -78124 -81903 -78068 -81859
rect -78024 -81903 -77968 -81859
rect -77924 -81903 -77868 -81859
rect -77824 -81903 -77768 -81859
rect -77724 -81903 -77668 -81859
rect -77624 -81903 -77568 -81859
rect -77524 -81903 -77468 -81859
rect -77424 -81903 -76968 -81859
rect -76924 -81903 -76868 -81859
rect -76824 -81903 -76768 -81859
rect -76724 -81903 -76668 -81859
rect -76624 -81903 -76568 -81859
rect -76524 -81903 -76468 -81859
rect -76424 -81903 -76368 -81859
rect -76324 -81903 -76268 -81859
rect -76224 -81903 -76168 -81859
rect -76124 -81903 -76068 -81859
rect -76024 -81903 -75968 -81859
rect -75924 -81903 -75868 -81859
rect -75824 -81903 -75768 -81859
rect -75724 -81903 -75668 -81859
rect -75624 -81903 -75568 -81859
rect -75524 -81903 -75468 -81859
rect -75424 -81861 80737 -81859
rect -75424 -81903 -50017 -81861
rect -109116 -81905 -50017 -81903
rect -49973 -81905 -49917 -81861
rect -49873 -81905 -49817 -81861
rect -49773 -81905 -49717 -81861
rect -49673 -81905 -49617 -81861
rect -49573 -81905 -49517 -81861
rect -49473 -81905 -49417 -81861
rect -49373 -81905 -49317 -81861
rect -49273 -81905 -49217 -81861
rect -49173 -81905 -49117 -81861
rect -49073 -81905 -49017 -81861
rect -48973 -81905 -48917 -81861
rect -48873 -81905 -48817 -81861
rect -48773 -81905 -48717 -81861
rect -48673 -81905 -48617 -81861
rect -48573 -81905 -48517 -81861
rect -48473 -81905 -48017 -81861
rect -47973 -81905 -47917 -81861
rect -47873 -81905 -47817 -81861
rect -47773 -81905 -47717 -81861
rect -47673 -81905 -47617 -81861
rect -47573 -81905 -47517 -81861
rect -47473 -81905 -47417 -81861
rect -47373 -81905 -47317 -81861
rect -47273 -81905 -47217 -81861
rect -47173 -81905 -47117 -81861
rect -47073 -81905 -47017 -81861
rect -46973 -81905 -46917 -81861
rect -46873 -81905 -46817 -81861
rect -46773 -81905 -46717 -81861
rect -46673 -81905 -46617 -81861
rect -46573 -81905 -46517 -81861
rect -46473 -81905 -46017 -81861
rect -45973 -81905 -45917 -81861
rect -45873 -81905 -45817 -81861
rect -45773 -81905 -45717 -81861
rect -45673 -81905 -45617 -81861
rect -45573 -81905 -45517 -81861
rect -45473 -81905 -45417 -81861
rect -45373 -81905 -45317 -81861
rect -45273 -81905 -45217 -81861
rect -45173 -81905 -45117 -81861
rect -45073 -81905 -45017 -81861
rect -44973 -81905 -44917 -81861
rect -44873 -81905 -44817 -81861
rect -44773 -81905 -44717 -81861
rect -44673 -81905 -44617 -81861
rect -44573 -81905 -44517 -81861
rect -44473 -81905 -44017 -81861
rect -43973 -81905 -43917 -81861
rect -43873 -81905 -43817 -81861
rect -43773 -81905 -43717 -81861
rect -43673 -81905 -43617 -81861
rect -43573 -81905 -43517 -81861
rect -43473 -81905 -43417 -81861
rect -43373 -81905 -43317 -81861
rect -43273 -81905 -43217 -81861
rect -43173 -81905 -43117 -81861
rect -43073 -81905 -43017 -81861
rect -42973 -81905 -42917 -81861
rect -42873 -81905 -42817 -81861
rect -42773 -81905 -42717 -81861
rect -42673 -81905 -42617 -81861
rect -42573 -81905 -42517 -81861
rect -42473 -81899 80737 -81861
rect 80781 -81899 80837 -81855
rect 80881 -81899 80937 -81855
rect 80981 -81899 81037 -81855
rect 81081 -81899 81137 -81855
rect 81181 -81899 81237 -81855
rect 81281 -81899 81337 -81855
rect 81381 -81899 81437 -81855
rect 81481 -81899 81537 -81855
rect 81581 -81899 81637 -81855
rect 81681 -81899 81737 -81855
rect 81781 -81899 81837 -81855
rect 81881 -81899 81937 -81855
rect 81981 -81899 82037 -81855
rect 82081 -81899 82137 -81855
rect 82181 -81899 82237 -81855
rect 82281 -81899 82737 -81855
rect 82781 -81899 82837 -81855
rect 82881 -81899 82937 -81855
rect 82981 -81899 83037 -81855
rect 83081 -81899 83137 -81855
rect 83181 -81899 83237 -81855
rect 83281 -81899 83337 -81855
rect 83381 -81899 83437 -81855
rect 83481 -81899 83537 -81855
rect 83581 -81899 83637 -81855
rect 83681 -81899 83737 -81855
rect 83781 -81899 83837 -81855
rect 83881 -81899 83937 -81855
rect 83981 -81899 84037 -81855
rect 84081 -81899 84137 -81855
rect 84181 -81899 84237 -81855
rect 84281 -81899 84737 -81855
rect 84781 -81899 84837 -81855
rect 84881 -81899 84937 -81855
rect 84981 -81899 85037 -81855
rect 85081 -81899 85137 -81855
rect 85181 -81899 85237 -81855
rect 85281 -81899 85337 -81855
rect 85381 -81899 85437 -81855
rect 85481 -81899 85537 -81855
rect 85581 -81899 85637 -81855
rect 85681 -81899 85737 -81855
rect 85781 -81899 85837 -81855
rect 85881 -81899 85937 -81855
rect 85981 -81899 86037 -81855
rect 86081 -81899 86137 -81855
rect 86181 -81899 86237 -81855
rect 86281 -81899 86737 -81855
rect 86781 -81899 86837 -81855
rect 86881 -81899 86937 -81855
rect 86981 -81899 87037 -81855
rect 87081 -81899 87137 -81855
rect 87181 -81899 87237 -81855
rect 87281 -81899 87337 -81855
rect 87381 -81899 87437 -81855
rect 87481 -81899 87537 -81855
rect 87581 -81899 87637 -81855
rect 87681 -81899 87737 -81855
rect 87781 -81899 87837 -81855
rect 87881 -81899 87937 -81855
rect 87981 -81899 88037 -81855
rect 88081 -81899 88137 -81855
rect 88181 -81899 88237 -81855
rect 88281 -81899 177360 -81855
rect -42473 -81905 177360 -81899
rect -109116 -81955 177360 -81905
rect -109116 -81959 80737 -81955
rect -109116 -82003 -82968 -81959
rect -82924 -82003 -82868 -81959
rect -82824 -82003 -82768 -81959
rect -82724 -82003 -82668 -81959
rect -82624 -82003 -82568 -81959
rect -82524 -82003 -82468 -81959
rect -82424 -82003 -82368 -81959
rect -82324 -82003 -82268 -81959
rect -82224 -82003 -82168 -81959
rect -82124 -82003 -82068 -81959
rect -82024 -82003 -81968 -81959
rect -81924 -82003 -81868 -81959
rect -81824 -82003 -81768 -81959
rect -81724 -82003 -81668 -81959
rect -81624 -82003 -81568 -81959
rect -81524 -82003 -81468 -81959
rect -81424 -82003 -80968 -81959
rect -80924 -82003 -80868 -81959
rect -80824 -82003 -80768 -81959
rect -80724 -82003 -80668 -81959
rect -80624 -82003 -80568 -81959
rect -80524 -82003 -80468 -81959
rect -80424 -82003 -80368 -81959
rect -80324 -82003 -80268 -81959
rect -80224 -82003 -80168 -81959
rect -80124 -82003 -80068 -81959
rect -80024 -82003 -79968 -81959
rect -79924 -82003 -79868 -81959
rect -79824 -82003 -79768 -81959
rect -79724 -82003 -79668 -81959
rect -79624 -82003 -79568 -81959
rect -79524 -82003 -79468 -81959
rect -79424 -82003 -78968 -81959
rect -78924 -82003 -78868 -81959
rect -78824 -82003 -78768 -81959
rect -78724 -82003 -78668 -81959
rect -78624 -82003 -78568 -81959
rect -78524 -82003 -78468 -81959
rect -78424 -82003 -78368 -81959
rect -78324 -82003 -78268 -81959
rect -78224 -82003 -78168 -81959
rect -78124 -82003 -78068 -81959
rect -78024 -82003 -77968 -81959
rect -77924 -82003 -77868 -81959
rect -77824 -82003 -77768 -81959
rect -77724 -82003 -77668 -81959
rect -77624 -82003 -77568 -81959
rect -77524 -82003 -77468 -81959
rect -77424 -82003 -76968 -81959
rect -76924 -82003 -76868 -81959
rect -76824 -82003 -76768 -81959
rect -76724 -82003 -76668 -81959
rect -76624 -82003 -76568 -81959
rect -76524 -82003 -76468 -81959
rect -76424 -82003 -76368 -81959
rect -76324 -82003 -76268 -81959
rect -76224 -82003 -76168 -81959
rect -76124 -82003 -76068 -81959
rect -76024 -82003 -75968 -81959
rect -75924 -82003 -75868 -81959
rect -75824 -82003 -75768 -81959
rect -75724 -82003 -75668 -81959
rect -75624 -82003 -75568 -81959
rect -75524 -82003 -75468 -81959
rect -75424 -81961 80737 -81959
rect -75424 -82003 -50017 -81961
rect -109116 -82005 -50017 -82003
rect -49973 -82005 -49917 -81961
rect -49873 -82005 -49817 -81961
rect -49773 -82005 -49717 -81961
rect -49673 -82005 -49617 -81961
rect -49573 -82005 -49517 -81961
rect -49473 -82005 -49417 -81961
rect -49373 -82005 -49317 -81961
rect -49273 -82005 -49217 -81961
rect -49173 -82005 -49117 -81961
rect -49073 -82005 -49017 -81961
rect -48973 -82005 -48917 -81961
rect -48873 -82005 -48817 -81961
rect -48773 -82005 -48717 -81961
rect -48673 -82005 -48617 -81961
rect -48573 -82005 -48517 -81961
rect -48473 -82005 -48017 -81961
rect -47973 -82005 -47917 -81961
rect -47873 -82005 -47817 -81961
rect -47773 -82005 -47717 -81961
rect -47673 -82005 -47617 -81961
rect -47573 -82005 -47517 -81961
rect -47473 -82005 -47417 -81961
rect -47373 -82005 -47317 -81961
rect -47273 -82005 -47217 -81961
rect -47173 -82005 -47117 -81961
rect -47073 -82005 -47017 -81961
rect -46973 -82005 -46917 -81961
rect -46873 -82005 -46817 -81961
rect -46773 -82005 -46717 -81961
rect -46673 -82005 -46617 -81961
rect -46573 -82005 -46517 -81961
rect -46473 -82005 -46017 -81961
rect -45973 -82005 -45917 -81961
rect -45873 -82005 -45817 -81961
rect -45773 -82005 -45717 -81961
rect -45673 -82005 -45617 -81961
rect -45573 -82005 -45517 -81961
rect -45473 -82005 -45417 -81961
rect -45373 -82005 -45317 -81961
rect -45273 -82005 -45217 -81961
rect -45173 -82005 -45117 -81961
rect -45073 -82005 -45017 -81961
rect -44973 -82005 -44917 -81961
rect -44873 -82005 -44817 -81961
rect -44773 -82005 -44717 -81961
rect -44673 -82005 -44617 -81961
rect -44573 -82005 -44517 -81961
rect -44473 -82005 -44017 -81961
rect -43973 -82005 -43917 -81961
rect -43873 -82005 -43817 -81961
rect -43773 -82005 -43717 -81961
rect -43673 -82005 -43617 -81961
rect -43573 -82005 -43517 -81961
rect -43473 -82005 -43417 -81961
rect -43373 -82005 -43317 -81961
rect -43273 -82005 -43217 -81961
rect -43173 -82005 -43117 -81961
rect -43073 -82005 -43017 -81961
rect -42973 -82005 -42917 -81961
rect -42873 -82005 -42817 -81961
rect -42773 -82005 -42717 -81961
rect -42673 -82005 -42617 -81961
rect -42573 -82005 -42517 -81961
rect -42473 -81999 80737 -81961
rect 80781 -81999 80837 -81955
rect 80881 -81999 80937 -81955
rect 80981 -81999 81037 -81955
rect 81081 -81999 81137 -81955
rect 81181 -81999 81237 -81955
rect 81281 -81999 81337 -81955
rect 81381 -81999 81437 -81955
rect 81481 -81999 81537 -81955
rect 81581 -81999 81637 -81955
rect 81681 -81999 81737 -81955
rect 81781 -81999 81837 -81955
rect 81881 -81999 81937 -81955
rect 81981 -81999 82037 -81955
rect 82081 -81999 82137 -81955
rect 82181 -81999 82237 -81955
rect 82281 -81999 82737 -81955
rect 82781 -81999 82837 -81955
rect 82881 -81999 82937 -81955
rect 82981 -81999 83037 -81955
rect 83081 -81999 83137 -81955
rect 83181 -81999 83237 -81955
rect 83281 -81999 83337 -81955
rect 83381 -81999 83437 -81955
rect 83481 -81999 83537 -81955
rect 83581 -81999 83637 -81955
rect 83681 -81999 83737 -81955
rect 83781 -81999 83837 -81955
rect 83881 -81999 83937 -81955
rect 83981 -81999 84037 -81955
rect 84081 -81999 84137 -81955
rect 84181 -81999 84237 -81955
rect 84281 -81999 84737 -81955
rect 84781 -81999 84837 -81955
rect 84881 -81999 84937 -81955
rect 84981 -81999 85037 -81955
rect 85081 -81999 85137 -81955
rect 85181 -81999 85237 -81955
rect 85281 -81999 85337 -81955
rect 85381 -81999 85437 -81955
rect 85481 -81999 85537 -81955
rect 85581 -81999 85637 -81955
rect 85681 -81999 85737 -81955
rect 85781 -81999 85837 -81955
rect 85881 -81999 85937 -81955
rect 85981 -81999 86037 -81955
rect 86081 -81999 86137 -81955
rect 86181 -81999 86237 -81955
rect 86281 -81999 86737 -81955
rect 86781 -81999 86837 -81955
rect 86881 -81999 86937 -81955
rect 86981 -81999 87037 -81955
rect 87081 -81999 87137 -81955
rect 87181 -81999 87237 -81955
rect 87281 -81999 87337 -81955
rect 87381 -81999 87437 -81955
rect 87481 -81999 87537 -81955
rect 87581 -81999 87637 -81955
rect 87681 -81999 87737 -81955
rect 87781 -81999 87837 -81955
rect 87881 -81999 87937 -81955
rect 87981 -81999 88037 -81955
rect 88081 -81999 88137 -81955
rect 88181 -81999 88237 -81955
rect 88281 -81999 177360 -81955
rect -42473 -82005 177360 -81999
rect -109116 -82203 177360 -82005
rect -109116 -83117 -109040 -82203
rect -108508 -83117 -108432 -82203
rect -107900 -83117 -107824 -82203
rect -107292 -83117 -107216 -82203
rect -106684 -83117 -106608 -82203
rect -106076 -83117 -106000 -82203
rect -105468 -83117 -105392 -82203
rect -104860 -83117 -104784 -82203
rect -104252 -83117 -104176 -82203
rect -103644 -83117 -103568 -82203
rect -103036 -83117 -102960 -82203
rect -102428 -83117 -102352 -82203
rect -101820 -83117 -101744 -82203
rect -101212 -83117 -101136 -82203
rect -100604 -83117 -100528 -82203
rect -99996 -83117 -99920 -82203
rect -99388 -83117 -99312 -82203
rect -98780 -83117 -98704 -82203
rect -98172 -83117 -98096 -82203
rect -97564 -83117 -97488 -82203
rect -96956 -83117 -96880 -82203
rect -96348 -83117 -96272 -82203
rect -95740 -83117 -95664 -82203
rect -95132 -83117 -95056 -82203
rect -94524 -83117 -94448 -82203
rect -93916 -83117 -93840 -82203
rect -93308 -83117 -93232 -82203
rect -92700 -83117 -92624 -82203
rect -92092 -83117 -92016 -82203
rect -91484 -83117 -91408 -82203
rect -90876 -83117 -90800 -82203
rect -90268 -83117 -90192 -82203
rect -89660 -83117 -89584 -82203
rect -89052 -83117 -88976 -82203
rect -88444 -83117 -88368 -82203
rect -87836 -83117 -87760 -82203
rect -87228 -83117 -87152 -82203
rect -86620 -83117 -86544 -82203
rect -86012 -83117 -85936 -82203
rect -85404 -83117 -85328 -82203
rect -84796 -83117 -84720 -82203
rect -84188 -83117 -84112 -82203
rect -83580 -83117 -83504 -82203
rect -82972 -83117 -82896 -82203
rect -82364 -83117 -82288 -82203
rect -81756 -83117 -81680 -82203
rect -81148 -83117 -81072 -82203
rect -80540 -83117 -80464 -82203
rect -79932 -83117 -79856 -82203
rect -79324 -83117 -79248 -82203
rect -78716 -83117 -78640 -82203
rect -77116 -83117 -77040 -82203
rect -76508 -83117 -76432 -82203
rect -75900 -83117 -75824 -82203
rect -75292 -83117 -75216 -82203
rect -74684 -83117 -74608 -82203
rect -74076 -83117 -74000 -82203
rect -73468 -83117 -73392 -82203
rect -72860 -83117 -72784 -82203
rect -72252 -83117 -72176 -82203
rect -71644 -83117 -71568 -82203
rect -71036 -83117 -70960 -82203
rect -70428 -83117 -70352 -82203
rect -69820 -83117 -69744 -82203
rect -69212 -83117 -69136 -82203
rect -68604 -83117 -68528 -82203
rect -67996 -83117 -67920 -82203
rect -67388 -83117 -67312 -82203
rect -66780 -83117 -66704 -82203
rect -66172 -83117 -66096 -82203
rect -65564 -83117 -65488 -82203
rect -64956 -83117 -64880 -82203
rect -64348 -83117 -64272 -82203
rect -63740 -83117 -63664 -82203
rect -63132 -83117 -63056 -82203
rect -62524 -83117 -62448 -82203
rect -61916 -83117 -61840 -82203
rect -61308 -83117 -61232 -82203
rect -60700 -83117 -60624 -82203
rect -60092 -83117 -60016 -82203
rect -59484 -83117 -59408 -82203
rect -58876 -83117 -58800 -82203
rect -58268 -83117 -58192 -82203
rect -57660 -83117 -57584 -82203
rect -57052 -83117 -56976 -82203
rect -56444 -83117 -56368 -82203
rect -55836 -83117 -55760 -82203
rect -55228 -83117 -55152 -82203
rect -54620 -83117 -54544 -82203
rect -54012 -83117 -53936 -82203
rect -53404 -83117 -53328 -82203
rect -52796 -83117 -52720 -82203
rect -52188 -83117 -52112 -82203
rect -51580 -83117 -51504 -82203
rect -50972 -83117 -50896 -82203
rect -50364 -83117 -50288 -82203
rect -49756 -83117 -49680 -82203
rect -49148 -83117 -49072 -82203
rect -48540 -83117 -48464 -82203
rect -47932 -83117 -47856 -82203
rect -47324 -83117 -47248 -82203
rect -46716 -83117 -46640 -82203
rect -45116 -83117 -45040 -82203
rect -44508 -83117 -44432 -82203
rect -43900 -83117 -43824 -82203
rect -43292 -83117 -43216 -82203
rect -42684 -83117 -42608 -82203
rect -42076 -83117 -42000 -82203
rect -41468 -83117 -41392 -82203
rect -40860 -83117 -40784 -82203
rect -40252 -83117 -40176 -82203
rect -39644 -83117 -39568 -82203
rect -39036 -83117 -38960 -82203
rect -38428 -83117 -38352 -82203
rect -37820 -83117 -37744 -82203
rect -37212 -83117 -37136 -82203
rect -36604 -83117 -36528 -82203
rect -35996 -83117 -35920 -82203
rect -35388 -83117 -35312 -82203
rect -34780 -83117 -34704 -82203
rect -34172 -83117 -34096 -82203
rect -33564 -83117 -33488 -82203
rect -32956 -83117 -32880 -82203
rect -32348 -83117 -32272 -82203
rect -31740 -83117 -31664 -82203
rect -31132 -83117 -31056 -82203
rect -30524 -83117 -30448 -82203
rect -29916 -83117 -29840 -82203
rect -29308 -83117 -29232 -82203
rect -28700 -83117 -28624 -82203
rect -28092 -83117 -28016 -82203
rect -27484 -83117 -27408 -82203
rect -26876 -83117 -26800 -82203
rect -26268 -83117 -26192 -82203
rect -25660 -83117 -25584 -82203
rect -25052 -83117 -24976 -82203
rect -24444 -83117 -24368 -82203
rect -23836 -83117 -23760 -82203
rect -23228 -83117 -23152 -82203
rect -22620 -83117 -22544 -82203
rect -22012 -83117 -21936 -82203
rect -21404 -83117 -21328 -82203
rect -20796 -83117 -20720 -82203
rect -20188 -83117 -20112 -82203
rect -19580 -83117 -19504 -82203
rect -18972 -83117 -18896 -82203
rect -18364 -83117 -18288 -82203
rect -17756 -83117 -17680 -82203
rect -17148 -83117 -17072 -82203
rect -16540 -83117 -16464 -82203
rect -15932 -83117 -15856 -82203
rect -15324 -83117 -15248 -82203
rect -14716 -83117 -14640 -82203
rect -13116 -83117 -13040 -82203
rect -12508 -83117 -12432 -82203
rect -11900 -83117 -11824 -82203
rect -11292 -83117 -11216 -82203
rect -10684 -83117 -10608 -82203
rect -10076 -83117 -10000 -82203
rect -9468 -83117 -9392 -82203
rect -8860 -83117 -8784 -82203
rect -8252 -83117 -8176 -82203
rect -7644 -83117 -7568 -82203
rect -7036 -83117 -6960 -82203
rect -6428 -83117 -6352 -82203
rect -5820 -83117 -5744 -82203
rect -5212 -83117 -5136 -82203
rect -4604 -83117 -4528 -82203
rect -3996 -83117 -3920 -82203
rect -3388 -83117 -3312 -82203
rect -2780 -83117 -2704 -82203
rect -2172 -83117 -2096 -82203
rect -1564 -83117 -1488 -82203
rect -956 -83117 -880 -82203
rect -348 -83117 -272 -82203
rect 260 -83117 336 -82203
rect 868 -83117 944 -82203
rect 1476 -83117 1552 -82203
rect 2084 -83117 2160 -82203
rect 2692 -83117 2768 -82203
rect 3300 -83117 3376 -82203
rect 3908 -83117 3984 -82203
rect 4516 -83117 4592 -82203
rect 5124 -83117 5200 -82203
rect 5732 -83117 5808 -82203
rect 6340 -83117 6416 -82203
rect 6948 -83117 7024 -82203
rect 7556 -83117 7632 -82203
rect 8164 -83117 8240 -82203
rect 8772 -83117 8848 -82203
rect 9380 -83117 9456 -82203
rect 9988 -83117 10064 -82203
rect 10596 -83117 10672 -82203
rect 11204 -83117 11280 -82203
rect 11812 -83117 11888 -82203
rect 12420 -83117 12496 -82203
rect 13028 -83117 13104 -82203
rect 13636 -83117 13712 -82203
rect 14244 -83117 14320 -82203
rect 14852 -83117 14928 -82203
rect 15460 -83117 15536 -82203
rect 16068 -83117 16144 -82203
rect 16676 -83117 16752 -82203
rect 17284 -83117 17360 -82203
rect 18884 -83117 18960 -82203
rect 19492 -83117 19568 -82203
rect 20100 -83117 20176 -82203
rect 20708 -83117 20784 -82203
rect 21316 -83117 21392 -82203
rect 21924 -83117 22000 -82203
rect 22532 -83117 22608 -82203
rect 23140 -83117 23216 -82203
rect 23748 -83117 23824 -82203
rect 24356 -83117 24432 -82203
rect 24964 -83117 25040 -82203
rect 25572 -83117 25648 -82203
rect 26180 -83117 26256 -82203
rect 26788 -83117 26864 -82203
rect 27396 -83117 27472 -82203
rect 28004 -83117 28080 -82203
rect 28612 -83117 28688 -82203
rect 29220 -83117 29296 -82203
rect 29828 -83117 29904 -82203
rect 30436 -83117 30512 -82203
rect 31044 -83117 31120 -82203
rect 31652 -83117 31728 -82203
rect 32260 -83117 32336 -82203
rect 32868 -83117 32944 -82203
rect 33476 -83117 33552 -82203
rect 34084 -83117 34160 -82203
rect 34692 -83117 34768 -82203
rect 35300 -83117 35376 -82203
rect 35908 -83117 35984 -82203
rect 36516 -83117 36592 -82203
rect 37124 -83117 37200 -82203
rect 37732 -83117 37808 -82203
rect 38340 -83117 38416 -82203
rect 38948 -83117 39024 -82203
rect 39556 -83117 39632 -82203
rect 40164 -83117 40240 -82203
rect 40772 -83117 40848 -82203
rect 41380 -83117 41456 -82203
rect 41988 -83117 42064 -82203
rect 42596 -83117 42672 -82203
rect 43204 -83117 43280 -82203
rect 43812 -83117 43888 -82203
rect 44420 -83117 44496 -82203
rect 45028 -83117 45104 -82203
rect 45636 -83117 45712 -82203
rect 46244 -83117 46320 -82203
rect 46852 -83117 46928 -82203
rect 47460 -83117 47536 -82203
rect 48068 -83117 48144 -82203
rect 48676 -83117 48752 -82203
rect 49284 -83117 49360 -82203
rect 50884 -83117 50960 -82203
rect 51492 -83117 51568 -82203
rect 52100 -83117 52176 -82203
rect 52708 -83117 52784 -82203
rect 53316 -83117 53392 -82203
rect 53924 -83117 54000 -82203
rect 54532 -83117 54608 -82203
rect 55140 -83117 55216 -82203
rect 55748 -83117 55824 -82203
rect 56356 -83117 56432 -82203
rect 56964 -83117 57040 -82203
rect 57572 -83117 57648 -82203
rect 58180 -83117 58256 -82203
rect 58788 -83117 58864 -82203
rect 59396 -83117 59472 -82203
rect 60004 -83117 60080 -82203
rect 60612 -83117 60688 -82203
rect 61220 -83117 61296 -82203
rect 61828 -83117 61904 -82203
rect 62436 -83117 62512 -82203
rect 63044 -83117 63120 -82203
rect 63652 -83117 63728 -82203
rect 64260 -83117 64336 -82203
rect 64868 -83117 64944 -82203
rect 65476 -83117 65552 -82203
rect 66084 -83117 66160 -82203
rect 66692 -83117 66768 -82203
rect 67300 -83117 67376 -82203
rect 67908 -83117 67984 -82203
rect 68516 -83117 68592 -82203
rect 69124 -83117 69200 -82203
rect 69732 -83117 69808 -82203
rect 70340 -83117 70416 -82203
rect 70948 -83117 71024 -82203
rect 71556 -83117 71632 -82203
rect 72164 -83117 72240 -82203
rect 72772 -83117 72848 -82203
rect 73380 -83117 73456 -82203
rect 73988 -83117 74064 -82203
rect 74596 -83117 74672 -82203
rect 75204 -83117 75280 -82203
rect 75812 -83117 75888 -82203
rect 76420 -83117 76496 -82203
rect 77028 -83117 77104 -82203
rect 77636 -83117 77712 -82203
rect 78244 -83117 78320 -82203
rect 78852 -83117 78928 -82203
rect 79460 -83117 79536 -82203
rect 80068 -83117 80144 -82203
rect 80676 -83117 80752 -82203
rect 81284 -83117 81360 -82203
rect 82884 -83117 82960 -82203
rect 83492 -83117 83568 -82203
rect 84100 -83117 84176 -82203
rect 84708 -83117 84784 -82203
rect 85316 -83117 85392 -82203
rect 85924 -83117 86000 -82203
rect 86532 -83117 86608 -82203
rect 87140 -83117 87216 -82203
rect 87748 -83117 87824 -82203
rect 88356 -83117 88432 -82203
rect 88964 -83117 89040 -82203
rect 89572 -83117 89648 -82203
rect 90180 -83117 90256 -82203
rect 90788 -83117 90864 -82203
rect 91396 -83117 91472 -82203
rect 92004 -83117 92080 -82203
rect 92612 -83117 92688 -82203
rect 93220 -83117 93296 -82203
rect 93828 -83117 93904 -82203
rect 94436 -83117 94512 -82203
rect 95044 -83117 95120 -82203
rect 95652 -83117 95728 -82203
rect 96260 -83117 96336 -82203
rect 96868 -83117 96944 -82203
rect 97476 -83117 97552 -82203
rect 98084 -83117 98160 -82203
rect 98692 -83117 98768 -82203
rect 99300 -83117 99376 -82203
rect 99908 -83117 99984 -82203
rect 100516 -83117 100592 -82203
rect 101124 -83117 101200 -82203
rect 101732 -83117 101808 -82203
rect 102340 -83117 102416 -82203
rect 102948 -83117 103024 -82203
rect 103556 -83117 103632 -82203
rect 104164 -83117 104240 -82203
rect 104772 -83117 104848 -82203
rect 105380 -83117 105456 -82203
rect 105988 -83117 106064 -82203
rect 106596 -83117 106672 -82203
rect 107204 -83117 107280 -82203
rect 107812 -83117 107888 -82203
rect 108420 -83117 108496 -82203
rect 109028 -83117 109104 -82203
rect 109636 -83117 109712 -82203
rect 110244 -83117 110320 -82203
rect 110852 -83117 110928 -82203
rect 111460 -83117 111536 -82203
rect 112068 -83117 112144 -82203
rect 112676 -83117 112752 -82203
rect 113284 -83117 113360 -82203
rect 114884 -83117 114960 -82203
rect 115492 -83117 115568 -82203
rect 116100 -83117 116176 -82203
rect 116708 -83117 116784 -82203
rect 117316 -83117 117392 -82203
rect 117924 -83117 118000 -82203
rect 118532 -83117 118608 -82203
rect 119140 -83117 119216 -82203
rect 119748 -83117 119824 -82203
rect 120356 -83117 120432 -82203
rect 120964 -83117 121040 -82203
rect 121572 -83117 121648 -82203
rect 122180 -83117 122256 -82203
rect 122788 -83117 122864 -82203
rect 123396 -83117 123472 -82203
rect 124004 -83117 124080 -82203
rect 124612 -83117 124688 -82203
rect 125220 -83117 125296 -82203
rect 125828 -83117 125904 -82203
rect 126436 -83117 126512 -82203
rect 127044 -83117 127120 -82203
rect 127652 -83117 127728 -82203
rect 128260 -83117 128336 -82203
rect 128868 -83117 128944 -82203
rect 129476 -83117 129552 -82203
rect 130084 -83117 130160 -82203
rect 130692 -83117 130768 -82203
rect 131300 -83117 131376 -82203
rect 131908 -83117 131984 -82203
rect 132516 -83117 132592 -82203
rect 133124 -83117 133200 -82203
rect 133732 -83117 133808 -82203
rect 134340 -83117 134416 -82203
rect 134948 -83117 135024 -82203
rect 135556 -83117 135632 -82203
rect 136164 -83117 136240 -82203
rect 136772 -83117 136848 -82203
rect 137380 -83117 137456 -82203
rect 137988 -83117 138064 -82203
rect 138596 -83117 138672 -82203
rect 139204 -83117 139280 -82203
rect 139812 -83117 139888 -82203
rect 140420 -83117 140496 -82203
rect 141028 -83117 141104 -82203
rect 141636 -83117 141712 -82203
rect 142244 -83117 142320 -82203
rect 142852 -83117 142928 -82203
rect 143460 -83117 143536 -82203
rect 144068 -83117 144144 -82203
rect 144676 -83117 144752 -82203
rect 145284 -83117 145360 -82203
rect 146884 -83117 146960 -82203
rect 147492 -83117 147568 -82203
rect 148100 -83117 148176 -82203
rect 148708 -83117 148784 -82203
rect 149316 -83117 149392 -82203
rect 149924 -83117 150000 -82203
rect 150532 -83117 150608 -82203
rect 151140 -83117 151216 -82203
rect 151748 -83117 151824 -82203
rect 152356 -83117 152432 -82203
rect 152964 -83117 153040 -82203
rect 153572 -83117 153648 -82203
rect 154180 -83117 154256 -82203
rect 154788 -83117 154864 -82203
rect 155396 -83117 155472 -82203
rect 156004 -83117 156080 -82203
rect 156612 -83117 156688 -82203
rect 157220 -83117 157296 -82203
rect 157828 -83117 157904 -82203
rect 158436 -83117 158512 -82203
rect 159044 -83117 159120 -82203
rect 159652 -83117 159728 -82203
rect 160260 -83117 160336 -82203
rect 160868 -83117 160944 -82203
rect 161476 -83117 161552 -82203
rect 162084 -83117 162160 -82203
rect 162692 -83117 162768 -82203
rect 163300 -83117 163376 -82203
rect 163908 -83117 163984 -82203
rect 164516 -83117 164592 -82203
rect 165124 -83117 165200 -82203
rect 165732 -83117 165808 -82203
rect 166340 -83117 166416 -82203
rect 166948 -83117 167024 -82203
rect 167556 -83117 167632 -82203
rect 168164 -83117 168240 -82203
rect 168772 -83117 168848 -82203
rect 169380 -83117 169456 -82203
rect 169988 -83117 170064 -82203
rect 170596 -83117 170672 -82203
rect 171204 -83117 171280 -82203
rect 171812 -83117 171888 -82203
rect 172420 -83117 172496 -82203
rect 173028 -83117 173104 -82203
rect 173636 -83117 173712 -82203
rect 174244 -83117 174320 -82203
rect 174852 -83117 174928 -82203
rect 175460 -83117 175536 -82203
rect 176068 -83117 176144 -82203
rect 176676 -83117 176752 -82203
rect 177284 -83117 177360 -82203
rect -77274 -103121 -77040 -83119
rect -45274 -103121 -45040 -83119
rect -13274 -103121 -13040 -83119
rect 18726 -103121 18960 -83119
rect 50726 -103121 50960 -83119
rect 82726 -103121 82960 -83119
rect 114726 -103121 114960 -83119
rect 146726 -103121 146960 -83119
rect 183526 -95506 188605 -92059
rect 183526 -96423 185033 -95506
rect 185843 -96423 188605 -95506
rect 183526 -98092 188605 -96423
rect -108812 -104035 -108736 -103121
rect -108204 -104035 -108128 -103121
rect -107596 -104035 -107520 -103121
rect -106988 -104035 -106912 -103121
rect -106380 -104035 -106304 -103121
rect -105772 -104035 -105696 -103121
rect -105164 -104035 -105088 -103121
rect -104556 -104035 -104480 -103121
rect -103948 -104035 -103872 -103121
rect -103340 -104035 -103264 -103121
rect -102732 -104035 -102656 -103121
rect -102124 -104035 -102048 -103121
rect -101516 -104035 -101440 -103121
rect -100908 -104035 -100832 -103121
rect -100300 -104035 -100224 -103121
rect -99692 -104035 -99616 -103121
rect -99084 -104035 -99008 -103121
rect -98476 -104035 -98400 -103121
rect -97868 -104035 -97792 -103121
rect -97260 -104035 -97184 -103121
rect -96652 -104035 -96576 -103121
rect -96044 -104035 -95968 -103121
rect -95436 -104035 -95360 -103121
rect -94828 -104035 -94752 -103121
rect -94220 -104035 -94144 -103121
rect -93612 -104035 -93536 -103121
rect -93004 -104035 -92928 -103121
rect -92396 -104035 -92320 -103121
rect -91788 -104035 -91712 -103121
rect -91180 -104035 -91104 -103121
rect -90572 -104035 -90496 -103121
rect -89964 -104035 -89888 -103121
rect -89356 -104035 -89280 -103121
rect -88748 -104035 -88672 -103121
rect -88140 -104035 -88064 -103121
rect -87532 -104035 -87456 -103121
rect -86924 -104035 -86848 -103121
rect -86316 -104035 -86240 -103121
rect -85708 -104035 -85632 -103121
rect -85100 -104035 -85024 -103121
rect -84492 -104035 -84416 -103121
rect -83884 -104035 -83808 -103121
rect -83276 -104035 -83200 -103121
rect -82668 -104035 -82592 -103121
rect -82060 -104035 -81984 -103121
rect -81452 -104035 -81376 -103121
rect -80844 -104035 -80768 -103121
rect -80236 -104035 -80160 -103121
rect -79628 -104035 -79552 -103121
rect -79020 -104035 -78944 -103121
rect -76812 -104035 -76736 -103121
rect -76204 -104035 -76128 -103121
rect -75596 -104035 -75520 -103121
rect -74988 -104035 -74912 -103121
rect -74380 -104035 -74304 -103121
rect -73772 -104035 -73696 -103121
rect -73164 -104035 -73088 -103121
rect -72556 -104035 -72480 -103121
rect -71948 -104035 -71872 -103121
rect -71340 -104035 -71264 -103121
rect -70732 -104035 -70656 -103121
rect -70124 -104035 -70048 -103121
rect -69516 -104035 -69440 -103121
rect -68908 -104035 -68832 -103121
rect -68300 -104035 -68224 -103121
rect -67692 -104035 -67616 -103121
rect -67084 -104035 -67008 -103121
rect -66476 -104035 -66400 -103121
rect -65868 -104035 -65792 -103121
rect -65260 -104035 -65184 -103121
rect -64652 -104035 -64576 -103121
rect -64044 -104035 -63968 -103121
rect -63436 -104035 -63360 -103121
rect -62828 -104035 -62752 -103121
rect -62220 -104035 -62144 -103121
rect -61612 -104035 -61536 -103121
rect -61004 -104035 -60928 -103121
rect -60396 -104035 -60320 -103121
rect -59788 -104035 -59712 -103121
rect -59180 -104035 -59104 -103121
rect -58572 -104035 -58496 -103121
rect -57964 -104035 -57888 -103121
rect -57356 -104035 -57280 -103121
rect -56748 -104035 -56672 -103121
rect -56140 -104035 -56064 -103121
rect -55532 -104035 -55456 -103121
rect -54924 -104035 -54848 -103121
rect -54316 -104035 -54240 -103121
rect -53708 -104035 -53632 -103121
rect -53100 -104035 -53024 -103121
rect -52492 -104035 -52416 -103121
rect -51884 -104035 -51808 -103121
rect -51276 -104035 -51200 -103121
rect -50668 -104035 -50592 -103121
rect -50060 -104035 -49984 -103121
rect -49452 -104035 -49376 -103121
rect -48844 -104035 -48768 -103121
rect -48236 -104035 -48160 -103121
rect -47628 -104035 -47552 -103121
rect -47020 -104035 -46944 -103121
rect -44812 -104035 -44736 -103121
rect -44204 -104035 -44128 -103121
rect -43596 -104035 -43520 -103121
rect -42988 -104035 -42912 -103121
rect -42380 -104035 -42304 -103121
rect -41772 -104035 -41696 -103121
rect -41164 -104035 -41088 -103121
rect -40556 -104035 -40480 -103121
rect -39948 -104035 -39872 -103121
rect -39340 -104035 -39264 -103121
rect -38732 -104035 -38656 -103121
rect -38124 -104035 -38048 -103121
rect -37516 -104035 -37440 -103121
rect -36908 -104035 -36832 -103121
rect -36300 -104035 -36224 -103121
rect -35692 -104035 -35616 -103121
rect -35084 -104035 -35008 -103121
rect -34476 -104035 -34400 -103121
rect -33868 -104035 -33792 -103121
rect -33260 -104035 -33184 -103121
rect -32652 -104035 -32576 -103121
rect -32044 -104035 -31968 -103121
rect -31436 -104035 -31360 -103121
rect -30828 -104035 -30752 -103121
rect -30220 -104035 -30144 -103121
rect -29612 -104035 -29536 -103121
rect -29004 -104035 -28928 -103121
rect -28396 -104035 -28320 -103121
rect -27788 -104035 -27712 -103121
rect -27180 -104035 -27104 -103121
rect -26572 -104035 -26496 -103121
rect -25964 -104035 -25888 -103121
rect -25356 -104035 -25280 -103121
rect -24748 -104035 -24672 -103121
rect -24140 -104035 -24064 -103121
rect -23532 -104035 -23456 -103121
rect -22924 -104035 -22848 -103121
rect -22316 -104035 -22240 -103121
rect -21708 -104035 -21632 -103121
rect -21100 -104035 -21024 -103121
rect -20492 -104035 -20416 -103121
rect -19884 -104035 -19808 -103121
rect -19276 -104035 -19200 -103121
rect -18668 -104035 -18592 -103121
rect -18060 -104035 -17984 -103121
rect -17452 -104035 -17376 -103121
rect -16844 -104035 -16768 -103121
rect -16236 -104035 -16160 -103121
rect -15628 -104035 -15552 -103121
rect -15020 -104035 -14944 -103121
rect -12812 -104035 -12736 -103121
rect -12204 -104035 -12128 -103121
rect -11596 -104035 -11520 -103121
rect -10988 -104035 -10912 -103121
rect -10380 -104035 -10304 -103121
rect -9772 -104035 -9696 -103121
rect -9164 -104035 -9088 -103121
rect -8556 -104035 -8480 -103121
rect -7948 -104035 -7872 -103121
rect -7340 -104035 -7264 -103121
rect -6732 -104035 -6656 -103121
rect -6124 -104035 -6048 -103121
rect -5516 -104035 -5440 -103121
rect -4908 -104035 -4832 -103121
rect -4300 -104035 -4224 -103121
rect -3692 -104035 -3616 -103121
rect -3084 -104035 -3008 -103121
rect -2476 -104035 -2400 -103121
rect -1868 -104035 -1792 -103121
rect -1260 -104035 -1184 -103121
rect -652 -104035 -576 -103121
rect -44 -104035 32 -103121
rect 564 -104035 640 -103121
rect 1172 -104035 1248 -103121
rect 1780 -104035 1856 -103121
rect 2388 -104035 2464 -103121
rect 2996 -104035 3072 -103121
rect 3604 -104035 3680 -103121
rect 4212 -104035 4288 -103121
rect 4820 -104035 4896 -103121
rect 5428 -104035 5504 -103121
rect 6036 -104035 6112 -103121
rect 6644 -104035 6720 -103121
rect 7252 -104035 7328 -103121
rect 7860 -104035 7936 -103121
rect 8468 -104035 8544 -103121
rect 9076 -104035 9152 -103121
rect 9684 -104035 9760 -103121
rect 10292 -104035 10368 -103121
rect 10900 -104035 10976 -103121
rect 11508 -104035 11584 -103121
rect 12116 -104035 12192 -103121
rect 12724 -104035 12800 -103121
rect 13332 -104035 13408 -103121
rect 13940 -104035 14016 -103121
rect 14548 -104035 14624 -103121
rect 15156 -104035 15232 -103121
rect 15764 -104035 15840 -103121
rect 16372 -104035 16448 -103121
rect 16980 -104035 17056 -103121
rect 19188 -104035 19264 -103121
rect 19796 -104035 19872 -103121
rect 20404 -104035 20480 -103121
rect 21012 -104035 21088 -103121
rect 21620 -104035 21696 -103121
rect 22228 -104035 22304 -103121
rect 22836 -104035 22912 -103121
rect 23444 -104035 23520 -103121
rect 24052 -104035 24128 -103121
rect 24660 -104035 24736 -103121
rect 25268 -104035 25344 -103121
rect 25876 -104035 25952 -103121
rect 26484 -104035 26560 -103121
rect 27092 -104035 27168 -103121
rect 27700 -104035 27776 -103121
rect 28308 -104035 28384 -103121
rect 28916 -104035 28992 -103121
rect 29524 -104035 29600 -103121
rect 30132 -104035 30208 -103121
rect 30740 -104035 30816 -103121
rect 31348 -104035 31424 -103121
rect 31956 -104035 32032 -103121
rect 32564 -104035 32640 -103121
rect 33172 -104035 33248 -103121
rect 33780 -104035 33856 -103121
rect 34388 -104035 34464 -103121
rect 34996 -104035 35072 -103121
rect 35604 -104035 35680 -103121
rect 36212 -104035 36288 -103121
rect 36820 -104035 36896 -103121
rect 37428 -104035 37504 -103121
rect 38036 -104035 38112 -103121
rect 38644 -104035 38720 -103121
rect 39252 -104035 39328 -103121
rect 39860 -104035 39936 -103121
rect 40468 -104035 40544 -103121
rect 41076 -104035 41152 -103121
rect 41684 -104035 41760 -103121
rect 42292 -104035 42368 -103121
rect 42900 -104035 42976 -103121
rect 43508 -104035 43584 -103121
rect 44116 -104035 44192 -103121
rect 44724 -104035 44800 -103121
rect 45332 -104035 45408 -103121
rect 45940 -104035 46016 -103121
rect 46548 -104035 46624 -103121
rect 47156 -104035 47232 -103121
rect 47764 -104035 47840 -103121
rect 48372 -104035 48448 -103121
rect 48980 -104035 49056 -103121
rect 51188 -104035 51264 -103121
rect 51796 -104035 51872 -103121
rect 52404 -104035 52480 -103121
rect 53012 -104035 53088 -103121
rect 53620 -104035 53696 -103121
rect 54228 -104035 54304 -103121
rect 54836 -104035 54912 -103121
rect 55444 -104035 55520 -103121
rect 56052 -104035 56128 -103121
rect 56660 -104035 56736 -103121
rect 57268 -104035 57344 -103121
rect 57876 -104035 57952 -103121
rect 58484 -104035 58560 -103121
rect 59092 -104035 59168 -103121
rect 59700 -104035 59776 -103121
rect 60308 -104035 60384 -103121
rect 60916 -104035 60992 -103121
rect 61524 -104035 61600 -103121
rect 62132 -104035 62208 -103121
rect 62740 -104035 62816 -103121
rect 63348 -104035 63424 -103121
rect 63956 -104035 64032 -103121
rect 64564 -104035 64640 -103121
rect 65172 -104035 65248 -103121
rect 65780 -104035 65856 -103121
rect 66388 -104035 66464 -103121
rect 66996 -104035 67072 -103121
rect 67604 -104035 67680 -103121
rect 68212 -104035 68288 -103121
rect 68820 -104035 68896 -103121
rect 69428 -104035 69504 -103121
rect 70036 -104035 70112 -103121
rect 70644 -104035 70720 -103121
rect 71252 -104035 71328 -103121
rect 71860 -104035 71936 -103121
rect 72468 -104035 72544 -103121
rect 73076 -104035 73152 -103121
rect 73684 -104035 73760 -103121
rect 74292 -104035 74368 -103121
rect 74900 -104035 74976 -103121
rect 75508 -104035 75584 -103121
rect 76116 -104035 76192 -103121
rect 76724 -104035 76800 -103121
rect 77332 -104035 77408 -103121
rect 77940 -104035 78016 -103121
rect 78548 -104035 78624 -103121
rect 79156 -104035 79232 -103121
rect 79764 -104035 79840 -103121
rect 80372 -104035 80448 -103121
rect 80980 -104035 81056 -103121
rect 83188 -104035 83264 -103121
rect 83796 -104035 83872 -103121
rect 84404 -104035 84480 -103121
rect 85012 -104035 85088 -103121
rect 85620 -104035 85696 -103121
rect 86228 -104035 86304 -103121
rect 86836 -104035 86912 -103121
rect 87444 -104035 87520 -103121
rect 88052 -104035 88128 -103121
rect 88660 -104035 88736 -103121
rect 89268 -104035 89344 -103121
rect 89876 -104035 89952 -103121
rect 90484 -104035 90560 -103121
rect 91092 -104035 91168 -103121
rect 91700 -104035 91776 -103121
rect 92308 -104035 92384 -103121
rect 92916 -104035 92992 -103121
rect 93524 -104035 93600 -103121
rect 94132 -104035 94208 -103121
rect 94740 -104035 94816 -103121
rect 95348 -104035 95424 -103121
rect 95956 -104035 96032 -103121
rect 96564 -104035 96640 -103121
rect 97172 -104035 97248 -103121
rect 97780 -104035 97856 -103121
rect 98388 -104035 98464 -103121
rect 98996 -104035 99072 -103121
rect 99604 -104035 99680 -103121
rect 100212 -104035 100288 -103121
rect 100820 -104035 100896 -103121
rect 101428 -104035 101504 -103121
rect 102036 -104035 102112 -103121
rect 102644 -104035 102720 -103121
rect 103252 -104035 103328 -103121
rect 103860 -104035 103936 -103121
rect 104468 -104035 104544 -103121
rect 105076 -104035 105152 -103121
rect 105684 -104035 105760 -103121
rect 106292 -104035 106368 -103121
rect 106900 -104035 106976 -103121
rect 107508 -104035 107584 -103121
rect 108116 -104035 108192 -103121
rect 108724 -104035 108800 -103121
rect 109332 -104035 109408 -103121
rect 109940 -104035 110016 -103121
rect 110548 -104035 110624 -103121
rect 111156 -104035 111232 -103121
rect 111764 -104035 111840 -103121
rect 112372 -104035 112448 -103121
rect 112980 -104035 113056 -103121
rect 115188 -104035 115264 -103121
rect 115796 -104035 115872 -103121
rect 116404 -104035 116480 -103121
rect 117012 -104035 117088 -103121
rect 117620 -104035 117696 -103121
rect 118228 -104035 118304 -103121
rect 118836 -104035 118912 -103121
rect 119444 -104035 119520 -103121
rect 120052 -104035 120128 -103121
rect 120660 -104035 120736 -103121
rect 121268 -104035 121344 -103121
rect 121876 -104035 121952 -103121
rect 122484 -104035 122560 -103121
rect 123092 -104035 123168 -103121
rect 123700 -104035 123776 -103121
rect 124308 -104035 124384 -103121
rect 124916 -104035 124992 -103121
rect 125524 -104035 125600 -103121
rect 126132 -104035 126208 -103121
rect 126740 -104035 126816 -103121
rect 127348 -104035 127424 -103121
rect 127956 -104035 128032 -103121
rect 128564 -104035 128640 -103121
rect 129172 -104035 129248 -103121
rect 129780 -104035 129856 -103121
rect 130388 -104035 130464 -103121
rect 130996 -104035 131072 -103121
rect 131604 -104035 131680 -103121
rect 132212 -104035 132288 -103121
rect 132820 -104035 132896 -103121
rect 133428 -104035 133504 -103121
rect 134036 -104035 134112 -103121
rect 134644 -104035 134720 -103121
rect 135252 -104035 135328 -103121
rect 135860 -104035 135936 -103121
rect 136468 -104035 136544 -103121
rect 137076 -104035 137152 -103121
rect 137684 -104035 137760 -103121
rect 138292 -104035 138368 -103121
rect 138900 -104035 138976 -103121
rect 139508 -104035 139584 -103121
rect 140116 -104035 140192 -103121
rect 140724 -104035 140800 -103121
rect 141332 -104035 141408 -103121
rect 141940 -104035 142016 -103121
rect 142548 -104035 142624 -103121
rect 143156 -104035 143232 -103121
rect 143764 -104035 143840 -103121
rect 144372 -104035 144448 -103121
rect 144980 -104035 145056 -103121
rect 147188 -104035 147264 -103121
rect 147796 -104035 147872 -103121
rect 148404 -104035 148480 -103121
rect 149012 -104035 149088 -103121
rect 149620 -104035 149696 -103121
rect 150228 -104035 150304 -103121
rect 150836 -104035 150912 -103121
rect 151444 -104035 151520 -103121
rect 152052 -104035 152128 -103121
rect 152660 -104035 152736 -103121
rect 153268 -104035 153344 -103121
rect 153876 -104035 153952 -103121
rect 154484 -104035 154560 -103121
rect 155092 -104035 155168 -103121
rect 155700 -104035 155776 -103121
rect 156308 -104035 156384 -103121
rect 156916 -104035 156992 -103121
rect 157524 -104035 157600 -103121
rect 158132 -104035 158208 -103121
rect 158740 -104035 158816 -103121
rect 159348 -104035 159424 -103121
rect 159956 -104035 160032 -103121
rect 160564 -104035 160640 -103121
rect 161172 -104035 161248 -103121
rect 161780 -104035 161856 -103121
rect 162388 -104035 162464 -103121
rect 162996 -104035 163072 -103121
rect 163604 -104035 163680 -103121
rect 164212 -104035 164288 -103121
rect 164820 -104035 164896 -103121
rect 165428 -104035 165504 -103121
rect 166036 -104035 166112 -103121
rect 166644 -104035 166720 -103121
rect 167252 -104035 167328 -103121
rect 167860 -104035 167936 -103121
rect 168468 -104035 168544 -103121
rect 169076 -104035 169152 -103121
rect 169684 -104035 169760 -103121
rect 170292 -104035 170368 -103121
rect 170900 -104035 170976 -103121
rect 171508 -104035 171584 -103121
rect 172116 -104035 172192 -103121
rect 172724 -104035 172800 -103121
rect 173332 -104035 173408 -103121
rect 173940 -104035 174016 -103121
rect 174548 -104035 174624 -103121
rect 175156 -104035 175232 -103121
rect 175764 -104035 175840 -103121
rect 176372 -104035 176448 -103121
rect 176980 -104035 177056 -103121
rect -108812 -104602 178308 -104035
rect -50768 -106193 -42000 -105630
rect -50768 -106237 -50075 -106193
rect -50031 -106237 -49975 -106193
rect -49931 -106237 -49875 -106193
rect -49831 -106237 -49775 -106193
rect -49731 -106237 -49675 -106193
rect -49631 -106237 -49575 -106193
rect -49531 -106237 -49475 -106193
rect -49431 -106237 -49375 -106193
rect -49331 -106237 -49275 -106193
rect -49231 -106237 -49175 -106193
rect -49131 -106237 -49075 -106193
rect -49031 -106237 -48975 -106193
rect -48931 -106237 -48875 -106193
rect -48831 -106237 -48775 -106193
rect -48731 -106237 -48675 -106193
rect -48631 -106237 -48575 -106193
rect -48531 -106237 -48075 -106193
rect -48031 -106237 -47975 -106193
rect -47931 -106237 -47875 -106193
rect -47831 -106237 -47775 -106193
rect -47731 -106237 -47675 -106193
rect -47631 -106237 -47575 -106193
rect -47531 -106237 -47475 -106193
rect -47431 -106237 -47375 -106193
rect -47331 -106237 -47275 -106193
rect -47231 -106237 -47175 -106193
rect -47131 -106237 -47075 -106193
rect -47031 -106237 -46975 -106193
rect -46931 -106237 -46875 -106193
rect -46831 -106237 -46775 -106193
rect -46731 -106237 -46675 -106193
rect -46631 -106237 -46575 -106193
rect -46531 -106237 -46075 -106193
rect -46031 -106237 -45975 -106193
rect -45931 -106237 -45875 -106193
rect -45831 -106237 -45775 -106193
rect -45731 -106237 -45675 -106193
rect -45631 -106237 -45575 -106193
rect -45531 -106237 -45475 -106193
rect -45431 -106237 -45375 -106193
rect -45331 -106237 -45275 -106193
rect -45231 -106237 -45175 -106193
rect -45131 -106237 -45075 -106193
rect -45031 -106237 -44975 -106193
rect -44931 -106237 -44875 -106193
rect -44831 -106237 -44775 -106193
rect -44731 -106237 -44675 -106193
rect -44631 -106237 -44575 -106193
rect -44531 -106237 -44075 -106193
rect -44031 -106237 -43975 -106193
rect -43931 -106237 -43875 -106193
rect -43831 -106237 -43775 -106193
rect -43731 -106237 -43675 -106193
rect -43631 -106237 -43575 -106193
rect -43531 -106237 -43475 -106193
rect -43431 -106237 -43375 -106193
rect -43331 -106237 -43275 -106193
rect -43231 -106237 -43175 -106193
rect -43131 -106237 -43075 -106193
rect -43031 -106237 -42975 -106193
rect -42931 -106237 -42875 -106193
rect -42831 -106237 -42775 -106193
rect -42731 -106237 -42675 -106193
rect -42631 -106237 -42575 -106193
rect -42531 -106237 -42000 -106193
rect -50768 -106293 -42000 -106237
rect -50768 -106337 -50075 -106293
rect -50031 -106337 -49975 -106293
rect -49931 -106337 -49875 -106293
rect -49831 -106337 -49775 -106293
rect -49731 -106337 -49675 -106293
rect -49631 -106337 -49575 -106293
rect -49531 -106337 -49475 -106293
rect -49431 -106337 -49375 -106293
rect -49331 -106337 -49275 -106293
rect -49231 -106337 -49175 -106293
rect -49131 -106337 -49075 -106293
rect -49031 -106337 -48975 -106293
rect -48931 -106337 -48875 -106293
rect -48831 -106337 -48775 -106293
rect -48731 -106337 -48675 -106293
rect -48631 -106337 -48575 -106293
rect -48531 -106337 -48075 -106293
rect -48031 -106337 -47975 -106293
rect -47931 -106337 -47875 -106293
rect -47831 -106337 -47775 -106293
rect -47731 -106337 -47675 -106293
rect -47631 -106337 -47575 -106293
rect -47531 -106337 -47475 -106293
rect -47431 -106337 -47375 -106293
rect -47331 -106337 -47275 -106293
rect -47231 -106337 -47175 -106293
rect -47131 -106337 -47075 -106293
rect -47031 -106337 -46975 -106293
rect -46931 -106337 -46875 -106293
rect -46831 -106337 -46775 -106293
rect -46731 -106337 -46675 -106293
rect -46631 -106337 -46575 -106293
rect -46531 -106337 -46075 -106293
rect -46031 -106337 -45975 -106293
rect -45931 -106337 -45875 -106293
rect -45831 -106337 -45775 -106293
rect -45731 -106337 -45675 -106293
rect -45631 -106337 -45575 -106293
rect -45531 -106337 -45475 -106293
rect -45431 -106337 -45375 -106293
rect -45331 -106337 -45275 -106293
rect -45231 -106337 -45175 -106293
rect -45131 -106337 -45075 -106293
rect -45031 -106337 -44975 -106293
rect -44931 -106337 -44875 -106293
rect -44831 -106337 -44775 -106293
rect -44731 -106337 -44675 -106293
rect -44631 -106337 -44575 -106293
rect -44531 -106337 -44075 -106293
rect -44031 -106337 -43975 -106293
rect -43931 -106337 -43875 -106293
rect -43831 -106337 -43775 -106293
rect -43731 -106337 -43675 -106293
rect -43631 -106337 -43575 -106293
rect -43531 -106337 -43475 -106293
rect -43431 -106337 -43375 -106293
rect -43331 -106337 -43275 -106293
rect -43231 -106337 -43175 -106293
rect -43131 -106337 -43075 -106293
rect -43031 -106337 -42975 -106293
rect -42931 -106337 -42875 -106293
rect -42831 -106337 -42775 -106293
rect -42731 -106337 -42675 -106293
rect -42631 -106337 -42575 -106293
rect -42531 -106337 -42000 -106293
rect -50768 -106393 -42000 -106337
rect -50768 -106437 -50075 -106393
rect -50031 -106437 -49975 -106393
rect -49931 -106437 -49875 -106393
rect -49831 -106437 -49775 -106393
rect -49731 -106437 -49675 -106393
rect -49631 -106437 -49575 -106393
rect -49531 -106437 -49475 -106393
rect -49431 -106437 -49375 -106393
rect -49331 -106437 -49275 -106393
rect -49231 -106437 -49175 -106393
rect -49131 -106437 -49075 -106393
rect -49031 -106437 -48975 -106393
rect -48931 -106437 -48875 -106393
rect -48831 -106437 -48775 -106393
rect -48731 -106437 -48675 -106393
rect -48631 -106437 -48575 -106393
rect -48531 -106437 -48075 -106393
rect -48031 -106437 -47975 -106393
rect -47931 -106437 -47875 -106393
rect -47831 -106437 -47775 -106393
rect -47731 -106437 -47675 -106393
rect -47631 -106437 -47575 -106393
rect -47531 -106437 -47475 -106393
rect -47431 -106437 -47375 -106393
rect -47331 -106437 -47275 -106393
rect -47231 -106437 -47175 -106393
rect -47131 -106437 -47075 -106393
rect -47031 -106437 -46975 -106393
rect -46931 -106437 -46875 -106393
rect -46831 -106437 -46775 -106393
rect -46731 -106437 -46675 -106393
rect -46631 -106437 -46575 -106393
rect -46531 -106437 -46075 -106393
rect -46031 -106437 -45975 -106393
rect -45931 -106437 -45875 -106393
rect -45831 -106437 -45775 -106393
rect -45731 -106437 -45675 -106393
rect -45631 -106437 -45575 -106393
rect -45531 -106437 -45475 -106393
rect -45431 -106437 -45375 -106393
rect -45331 -106437 -45275 -106393
rect -45231 -106437 -45175 -106393
rect -45131 -106437 -45075 -106393
rect -45031 -106437 -44975 -106393
rect -44931 -106437 -44875 -106393
rect -44831 -106437 -44775 -106393
rect -44731 -106437 -44675 -106393
rect -44631 -106437 -44575 -106393
rect -44531 -106437 -44075 -106393
rect -44031 -106437 -43975 -106393
rect -43931 -106437 -43875 -106393
rect -43831 -106437 -43775 -106393
rect -43731 -106437 -43675 -106393
rect -43631 -106437 -43575 -106393
rect -43531 -106437 -43475 -106393
rect -43431 -106437 -43375 -106393
rect -43331 -106437 -43275 -106393
rect -43231 -106437 -43175 -106393
rect -43131 -106437 -43075 -106393
rect -43031 -106437 -42975 -106393
rect -42931 -106437 -42875 -106393
rect -42831 -106437 -42775 -106393
rect -42731 -106437 -42675 -106393
rect -42631 -106437 -42575 -106393
rect -42531 -106437 -42000 -106393
rect -50768 -106493 -42000 -106437
rect -50768 -106537 -50075 -106493
rect -50031 -106537 -49975 -106493
rect -49931 -106537 -49875 -106493
rect -49831 -106537 -49775 -106493
rect -49731 -106537 -49675 -106493
rect -49631 -106537 -49575 -106493
rect -49531 -106537 -49475 -106493
rect -49431 -106537 -49375 -106493
rect -49331 -106537 -49275 -106493
rect -49231 -106537 -49175 -106493
rect -49131 -106537 -49075 -106493
rect -49031 -106537 -48975 -106493
rect -48931 -106537 -48875 -106493
rect -48831 -106537 -48775 -106493
rect -48731 -106537 -48675 -106493
rect -48631 -106537 -48575 -106493
rect -48531 -106537 -48075 -106493
rect -48031 -106537 -47975 -106493
rect -47931 -106537 -47875 -106493
rect -47831 -106537 -47775 -106493
rect -47731 -106537 -47675 -106493
rect -47631 -106537 -47575 -106493
rect -47531 -106537 -47475 -106493
rect -47431 -106537 -47375 -106493
rect -47331 -106537 -47275 -106493
rect -47231 -106537 -47175 -106493
rect -47131 -106537 -47075 -106493
rect -47031 -106537 -46975 -106493
rect -46931 -106537 -46875 -106493
rect -46831 -106537 -46775 -106493
rect -46731 -106537 -46675 -106493
rect -46631 -106537 -46575 -106493
rect -46531 -106537 -46075 -106493
rect -46031 -106537 -45975 -106493
rect -45931 -106537 -45875 -106493
rect -45831 -106537 -45775 -106493
rect -45731 -106537 -45675 -106493
rect -45631 -106537 -45575 -106493
rect -45531 -106537 -45475 -106493
rect -45431 -106537 -45375 -106493
rect -45331 -106537 -45275 -106493
rect -45231 -106537 -45175 -106493
rect -45131 -106537 -45075 -106493
rect -45031 -106537 -44975 -106493
rect -44931 -106537 -44875 -106493
rect -44831 -106537 -44775 -106493
rect -44731 -106537 -44675 -106493
rect -44631 -106537 -44575 -106493
rect -44531 -106537 -44075 -106493
rect -44031 -106537 -43975 -106493
rect -43931 -106537 -43875 -106493
rect -43831 -106537 -43775 -106493
rect -43731 -106537 -43675 -106493
rect -43631 -106537 -43575 -106493
rect -43531 -106537 -43475 -106493
rect -43431 -106537 -43375 -106493
rect -43331 -106537 -43275 -106493
rect -43231 -106537 -43175 -106493
rect -43131 -106537 -43075 -106493
rect -43031 -106537 -42975 -106493
rect -42931 -106537 -42875 -106493
rect -42831 -106537 -42775 -106493
rect -42731 -106537 -42675 -106493
rect -42631 -106537 -42575 -106493
rect -42531 -106537 -42000 -106493
rect -50768 -106593 -42000 -106537
rect -50768 -106637 -50075 -106593
rect -50031 -106637 -49975 -106593
rect -49931 -106637 -49875 -106593
rect -49831 -106637 -49775 -106593
rect -49731 -106637 -49675 -106593
rect -49631 -106637 -49575 -106593
rect -49531 -106637 -49475 -106593
rect -49431 -106637 -49375 -106593
rect -49331 -106637 -49275 -106593
rect -49231 -106637 -49175 -106593
rect -49131 -106637 -49075 -106593
rect -49031 -106637 -48975 -106593
rect -48931 -106637 -48875 -106593
rect -48831 -106637 -48775 -106593
rect -48731 -106637 -48675 -106593
rect -48631 -106637 -48575 -106593
rect -48531 -106637 -48075 -106593
rect -48031 -106637 -47975 -106593
rect -47931 -106637 -47875 -106593
rect -47831 -106637 -47775 -106593
rect -47731 -106637 -47675 -106593
rect -47631 -106637 -47575 -106593
rect -47531 -106637 -47475 -106593
rect -47431 -106637 -47375 -106593
rect -47331 -106637 -47275 -106593
rect -47231 -106637 -47175 -106593
rect -47131 -106637 -47075 -106593
rect -47031 -106637 -46975 -106593
rect -46931 -106637 -46875 -106593
rect -46831 -106637 -46775 -106593
rect -46731 -106637 -46675 -106593
rect -46631 -106637 -46575 -106593
rect -46531 -106637 -46075 -106593
rect -46031 -106637 -45975 -106593
rect -45931 -106637 -45875 -106593
rect -45831 -106637 -45775 -106593
rect -45731 -106637 -45675 -106593
rect -45631 -106637 -45575 -106593
rect -45531 -106637 -45475 -106593
rect -45431 -106637 -45375 -106593
rect -45331 -106637 -45275 -106593
rect -45231 -106637 -45175 -106593
rect -45131 -106637 -45075 -106593
rect -45031 -106637 -44975 -106593
rect -44931 -106637 -44875 -106593
rect -44831 -106637 -44775 -106593
rect -44731 -106637 -44675 -106593
rect -44631 -106637 -44575 -106593
rect -44531 -106637 -44075 -106593
rect -44031 -106637 -43975 -106593
rect -43931 -106637 -43875 -106593
rect -43831 -106637 -43775 -106593
rect -43731 -106637 -43675 -106593
rect -43631 -106637 -43575 -106593
rect -43531 -106637 -43475 -106593
rect -43431 -106637 -43375 -106593
rect -43331 -106637 -43275 -106593
rect -43231 -106637 -43175 -106593
rect -43131 -106637 -43075 -106593
rect -43031 -106637 -42975 -106593
rect -42931 -106637 -42875 -106593
rect -42831 -106637 -42775 -106593
rect -42731 -106637 -42675 -106593
rect -42631 -106637 -42575 -106593
rect -42531 -106637 -42000 -106593
rect -50768 -106693 -42000 -106637
rect -50768 -106737 -50075 -106693
rect -50031 -106737 -49975 -106693
rect -49931 -106737 -49875 -106693
rect -49831 -106737 -49775 -106693
rect -49731 -106737 -49675 -106693
rect -49631 -106737 -49575 -106693
rect -49531 -106737 -49475 -106693
rect -49431 -106737 -49375 -106693
rect -49331 -106737 -49275 -106693
rect -49231 -106737 -49175 -106693
rect -49131 -106737 -49075 -106693
rect -49031 -106737 -48975 -106693
rect -48931 -106737 -48875 -106693
rect -48831 -106737 -48775 -106693
rect -48731 -106737 -48675 -106693
rect -48631 -106737 -48575 -106693
rect -48531 -106737 -48075 -106693
rect -48031 -106737 -47975 -106693
rect -47931 -106737 -47875 -106693
rect -47831 -106737 -47775 -106693
rect -47731 -106737 -47675 -106693
rect -47631 -106737 -47575 -106693
rect -47531 -106737 -47475 -106693
rect -47431 -106737 -47375 -106693
rect -47331 -106737 -47275 -106693
rect -47231 -106737 -47175 -106693
rect -47131 -106737 -47075 -106693
rect -47031 -106737 -46975 -106693
rect -46931 -106737 -46875 -106693
rect -46831 -106737 -46775 -106693
rect -46731 -106737 -46675 -106693
rect -46631 -106737 -46575 -106693
rect -46531 -106737 -46075 -106693
rect -46031 -106737 -45975 -106693
rect -45931 -106737 -45875 -106693
rect -45831 -106737 -45775 -106693
rect -45731 -106737 -45675 -106693
rect -45631 -106737 -45575 -106693
rect -45531 -106737 -45475 -106693
rect -45431 -106737 -45375 -106693
rect -45331 -106737 -45275 -106693
rect -45231 -106737 -45175 -106693
rect -45131 -106737 -45075 -106693
rect -45031 -106737 -44975 -106693
rect -44931 -106737 -44875 -106693
rect -44831 -106737 -44775 -106693
rect -44731 -106737 -44675 -106693
rect -44631 -106737 -44575 -106693
rect -44531 -106737 -44075 -106693
rect -44031 -106737 -43975 -106693
rect -43931 -106737 -43875 -106693
rect -43831 -106737 -43775 -106693
rect -43731 -106737 -43675 -106693
rect -43631 -106737 -43575 -106693
rect -43531 -106737 -43475 -106693
rect -43431 -106737 -43375 -106693
rect -43331 -106737 -43275 -106693
rect -43231 -106737 -43175 -106693
rect -43131 -106737 -43075 -106693
rect -43031 -106737 -42975 -106693
rect -42931 -106737 -42875 -106693
rect -42831 -106737 -42775 -106693
rect -42731 -106737 -42675 -106693
rect -42631 -106737 -42575 -106693
rect -42531 -106737 -42000 -106693
rect -50768 -106793 -42000 -106737
rect -50768 -106837 -50075 -106793
rect -50031 -106837 -49975 -106793
rect -49931 -106837 -49875 -106793
rect -49831 -106837 -49775 -106793
rect -49731 -106837 -49675 -106793
rect -49631 -106837 -49575 -106793
rect -49531 -106837 -49475 -106793
rect -49431 -106837 -49375 -106793
rect -49331 -106837 -49275 -106793
rect -49231 -106837 -49175 -106793
rect -49131 -106837 -49075 -106793
rect -49031 -106837 -48975 -106793
rect -48931 -106837 -48875 -106793
rect -48831 -106837 -48775 -106793
rect -48731 -106837 -48675 -106793
rect -48631 -106837 -48575 -106793
rect -48531 -106837 -48075 -106793
rect -48031 -106837 -47975 -106793
rect -47931 -106837 -47875 -106793
rect -47831 -106837 -47775 -106793
rect -47731 -106837 -47675 -106793
rect -47631 -106837 -47575 -106793
rect -47531 -106837 -47475 -106793
rect -47431 -106837 -47375 -106793
rect -47331 -106837 -47275 -106793
rect -47231 -106837 -47175 -106793
rect -47131 -106837 -47075 -106793
rect -47031 -106837 -46975 -106793
rect -46931 -106837 -46875 -106793
rect -46831 -106837 -46775 -106793
rect -46731 -106837 -46675 -106793
rect -46631 -106837 -46575 -106793
rect -46531 -106837 -46075 -106793
rect -46031 -106837 -45975 -106793
rect -45931 -106837 -45875 -106793
rect -45831 -106837 -45775 -106793
rect -45731 -106837 -45675 -106793
rect -45631 -106837 -45575 -106793
rect -45531 -106837 -45475 -106793
rect -45431 -106837 -45375 -106793
rect -45331 -106837 -45275 -106793
rect -45231 -106837 -45175 -106793
rect -45131 -106837 -45075 -106793
rect -45031 -106837 -44975 -106793
rect -44931 -106837 -44875 -106793
rect -44831 -106837 -44775 -106793
rect -44731 -106837 -44675 -106793
rect -44631 -106837 -44575 -106793
rect -44531 -106837 -44075 -106793
rect -44031 -106837 -43975 -106793
rect -43931 -106837 -43875 -106793
rect -43831 -106837 -43775 -106793
rect -43731 -106837 -43675 -106793
rect -43631 -106837 -43575 -106793
rect -43531 -106837 -43475 -106793
rect -43431 -106837 -43375 -106793
rect -43331 -106837 -43275 -106793
rect -43231 -106837 -43175 -106793
rect -43131 -106837 -43075 -106793
rect -43031 -106837 -42975 -106793
rect -42931 -106837 -42875 -106793
rect -42831 -106837 -42775 -106793
rect -42731 -106837 -42675 -106793
rect -42631 -106837 -42575 -106793
rect -42531 -106837 -42000 -106793
rect -50768 -106893 -42000 -106837
rect -50768 -106937 -50075 -106893
rect -50031 -106937 -49975 -106893
rect -49931 -106937 -49875 -106893
rect -49831 -106937 -49775 -106893
rect -49731 -106937 -49675 -106893
rect -49631 -106937 -49575 -106893
rect -49531 -106937 -49475 -106893
rect -49431 -106937 -49375 -106893
rect -49331 -106937 -49275 -106893
rect -49231 -106937 -49175 -106893
rect -49131 -106937 -49075 -106893
rect -49031 -106937 -48975 -106893
rect -48931 -106937 -48875 -106893
rect -48831 -106937 -48775 -106893
rect -48731 -106937 -48675 -106893
rect -48631 -106937 -48575 -106893
rect -48531 -106937 -48075 -106893
rect -48031 -106937 -47975 -106893
rect -47931 -106937 -47875 -106893
rect -47831 -106937 -47775 -106893
rect -47731 -106937 -47675 -106893
rect -47631 -106937 -47575 -106893
rect -47531 -106937 -47475 -106893
rect -47431 -106937 -47375 -106893
rect -47331 -106937 -47275 -106893
rect -47231 -106937 -47175 -106893
rect -47131 -106937 -47075 -106893
rect -47031 -106937 -46975 -106893
rect -46931 -106937 -46875 -106893
rect -46831 -106937 -46775 -106893
rect -46731 -106937 -46675 -106893
rect -46631 -106937 -46575 -106893
rect -46531 -106937 -46075 -106893
rect -46031 -106937 -45975 -106893
rect -45931 -106937 -45875 -106893
rect -45831 -106937 -45775 -106893
rect -45731 -106937 -45675 -106893
rect -45631 -106937 -45575 -106893
rect -45531 -106937 -45475 -106893
rect -45431 -106937 -45375 -106893
rect -45331 -106937 -45275 -106893
rect -45231 -106937 -45175 -106893
rect -45131 -106937 -45075 -106893
rect -45031 -106937 -44975 -106893
rect -44931 -106937 -44875 -106893
rect -44831 -106937 -44775 -106893
rect -44731 -106937 -44675 -106893
rect -44631 -106937 -44575 -106893
rect -44531 -106937 -44075 -106893
rect -44031 -106937 -43975 -106893
rect -43931 -106937 -43875 -106893
rect -43831 -106937 -43775 -106893
rect -43731 -106937 -43675 -106893
rect -43631 -106937 -43575 -106893
rect -43531 -106937 -43475 -106893
rect -43431 -106937 -43375 -106893
rect -43331 -106937 -43275 -106893
rect -43231 -106937 -43175 -106893
rect -43131 -106937 -43075 -106893
rect -43031 -106937 -42975 -106893
rect -42931 -106937 -42875 -106893
rect -42831 -106937 -42775 -106893
rect -42731 -106937 -42675 -106893
rect -42631 -106937 -42575 -106893
rect -42531 -106937 -42000 -106893
rect -50768 -106993 -42000 -106937
rect -50768 -107037 -50075 -106993
rect -50031 -107037 -49975 -106993
rect -49931 -107037 -49875 -106993
rect -49831 -107037 -49775 -106993
rect -49731 -107037 -49675 -106993
rect -49631 -107037 -49575 -106993
rect -49531 -107037 -49475 -106993
rect -49431 -107037 -49375 -106993
rect -49331 -107037 -49275 -106993
rect -49231 -107037 -49175 -106993
rect -49131 -107037 -49075 -106993
rect -49031 -107037 -48975 -106993
rect -48931 -107037 -48875 -106993
rect -48831 -107037 -48775 -106993
rect -48731 -107037 -48675 -106993
rect -48631 -107037 -48575 -106993
rect -48531 -107037 -48075 -106993
rect -48031 -107037 -47975 -106993
rect -47931 -107037 -47875 -106993
rect -47831 -107037 -47775 -106993
rect -47731 -107037 -47675 -106993
rect -47631 -107037 -47575 -106993
rect -47531 -107037 -47475 -106993
rect -47431 -107037 -47375 -106993
rect -47331 -107037 -47275 -106993
rect -47231 -107037 -47175 -106993
rect -47131 -107037 -47075 -106993
rect -47031 -107037 -46975 -106993
rect -46931 -107037 -46875 -106993
rect -46831 -107037 -46775 -106993
rect -46731 -107037 -46675 -106993
rect -46631 -107037 -46575 -106993
rect -46531 -107037 -46075 -106993
rect -46031 -107037 -45975 -106993
rect -45931 -107037 -45875 -106993
rect -45831 -107037 -45775 -106993
rect -45731 -107037 -45675 -106993
rect -45631 -107037 -45575 -106993
rect -45531 -107037 -45475 -106993
rect -45431 -107037 -45375 -106993
rect -45331 -107037 -45275 -106993
rect -45231 -107037 -45175 -106993
rect -45131 -107037 -45075 -106993
rect -45031 -107037 -44975 -106993
rect -44931 -107037 -44875 -106993
rect -44831 -107037 -44775 -106993
rect -44731 -107037 -44675 -106993
rect -44631 -107037 -44575 -106993
rect -44531 -107037 -44075 -106993
rect -44031 -107037 -43975 -106993
rect -43931 -107037 -43875 -106993
rect -43831 -107037 -43775 -106993
rect -43731 -107037 -43675 -106993
rect -43631 -107037 -43575 -106993
rect -43531 -107037 -43475 -106993
rect -43431 -107037 -43375 -106993
rect -43331 -107037 -43275 -106993
rect -43231 -107037 -43175 -106993
rect -43131 -107037 -43075 -106993
rect -43031 -107037 -42975 -106993
rect -42931 -107037 -42875 -106993
rect -42831 -107037 -42775 -106993
rect -42731 -107037 -42675 -106993
rect -42631 -107037 -42575 -106993
rect -42531 -107037 -42000 -106993
rect -50768 -107093 -42000 -107037
rect -50768 -107137 -50075 -107093
rect -50031 -107137 -49975 -107093
rect -49931 -107137 -49875 -107093
rect -49831 -107137 -49775 -107093
rect -49731 -107137 -49675 -107093
rect -49631 -107137 -49575 -107093
rect -49531 -107137 -49475 -107093
rect -49431 -107137 -49375 -107093
rect -49331 -107137 -49275 -107093
rect -49231 -107137 -49175 -107093
rect -49131 -107137 -49075 -107093
rect -49031 -107137 -48975 -107093
rect -48931 -107137 -48875 -107093
rect -48831 -107137 -48775 -107093
rect -48731 -107137 -48675 -107093
rect -48631 -107137 -48575 -107093
rect -48531 -107137 -48075 -107093
rect -48031 -107137 -47975 -107093
rect -47931 -107137 -47875 -107093
rect -47831 -107137 -47775 -107093
rect -47731 -107137 -47675 -107093
rect -47631 -107137 -47575 -107093
rect -47531 -107137 -47475 -107093
rect -47431 -107137 -47375 -107093
rect -47331 -107137 -47275 -107093
rect -47231 -107137 -47175 -107093
rect -47131 -107137 -47075 -107093
rect -47031 -107137 -46975 -107093
rect -46931 -107137 -46875 -107093
rect -46831 -107137 -46775 -107093
rect -46731 -107137 -46675 -107093
rect -46631 -107137 -46575 -107093
rect -46531 -107137 -46075 -107093
rect -46031 -107137 -45975 -107093
rect -45931 -107137 -45875 -107093
rect -45831 -107137 -45775 -107093
rect -45731 -107137 -45675 -107093
rect -45631 -107137 -45575 -107093
rect -45531 -107137 -45475 -107093
rect -45431 -107137 -45375 -107093
rect -45331 -107137 -45275 -107093
rect -45231 -107137 -45175 -107093
rect -45131 -107137 -45075 -107093
rect -45031 -107137 -44975 -107093
rect -44931 -107137 -44875 -107093
rect -44831 -107137 -44775 -107093
rect -44731 -107137 -44675 -107093
rect -44631 -107137 -44575 -107093
rect -44531 -107137 -44075 -107093
rect -44031 -107137 -43975 -107093
rect -43931 -107137 -43875 -107093
rect -43831 -107137 -43775 -107093
rect -43731 -107137 -43675 -107093
rect -43631 -107137 -43575 -107093
rect -43531 -107137 -43475 -107093
rect -43431 -107137 -43375 -107093
rect -43331 -107137 -43275 -107093
rect -43231 -107137 -43175 -107093
rect -43131 -107137 -43075 -107093
rect -43031 -107137 -42975 -107093
rect -42931 -107137 -42875 -107093
rect -42831 -107137 -42775 -107093
rect -42731 -107137 -42675 -107093
rect -42631 -107137 -42575 -107093
rect -42531 -107137 -42000 -107093
rect -50768 -107193 -42000 -107137
rect -50768 -107237 -50075 -107193
rect -50031 -107237 -49975 -107193
rect -49931 -107237 -49875 -107193
rect -49831 -107237 -49775 -107193
rect -49731 -107237 -49675 -107193
rect -49631 -107237 -49575 -107193
rect -49531 -107237 -49475 -107193
rect -49431 -107237 -49375 -107193
rect -49331 -107237 -49275 -107193
rect -49231 -107237 -49175 -107193
rect -49131 -107237 -49075 -107193
rect -49031 -107237 -48975 -107193
rect -48931 -107237 -48875 -107193
rect -48831 -107237 -48775 -107193
rect -48731 -107237 -48675 -107193
rect -48631 -107237 -48575 -107193
rect -48531 -107237 -48075 -107193
rect -48031 -107237 -47975 -107193
rect -47931 -107237 -47875 -107193
rect -47831 -107237 -47775 -107193
rect -47731 -107237 -47675 -107193
rect -47631 -107237 -47575 -107193
rect -47531 -107237 -47475 -107193
rect -47431 -107237 -47375 -107193
rect -47331 -107237 -47275 -107193
rect -47231 -107237 -47175 -107193
rect -47131 -107237 -47075 -107193
rect -47031 -107237 -46975 -107193
rect -46931 -107237 -46875 -107193
rect -46831 -107237 -46775 -107193
rect -46731 -107237 -46675 -107193
rect -46631 -107237 -46575 -107193
rect -46531 -107237 -46075 -107193
rect -46031 -107237 -45975 -107193
rect -45931 -107237 -45875 -107193
rect -45831 -107237 -45775 -107193
rect -45731 -107237 -45675 -107193
rect -45631 -107237 -45575 -107193
rect -45531 -107237 -45475 -107193
rect -45431 -107237 -45375 -107193
rect -45331 -107237 -45275 -107193
rect -45231 -107237 -45175 -107193
rect -45131 -107237 -45075 -107193
rect -45031 -107237 -44975 -107193
rect -44931 -107237 -44875 -107193
rect -44831 -107237 -44775 -107193
rect -44731 -107237 -44675 -107193
rect -44631 -107237 -44575 -107193
rect -44531 -107237 -44075 -107193
rect -44031 -107237 -43975 -107193
rect -43931 -107237 -43875 -107193
rect -43831 -107237 -43775 -107193
rect -43731 -107237 -43675 -107193
rect -43631 -107237 -43575 -107193
rect -43531 -107237 -43475 -107193
rect -43431 -107237 -43375 -107193
rect -43331 -107237 -43275 -107193
rect -43231 -107237 -43175 -107193
rect -43131 -107237 -43075 -107193
rect -43031 -107237 -42975 -107193
rect -42931 -107237 -42875 -107193
rect -42831 -107237 -42775 -107193
rect -42731 -107237 -42675 -107193
rect -42631 -107237 -42575 -107193
rect -42531 -107237 -42000 -107193
rect -50768 -107293 -42000 -107237
rect -50768 -107337 -50075 -107293
rect -50031 -107337 -49975 -107293
rect -49931 -107337 -49875 -107293
rect -49831 -107337 -49775 -107293
rect -49731 -107337 -49675 -107293
rect -49631 -107337 -49575 -107293
rect -49531 -107337 -49475 -107293
rect -49431 -107337 -49375 -107293
rect -49331 -107337 -49275 -107293
rect -49231 -107337 -49175 -107293
rect -49131 -107337 -49075 -107293
rect -49031 -107337 -48975 -107293
rect -48931 -107337 -48875 -107293
rect -48831 -107337 -48775 -107293
rect -48731 -107337 -48675 -107293
rect -48631 -107337 -48575 -107293
rect -48531 -107337 -48075 -107293
rect -48031 -107337 -47975 -107293
rect -47931 -107337 -47875 -107293
rect -47831 -107337 -47775 -107293
rect -47731 -107337 -47675 -107293
rect -47631 -107337 -47575 -107293
rect -47531 -107337 -47475 -107293
rect -47431 -107337 -47375 -107293
rect -47331 -107337 -47275 -107293
rect -47231 -107337 -47175 -107293
rect -47131 -107337 -47075 -107293
rect -47031 -107337 -46975 -107293
rect -46931 -107337 -46875 -107293
rect -46831 -107337 -46775 -107293
rect -46731 -107337 -46675 -107293
rect -46631 -107337 -46575 -107293
rect -46531 -107337 -46075 -107293
rect -46031 -107337 -45975 -107293
rect -45931 -107337 -45875 -107293
rect -45831 -107337 -45775 -107293
rect -45731 -107337 -45675 -107293
rect -45631 -107337 -45575 -107293
rect -45531 -107337 -45475 -107293
rect -45431 -107337 -45375 -107293
rect -45331 -107337 -45275 -107293
rect -45231 -107337 -45175 -107293
rect -45131 -107337 -45075 -107293
rect -45031 -107337 -44975 -107293
rect -44931 -107337 -44875 -107293
rect -44831 -107337 -44775 -107293
rect -44731 -107337 -44675 -107293
rect -44631 -107337 -44575 -107293
rect -44531 -107337 -44075 -107293
rect -44031 -107337 -43975 -107293
rect -43931 -107337 -43875 -107293
rect -43831 -107337 -43775 -107293
rect -43731 -107337 -43675 -107293
rect -43631 -107337 -43575 -107293
rect -43531 -107337 -43475 -107293
rect -43431 -107337 -43375 -107293
rect -43331 -107337 -43275 -107293
rect -43231 -107337 -43175 -107293
rect -43131 -107337 -43075 -107293
rect -43031 -107337 -42975 -107293
rect -42931 -107337 -42875 -107293
rect -42831 -107337 -42775 -107293
rect -42731 -107337 -42675 -107293
rect -42631 -107337 -42575 -107293
rect -42531 -107337 -42000 -107293
rect -50768 -107393 -42000 -107337
rect -50768 -107437 -50075 -107393
rect -50031 -107437 -49975 -107393
rect -49931 -107437 -49875 -107393
rect -49831 -107437 -49775 -107393
rect -49731 -107437 -49675 -107393
rect -49631 -107437 -49575 -107393
rect -49531 -107437 -49475 -107393
rect -49431 -107437 -49375 -107393
rect -49331 -107437 -49275 -107393
rect -49231 -107437 -49175 -107393
rect -49131 -107437 -49075 -107393
rect -49031 -107437 -48975 -107393
rect -48931 -107437 -48875 -107393
rect -48831 -107437 -48775 -107393
rect -48731 -107437 -48675 -107393
rect -48631 -107437 -48575 -107393
rect -48531 -107437 -48075 -107393
rect -48031 -107437 -47975 -107393
rect -47931 -107437 -47875 -107393
rect -47831 -107437 -47775 -107393
rect -47731 -107437 -47675 -107393
rect -47631 -107437 -47575 -107393
rect -47531 -107437 -47475 -107393
rect -47431 -107437 -47375 -107393
rect -47331 -107437 -47275 -107393
rect -47231 -107437 -47175 -107393
rect -47131 -107437 -47075 -107393
rect -47031 -107437 -46975 -107393
rect -46931 -107437 -46875 -107393
rect -46831 -107437 -46775 -107393
rect -46731 -107437 -46675 -107393
rect -46631 -107437 -46575 -107393
rect -46531 -107437 -46075 -107393
rect -46031 -107437 -45975 -107393
rect -45931 -107437 -45875 -107393
rect -45831 -107437 -45775 -107393
rect -45731 -107437 -45675 -107393
rect -45631 -107437 -45575 -107393
rect -45531 -107437 -45475 -107393
rect -45431 -107437 -45375 -107393
rect -45331 -107437 -45275 -107393
rect -45231 -107437 -45175 -107393
rect -45131 -107437 -45075 -107393
rect -45031 -107437 -44975 -107393
rect -44931 -107437 -44875 -107393
rect -44831 -107437 -44775 -107393
rect -44731 -107437 -44675 -107393
rect -44631 -107437 -44575 -107393
rect -44531 -107437 -44075 -107393
rect -44031 -107437 -43975 -107393
rect -43931 -107437 -43875 -107393
rect -43831 -107437 -43775 -107393
rect -43731 -107437 -43675 -107393
rect -43631 -107437 -43575 -107393
rect -43531 -107437 -43475 -107393
rect -43431 -107437 -43375 -107393
rect -43331 -107437 -43275 -107393
rect -43231 -107437 -43175 -107393
rect -43131 -107437 -43075 -107393
rect -43031 -107437 -42975 -107393
rect -42931 -107437 -42875 -107393
rect -42831 -107437 -42775 -107393
rect -42731 -107437 -42675 -107393
rect -42631 -107437 -42575 -107393
rect -42531 -107437 -42000 -107393
rect -50768 -107493 -42000 -107437
rect -50768 -107537 -50075 -107493
rect -50031 -107537 -49975 -107493
rect -49931 -107537 -49875 -107493
rect -49831 -107537 -49775 -107493
rect -49731 -107537 -49675 -107493
rect -49631 -107537 -49575 -107493
rect -49531 -107537 -49475 -107493
rect -49431 -107537 -49375 -107493
rect -49331 -107537 -49275 -107493
rect -49231 -107537 -49175 -107493
rect -49131 -107537 -49075 -107493
rect -49031 -107537 -48975 -107493
rect -48931 -107537 -48875 -107493
rect -48831 -107537 -48775 -107493
rect -48731 -107537 -48675 -107493
rect -48631 -107537 -48575 -107493
rect -48531 -107537 -48075 -107493
rect -48031 -107537 -47975 -107493
rect -47931 -107537 -47875 -107493
rect -47831 -107537 -47775 -107493
rect -47731 -107537 -47675 -107493
rect -47631 -107537 -47575 -107493
rect -47531 -107537 -47475 -107493
rect -47431 -107537 -47375 -107493
rect -47331 -107537 -47275 -107493
rect -47231 -107537 -47175 -107493
rect -47131 -107537 -47075 -107493
rect -47031 -107537 -46975 -107493
rect -46931 -107537 -46875 -107493
rect -46831 -107537 -46775 -107493
rect -46731 -107537 -46675 -107493
rect -46631 -107537 -46575 -107493
rect -46531 -107537 -46075 -107493
rect -46031 -107537 -45975 -107493
rect -45931 -107537 -45875 -107493
rect -45831 -107537 -45775 -107493
rect -45731 -107537 -45675 -107493
rect -45631 -107537 -45575 -107493
rect -45531 -107537 -45475 -107493
rect -45431 -107537 -45375 -107493
rect -45331 -107537 -45275 -107493
rect -45231 -107537 -45175 -107493
rect -45131 -107537 -45075 -107493
rect -45031 -107537 -44975 -107493
rect -44931 -107537 -44875 -107493
rect -44831 -107537 -44775 -107493
rect -44731 -107537 -44675 -107493
rect -44631 -107537 -44575 -107493
rect -44531 -107537 -44075 -107493
rect -44031 -107537 -43975 -107493
rect -43931 -107537 -43875 -107493
rect -43831 -107537 -43775 -107493
rect -43731 -107537 -43675 -107493
rect -43631 -107537 -43575 -107493
rect -43531 -107537 -43475 -107493
rect -43431 -107537 -43375 -107493
rect -43331 -107537 -43275 -107493
rect -43231 -107537 -43175 -107493
rect -43131 -107537 -43075 -107493
rect -43031 -107537 -42975 -107493
rect -42931 -107537 -42875 -107493
rect -42831 -107537 -42775 -107493
rect -42731 -107537 -42675 -107493
rect -42631 -107537 -42575 -107493
rect -42531 -107537 -42000 -107493
rect -50768 -107593 -42000 -107537
rect -50768 -107636 -50075 -107593
rect -109116 -107637 -50075 -107636
rect -50031 -107637 -49975 -107593
rect -49931 -107637 -49875 -107593
rect -49831 -107637 -49775 -107593
rect -49731 -107637 -49675 -107593
rect -49631 -107637 -49575 -107593
rect -49531 -107637 -49475 -107593
rect -49431 -107637 -49375 -107593
rect -49331 -107637 -49275 -107593
rect -49231 -107637 -49175 -107593
rect -49131 -107637 -49075 -107593
rect -49031 -107637 -48975 -107593
rect -48931 -107637 -48875 -107593
rect -48831 -107637 -48775 -107593
rect -48731 -107637 -48675 -107593
rect -48631 -107637 -48575 -107593
rect -48531 -107637 -48075 -107593
rect -48031 -107637 -47975 -107593
rect -47931 -107637 -47875 -107593
rect -47831 -107637 -47775 -107593
rect -47731 -107637 -47675 -107593
rect -47631 -107637 -47575 -107593
rect -47531 -107637 -47475 -107593
rect -47431 -107637 -47375 -107593
rect -47331 -107637 -47275 -107593
rect -47231 -107637 -47175 -107593
rect -47131 -107637 -47075 -107593
rect -47031 -107637 -46975 -107593
rect -46931 -107637 -46875 -107593
rect -46831 -107637 -46775 -107593
rect -46731 -107637 -46675 -107593
rect -46631 -107637 -46575 -107593
rect -46531 -107637 -46075 -107593
rect -46031 -107637 -45975 -107593
rect -45931 -107637 -45875 -107593
rect -45831 -107637 -45775 -107593
rect -45731 -107637 -45675 -107593
rect -45631 -107637 -45575 -107593
rect -45531 -107637 -45475 -107593
rect -45431 -107637 -45375 -107593
rect -45331 -107637 -45275 -107593
rect -45231 -107637 -45175 -107593
rect -45131 -107637 -45075 -107593
rect -45031 -107637 -44975 -107593
rect -44931 -107637 -44875 -107593
rect -44831 -107637 -44775 -107593
rect -44731 -107637 -44675 -107593
rect -44631 -107637 -44575 -107593
rect -44531 -107637 -44075 -107593
rect -44031 -107637 -43975 -107593
rect -43931 -107637 -43875 -107593
rect -43831 -107637 -43775 -107593
rect -43731 -107637 -43675 -107593
rect -43631 -107637 -43575 -107593
rect -43531 -107637 -43475 -107593
rect -43431 -107637 -43375 -107593
rect -43331 -107637 -43275 -107593
rect -43231 -107637 -43175 -107593
rect -43131 -107637 -43075 -107593
rect -43031 -107637 -42975 -107593
rect -42931 -107637 -42875 -107593
rect -42831 -107637 -42775 -107593
rect -42731 -107637 -42675 -107593
rect -42631 -107637 -42575 -107593
rect -42531 -107636 -42000 -107593
rect -42531 -107637 177360 -107636
rect -109116 -107693 177360 -107637
rect -109116 -107737 -50075 -107693
rect -50031 -107737 -49975 -107693
rect -49931 -107737 -49875 -107693
rect -49831 -107737 -49775 -107693
rect -49731 -107737 -49675 -107693
rect -49631 -107737 -49575 -107693
rect -49531 -107737 -49475 -107693
rect -49431 -107737 -49375 -107693
rect -49331 -107737 -49275 -107693
rect -49231 -107737 -49175 -107693
rect -49131 -107737 -49075 -107693
rect -49031 -107737 -48975 -107693
rect -48931 -107737 -48875 -107693
rect -48831 -107737 -48775 -107693
rect -48731 -107737 -48675 -107693
rect -48631 -107737 -48575 -107693
rect -48531 -107737 -48075 -107693
rect -48031 -107737 -47975 -107693
rect -47931 -107737 -47875 -107693
rect -47831 -107737 -47775 -107693
rect -47731 -107737 -47675 -107693
rect -47631 -107737 -47575 -107693
rect -47531 -107737 -47475 -107693
rect -47431 -107737 -47375 -107693
rect -47331 -107737 -47275 -107693
rect -47231 -107737 -47175 -107693
rect -47131 -107737 -47075 -107693
rect -47031 -107737 -46975 -107693
rect -46931 -107737 -46875 -107693
rect -46831 -107737 -46775 -107693
rect -46731 -107737 -46675 -107693
rect -46631 -107737 -46575 -107693
rect -46531 -107737 -46075 -107693
rect -46031 -107737 -45975 -107693
rect -45931 -107737 -45875 -107693
rect -45831 -107737 -45775 -107693
rect -45731 -107737 -45675 -107693
rect -45631 -107737 -45575 -107693
rect -45531 -107737 -45475 -107693
rect -45431 -107737 -45375 -107693
rect -45331 -107737 -45275 -107693
rect -45231 -107737 -45175 -107693
rect -45131 -107737 -45075 -107693
rect -45031 -107737 -44975 -107693
rect -44931 -107737 -44875 -107693
rect -44831 -107737 -44775 -107693
rect -44731 -107737 -44675 -107693
rect -44631 -107737 -44575 -107693
rect -44531 -107737 -44075 -107693
rect -44031 -107737 -43975 -107693
rect -43931 -107737 -43875 -107693
rect -43831 -107737 -43775 -107693
rect -43731 -107737 -43675 -107693
rect -43631 -107737 -43575 -107693
rect -43531 -107737 -43475 -107693
rect -43431 -107737 -43375 -107693
rect -43331 -107737 -43275 -107693
rect -43231 -107737 -43175 -107693
rect -43131 -107737 -43075 -107693
rect -43031 -107737 -42975 -107693
rect -42931 -107737 -42875 -107693
rect -42831 -107737 -42775 -107693
rect -42731 -107737 -42675 -107693
rect -42631 -107737 -42575 -107693
rect -42531 -107737 177360 -107693
rect -109116 -108203 177360 -107737
rect -109116 -109117 -109040 -108203
rect -108508 -109117 -108432 -108203
rect -107900 -109117 -107824 -108203
rect -107292 -109117 -107216 -108203
rect -106684 -109117 -106608 -108203
rect -106076 -109117 -106000 -108203
rect -105468 -109117 -105392 -108203
rect -104860 -109117 -104784 -108203
rect -104252 -109117 -104176 -108203
rect -103644 -109117 -103568 -108203
rect -103036 -109117 -102960 -108203
rect -102428 -109117 -102352 -108203
rect -101820 -109117 -101744 -108203
rect -101212 -109117 -101136 -108203
rect -100604 -109117 -100528 -108203
rect -99996 -109117 -99920 -108203
rect -99388 -109117 -99312 -108203
rect -98780 -109117 -98704 -108203
rect -98172 -109117 -98096 -108203
rect -97564 -109117 -97488 -108203
rect -96956 -109117 -96880 -108203
rect -96348 -109117 -96272 -108203
rect -95740 -109117 -95664 -108203
rect -95132 -109117 -95056 -108203
rect -94524 -109117 -94448 -108203
rect -93916 -109117 -93840 -108203
rect -93308 -109117 -93232 -108203
rect -92700 -109117 -92624 -108203
rect -92092 -109117 -92016 -108203
rect -91484 -109117 -91408 -108203
rect -90876 -109117 -90800 -108203
rect -90268 -109117 -90192 -108203
rect -89660 -109117 -89584 -108203
rect -89052 -109117 -88976 -108203
rect -88444 -109117 -88368 -108203
rect -87836 -109117 -87760 -108203
rect -87228 -109117 -87152 -108203
rect -86620 -109117 -86544 -108203
rect -86012 -109117 -85936 -108203
rect -85404 -109117 -85328 -108203
rect -84796 -109117 -84720 -108203
rect -84188 -109117 -84112 -108203
rect -83580 -109117 -83504 -108203
rect -82972 -109117 -82896 -108203
rect -82364 -109117 -82288 -108203
rect -81756 -109117 -81680 -108203
rect -81148 -109117 -81072 -108203
rect -80540 -109117 -80464 -108203
rect -79932 -109117 -79856 -108203
rect -79324 -109117 -79248 -108203
rect -78716 -109117 -78640 -108203
rect -77116 -109117 -77040 -108203
rect -76508 -109117 -76432 -108203
rect -75900 -109117 -75824 -108203
rect -75292 -109117 -75216 -108203
rect -74684 -109117 -74608 -108203
rect -74076 -109117 -74000 -108203
rect -73468 -109117 -73392 -108203
rect -72860 -109117 -72784 -108203
rect -72252 -109117 -72176 -108203
rect -71644 -109117 -71568 -108203
rect -71036 -109117 -70960 -108203
rect -70428 -109117 -70352 -108203
rect -69820 -109117 -69744 -108203
rect -69212 -109117 -69136 -108203
rect -68604 -109117 -68528 -108203
rect -67996 -109117 -67920 -108203
rect -67388 -109117 -67312 -108203
rect -66780 -109117 -66704 -108203
rect -66172 -109117 -66096 -108203
rect -65564 -109117 -65488 -108203
rect -64956 -109117 -64880 -108203
rect -64348 -109117 -64272 -108203
rect -63740 -109117 -63664 -108203
rect -63132 -109117 -63056 -108203
rect -62524 -109117 -62448 -108203
rect -61916 -109117 -61840 -108203
rect -61308 -109117 -61232 -108203
rect -60700 -109117 -60624 -108203
rect -60092 -109117 -60016 -108203
rect -59484 -109117 -59408 -108203
rect -58876 -109117 -58800 -108203
rect -58268 -109117 -58192 -108203
rect -57660 -109117 -57584 -108203
rect -57052 -109117 -56976 -108203
rect -56444 -109117 -56368 -108203
rect -55836 -109117 -55760 -108203
rect -55228 -109117 -55152 -108203
rect -54620 -109117 -54544 -108203
rect -54012 -109117 -53936 -108203
rect -53404 -109117 -53328 -108203
rect -52796 -109117 -52720 -108203
rect -52188 -109117 -52112 -108203
rect -51580 -109117 -51504 -108203
rect -50972 -109117 -50896 -108203
rect -50364 -109117 -50288 -108203
rect -49756 -109117 -49680 -108203
rect -49148 -109117 -49072 -108203
rect -48540 -109117 -48464 -108203
rect -47932 -109117 -47856 -108203
rect -47324 -109117 -47248 -108203
rect -46716 -109117 -46640 -108203
rect -45116 -109117 -45040 -108203
rect -44508 -109117 -44432 -108203
rect -43900 -109117 -43824 -108203
rect -43292 -109117 -43216 -108203
rect -42684 -109117 -42608 -108203
rect -42076 -109117 -42000 -108203
rect -41468 -109117 -41392 -108203
rect -40860 -109117 -40784 -108203
rect -40252 -109117 -40176 -108203
rect -39644 -109117 -39568 -108203
rect -39036 -109117 -38960 -108203
rect -38428 -109117 -38352 -108203
rect -37820 -109117 -37744 -108203
rect -37212 -109117 -37136 -108203
rect -36604 -109117 -36528 -108203
rect -35996 -109117 -35920 -108203
rect -35388 -109117 -35312 -108203
rect -34780 -109117 -34704 -108203
rect -34172 -109117 -34096 -108203
rect -33564 -109117 -33488 -108203
rect -32956 -109117 -32880 -108203
rect -32348 -109117 -32272 -108203
rect -31740 -109117 -31664 -108203
rect -31132 -109117 -31056 -108203
rect -30524 -109117 -30448 -108203
rect -29916 -109117 -29840 -108203
rect -29308 -109117 -29232 -108203
rect -28700 -109117 -28624 -108203
rect -28092 -109117 -28016 -108203
rect -27484 -109117 -27408 -108203
rect -26876 -109117 -26800 -108203
rect -26268 -109117 -26192 -108203
rect -25660 -109117 -25584 -108203
rect -25052 -109117 -24976 -108203
rect -24444 -109117 -24368 -108203
rect -23836 -109117 -23760 -108203
rect -23228 -109117 -23152 -108203
rect -22620 -109117 -22544 -108203
rect -22012 -109117 -21936 -108203
rect -21404 -109117 -21328 -108203
rect -20796 -109117 -20720 -108203
rect -20188 -109117 -20112 -108203
rect -19580 -109117 -19504 -108203
rect -18972 -109117 -18896 -108203
rect -18364 -109117 -18288 -108203
rect -17756 -109117 -17680 -108203
rect -17148 -109117 -17072 -108203
rect -16540 -109117 -16464 -108203
rect -15932 -109117 -15856 -108203
rect -15324 -109117 -15248 -108203
rect -14716 -109117 -14640 -108203
rect -13116 -109117 -13040 -108203
rect -12508 -109117 -12432 -108203
rect -11900 -109117 -11824 -108203
rect -11292 -109117 -11216 -108203
rect -10684 -109117 -10608 -108203
rect -10076 -109117 -10000 -108203
rect -9468 -109117 -9392 -108203
rect -8860 -109117 -8784 -108203
rect -8252 -109117 -8176 -108203
rect -7644 -109117 -7568 -108203
rect -7036 -109117 -6960 -108203
rect -6428 -109117 -6352 -108203
rect -5820 -109117 -5744 -108203
rect -5212 -109117 -5136 -108203
rect -4604 -109117 -4528 -108203
rect -3996 -109117 -3920 -108203
rect -3388 -109117 -3312 -108203
rect -2780 -109117 -2704 -108203
rect -2172 -109117 -2096 -108203
rect -1564 -109117 -1488 -108203
rect -956 -109117 -880 -108203
rect -348 -109117 -272 -108203
rect 260 -109117 336 -108203
rect 868 -109117 944 -108203
rect 1476 -109117 1552 -108203
rect 2084 -109117 2160 -108203
rect 2692 -109117 2768 -108203
rect 3300 -109117 3376 -108203
rect 3908 -109117 3984 -108203
rect 4516 -109117 4592 -108203
rect 5124 -109117 5200 -108203
rect 5732 -109117 5808 -108203
rect 6340 -109117 6416 -108203
rect 6948 -109117 7024 -108203
rect 7556 -109117 7632 -108203
rect 8164 -109117 8240 -108203
rect 8772 -109117 8848 -108203
rect 9380 -109117 9456 -108203
rect 9988 -109117 10064 -108203
rect 10596 -109117 10672 -108203
rect 11204 -109117 11280 -108203
rect 11812 -109117 11888 -108203
rect 12420 -109117 12496 -108203
rect 13028 -109117 13104 -108203
rect 13636 -109117 13712 -108203
rect 14244 -109117 14320 -108203
rect 14852 -109117 14928 -108203
rect 15460 -109117 15536 -108203
rect 16068 -109117 16144 -108203
rect 16676 -109117 16752 -108203
rect 17284 -109117 17360 -108203
rect 18884 -109117 18960 -108203
rect 19492 -109117 19568 -108203
rect 20100 -109117 20176 -108203
rect 20708 -109117 20784 -108203
rect 21316 -109117 21392 -108203
rect 21924 -109117 22000 -108203
rect 22532 -109117 22608 -108203
rect 23140 -109117 23216 -108203
rect 23748 -109117 23824 -108203
rect 24356 -109117 24432 -108203
rect 24964 -109117 25040 -108203
rect 25572 -109117 25648 -108203
rect 26180 -109117 26256 -108203
rect 26788 -109117 26864 -108203
rect 27396 -109117 27472 -108203
rect 28004 -109117 28080 -108203
rect 28612 -109117 28688 -108203
rect 29220 -109117 29296 -108203
rect 29828 -109117 29904 -108203
rect 30436 -109117 30512 -108203
rect 31044 -109117 31120 -108203
rect 31652 -109117 31728 -108203
rect 32260 -109117 32336 -108203
rect 32868 -109117 32944 -108203
rect 33476 -109117 33552 -108203
rect 34084 -109117 34160 -108203
rect 34692 -109117 34768 -108203
rect 35300 -109117 35376 -108203
rect 35908 -109117 35984 -108203
rect 36516 -109117 36592 -108203
rect 37124 -109117 37200 -108203
rect 37732 -109117 37808 -108203
rect 38340 -109117 38416 -108203
rect 38948 -109117 39024 -108203
rect 39556 -109117 39632 -108203
rect 40164 -109117 40240 -108203
rect 40772 -109117 40848 -108203
rect 41380 -109117 41456 -108203
rect 41988 -109117 42064 -108203
rect 42596 -109117 42672 -108203
rect 43204 -109117 43280 -108203
rect 43812 -109117 43888 -108203
rect 44420 -109117 44496 -108203
rect 45028 -109117 45104 -108203
rect 45636 -109117 45712 -108203
rect 46244 -109117 46320 -108203
rect 46852 -109117 46928 -108203
rect 47460 -109117 47536 -108203
rect 48068 -109117 48144 -108203
rect 48676 -109117 48752 -108203
rect 49284 -109117 49360 -108203
rect 50884 -109117 50960 -108203
rect 51492 -109117 51568 -108203
rect 52100 -109117 52176 -108203
rect 52708 -109117 52784 -108203
rect 53316 -109117 53392 -108203
rect 53924 -109117 54000 -108203
rect 54532 -109117 54608 -108203
rect 55140 -109117 55216 -108203
rect 55748 -109117 55824 -108203
rect 56356 -109117 56432 -108203
rect 56964 -109117 57040 -108203
rect 57572 -109117 57648 -108203
rect 58180 -109117 58256 -108203
rect 58788 -109117 58864 -108203
rect 59396 -109117 59472 -108203
rect 60004 -109117 60080 -108203
rect 60612 -109117 60688 -108203
rect 61220 -109117 61296 -108203
rect 61828 -109117 61904 -108203
rect 62436 -109117 62512 -108203
rect 63044 -109117 63120 -108203
rect 63652 -109117 63728 -108203
rect 64260 -109117 64336 -108203
rect 64868 -109117 64944 -108203
rect 65476 -109117 65552 -108203
rect 66084 -109117 66160 -108203
rect 66692 -109117 66768 -108203
rect 67300 -109117 67376 -108203
rect 67908 -109117 67984 -108203
rect 68516 -109117 68592 -108203
rect 69124 -109117 69200 -108203
rect 69732 -109117 69808 -108203
rect 70340 -109117 70416 -108203
rect 70948 -109117 71024 -108203
rect 71556 -109117 71632 -108203
rect 72164 -109117 72240 -108203
rect 72772 -109117 72848 -108203
rect 73380 -109117 73456 -108203
rect 73988 -109117 74064 -108203
rect 74596 -109117 74672 -108203
rect 75204 -109117 75280 -108203
rect 75812 -109117 75888 -108203
rect 76420 -109117 76496 -108203
rect 77028 -109117 77104 -108203
rect 77636 -109117 77712 -108203
rect 78244 -109117 78320 -108203
rect 78852 -109117 78928 -108203
rect 79460 -109117 79536 -108203
rect 80068 -109117 80144 -108203
rect 80676 -109117 80752 -108203
rect 81284 -109117 81360 -108203
rect 82884 -109117 82960 -108203
rect 83492 -109117 83568 -108203
rect 84100 -109117 84176 -108203
rect 84708 -109117 84784 -108203
rect 85316 -109117 85392 -108203
rect 85924 -109117 86000 -108203
rect 86532 -109117 86608 -108203
rect 87140 -109117 87216 -108203
rect 87748 -109117 87824 -108203
rect 88356 -109117 88432 -108203
rect 88964 -109117 89040 -108203
rect 89572 -109117 89648 -108203
rect 90180 -109117 90256 -108203
rect 90788 -109117 90864 -108203
rect 91396 -109117 91472 -108203
rect 92004 -109117 92080 -108203
rect 92612 -109117 92688 -108203
rect 93220 -109117 93296 -108203
rect 93828 -109117 93904 -108203
rect 94436 -109117 94512 -108203
rect 95044 -109117 95120 -108203
rect 95652 -109117 95728 -108203
rect 96260 -109117 96336 -108203
rect 96868 -109117 96944 -108203
rect 97476 -109117 97552 -108203
rect 98084 -109117 98160 -108203
rect 98692 -109117 98768 -108203
rect 99300 -109117 99376 -108203
rect 99908 -109117 99984 -108203
rect 100516 -109117 100592 -108203
rect 101124 -109117 101200 -108203
rect 101732 -109117 101808 -108203
rect 102340 -109117 102416 -108203
rect 102948 -109117 103024 -108203
rect 103556 -109117 103632 -108203
rect 104164 -109117 104240 -108203
rect 104772 -109117 104848 -108203
rect 105380 -109117 105456 -108203
rect 105988 -109117 106064 -108203
rect 106596 -109117 106672 -108203
rect 107204 -109117 107280 -108203
rect 107812 -109117 107888 -108203
rect 108420 -109117 108496 -108203
rect 109028 -109117 109104 -108203
rect 109636 -109117 109712 -108203
rect 110244 -109117 110320 -108203
rect 110852 -109117 110928 -108203
rect 111460 -109117 111536 -108203
rect 112068 -109117 112144 -108203
rect 112676 -109117 112752 -108203
rect 113284 -109117 113360 -108203
rect 114884 -109117 114960 -108203
rect 115492 -109117 115568 -108203
rect 116100 -109117 116176 -108203
rect 116708 -109117 116784 -108203
rect 117316 -109117 117392 -108203
rect 117924 -109117 118000 -108203
rect 118532 -109117 118608 -108203
rect 119140 -109117 119216 -108203
rect 119748 -109117 119824 -108203
rect 120356 -109117 120432 -108203
rect 120964 -109117 121040 -108203
rect 121572 -109117 121648 -108203
rect 122180 -109117 122256 -108203
rect 122788 -109117 122864 -108203
rect 123396 -109117 123472 -108203
rect 124004 -109117 124080 -108203
rect 124612 -109117 124688 -108203
rect 125220 -109117 125296 -108203
rect 125828 -109117 125904 -108203
rect 126436 -109117 126512 -108203
rect 127044 -109117 127120 -108203
rect 127652 -109117 127728 -108203
rect 128260 -109117 128336 -108203
rect 128868 -109117 128944 -108203
rect 129476 -109117 129552 -108203
rect 130084 -109117 130160 -108203
rect 130692 -109117 130768 -108203
rect 131300 -109117 131376 -108203
rect 131908 -109117 131984 -108203
rect 132516 -109117 132592 -108203
rect 133124 -109117 133200 -108203
rect 133732 -109117 133808 -108203
rect 134340 -109117 134416 -108203
rect 134948 -109117 135024 -108203
rect 135556 -109117 135632 -108203
rect 136164 -109117 136240 -108203
rect 136772 -109117 136848 -108203
rect 137380 -109117 137456 -108203
rect 137988 -109117 138064 -108203
rect 138596 -109117 138672 -108203
rect 139204 -109117 139280 -108203
rect 139812 -109117 139888 -108203
rect 140420 -109117 140496 -108203
rect 141028 -109117 141104 -108203
rect 141636 -109117 141712 -108203
rect 142244 -109117 142320 -108203
rect 142852 -109117 142928 -108203
rect 143460 -109117 143536 -108203
rect 144068 -109117 144144 -108203
rect 144676 -109117 144752 -108203
rect 145284 -109117 145360 -108203
rect 146884 -109117 146960 -108203
rect 147492 -109117 147568 -108203
rect 148100 -109117 148176 -108203
rect 148708 -109117 148784 -108203
rect 149316 -109117 149392 -108203
rect 149924 -109117 150000 -108203
rect 150532 -109117 150608 -108203
rect 151140 -109117 151216 -108203
rect 151748 -109117 151824 -108203
rect 152356 -109117 152432 -108203
rect 152964 -109117 153040 -108203
rect 153572 -109117 153648 -108203
rect 154180 -109117 154256 -108203
rect 154788 -109117 154864 -108203
rect 155396 -109117 155472 -108203
rect 156004 -109117 156080 -108203
rect 156612 -109117 156688 -108203
rect 157220 -109117 157296 -108203
rect 157828 -109117 157904 -108203
rect 158436 -109117 158512 -108203
rect 159044 -109117 159120 -108203
rect 159652 -109117 159728 -108203
rect 160260 -109117 160336 -108203
rect 160868 -109117 160944 -108203
rect 161476 -109117 161552 -108203
rect 162084 -109117 162160 -108203
rect 162692 -109117 162768 -108203
rect 163300 -109117 163376 -108203
rect 163908 -109117 163984 -108203
rect 164516 -109117 164592 -108203
rect 165124 -109117 165200 -108203
rect 165732 -109117 165808 -108203
rect 166340 -109117 166416 -108203
rect 166948 -109117 167024 -108203
rect 167556 -109117 167632 -108203
rect 168164 -109117 168240 -108203
rect 168772 -109117 168848 -108203
rect 169380 -109117 169456 -108203
rect 169988 -109117 170064 -108203
rect 170596 -109117 170672 -108203
rect 171204 -109117 171280 -108203
rect 171812 -109117 171888 -108203
rect 172420 -109117 172496 -108203
rect 173028 -109117 173104 -108203
rect 173636 -109117 173712 -108203
rect 174244 -109117 174320 -108203
rect 174852 -109117 174928 -108203
rect 175460 -109117 175536 -108203
rect 176068 -109117 176144 -108203
rect 176676 -109117 176752 -108203
rect 177284 -109117 177360 -108203
rect -77274 -129121 -77040 -109119
rect -45274 -129121 -45040 -109119
rect -13274 -129121 -13040 -109119
rect 18726 -129121 18960 -109119
rect 50726 -129121 50960 -109119
rect 82726 -129121 82960 -109119
rect 114726 -129121 114960 -109119
rect 146726 -129121 146960 -109119
rect -108812 -130035 -108736 -129121
rect -108204 -130035 -108128 -129121
rect -107596 -130035 -107520 -129121
rect -106988 -130035 -106912 -129121
rect -106380 -130035 -106304 -129121
rect -105772 -130035 -105696 -129121
rect -105164 -130035 -105088 -129121
rect -104556 -130035 -104480 -129121
rect -103948 -130035 -103872 -129121
rect -103340 -130035 -103264 -129121
rect -102732 -130035 -102656 -129121
rect -102124 -130035 -102048 -129121
rect -101516 -130035 -101440 -129121
rect -100908 -130035 -100832 -129121
rect -100300 -130035 -100224 -129121
rect -99692 -130035 -99616 -129121
rect -99084 -130035 -99008 -129121
rect -98476 -130035 -98400 -129121
rect -97868 -130035 -97792 -129121
rect -97260 -130035 -97184 -129121
rect -96652 -130035 -96576 -129121
rect -96044 -130035 -95968 -129121
rect -95436 -130035 -95360 -129121
rect -94828 -130035 -94752 -129121
rect -94220 -130035 -94144 -129121
rect -93612 -130035 -93536 -129121
rect -93004 -130035 -92928 -129121
rect -92396 -130035 -92320 -129121
rect -91788 -130035 -91712 -129121
rect -91180 -130035 -91104 -129121
rect -90572 -130035 -90496 -129121
rect -89964 -130035 -89888 -129121
rect -89356 -130035 -89280 -129121
rect -88748 -130035 -88672 -129121
rect -88140 -130035 -88064 -129121
rect -87532 -130035 -87456 -129121
rect -86924 -130035 -86848 -129121
rect -86316 -130035 -86240 -129121
rect -85708 -130035 -85632 -129121
rect -85100 -130035 -85024 -129121
rect -84492 -130035 -84416 -129121
rect -83884 -130035 -83808 -129121
rect -83276 -130035 -83200 -129121
rect -82668 -130035 -82592 -129121
rect -82060 -130035 -81984 -129121
rect -81452 -130035 -81376 -129121
rect -80844 -130035 -80768 -129121
rect -80236 -130035 -80160 -129121
rect -79628 -130035 -79552 -129121
rect -79020 -130035 -78944 -129121
rect -76812 -130035 -76736 -129121
rect -76204 -130035 -76128 -129121
rect -75596 -130035 -75520 -129121
rect -74988 -130035 -74912 -129121
rect -74380 -130035 -74304 -129121
rect -73772 -130035 -73696 -129121
rect -73164 -130035 -73088 -129121
rect -72556 -130035 -72480 -129121
rect -71948 -130035 -71872 -129121
rect -71340 -130035 -71264 -129121
rect -70732 -130035 -70656 -129121
rect -70124 -130035 -70048 -129121
rect -69516 -130035 -69440 -129121
rect -68908 -130035 -68832 -129121
rect -68300 -130035 -68224 -129121
rect -67692 -130035 -67616 -129121
rect -67084 -130035 -67008 -129121
rect -66476 -130035 -66400 -129121
rect -65868 -130035 -65792 -129121
rect -65260 -130035 -65184 -129121
rect -64652 -130035 -64576 -129121
rect -64044 -130035 -63968 -129121
rect -63436 -130035 -63360 -129121
rect -62828 -130035 -62752 -129121
rect -62220 -130035 -62144 -129121
rect -61612 -130035 -61536 -129121
rect -61004 -130035 -60928 -129121
rect -60396 -130035 -60320 -129121
rect -59788 -130035 -59712 -129121
rect -59180 -130035 -59104 -129121
rect -58572 -130035 -58496 -129121
rect -57964 -130035 -57888 -129121
rect -57356 -130035 -57280 -129121
rect -56748 -130035 -56672 -129121
rect -56140 -130035 -56064 -129121
rect -55532 -130035 -55456 -129121
rect -54924 -130035 -54848 -129121
rect -54316 -130035 -54240 -129121
rect -53708 -130035 -53632 -129121
rect -53100 -130035 -53024 -129121
rect -52492 -130035 -52416 -129121
rect -51884 -130035 -51808 -129121
rect -51276 -130035 -51200 -129121
rect -50668 -130035 -50592 -129121
rect -50060 -130035 -49984 -129121
rect -49452 -130035 -49376 -129121
rect -48844 -130035 -48768 -129121
rect -48236 -130035 -48160 -129121
rect -47628 -130035 -47552 -129121
rect -47020 -130035 -46944 -129121
rect -44812 -130035 -44736 -129121
rect -44204 -130035 -44128 -129121
rect -43596 -130035 -43520 -129121
rect -42988 -130035 -42912 -129121
rect -42380 -130035 -42304 -129121
rect -41772 -130035 -41696 -129121
rect -41164 -130035 -41088 -129121
rect -40556 -130035 -40480 -129121
rect -39948 -130035 -39872 -129121
rect -39340 -130035 -39264 -129121
rect -38732 -130035 -38656 -129121
rect -38124 -130035 -38048 -129121
rect -37516 -130035 -37440 -129121
rect -36908 -130035 -36832 -129121
rect -36300 -130035 -36224 -129121
rect -35692 -130035 -35616 -129121
rect -35084 -130035 -35008 -129121
rect -34476 -130035 -34400 -129121
rect -33868 -130035 -33792 -129121
rect -33260 -130035 -33184 -129121
rect -32652 -130035 -32576 -129121
rect -32044 -130035 -31968 -129121
rect -31436 -130035 -31360 -129121
rect -30828 -130035 -30752 -129121
rect -30220 -130035 -30144 -129121
rect -29612 -130035 -29536 -129121
rect -29004 -130035 -28928 -129121
rect -28396 -130035 -28320 -129121
rect -27788 -130035 -27712 -129121
rect -27180 -130035 -27104 -129121
rect -26572 -130035 -26496 -129121
rect -25964 -130035 -25888 -129121
rect -25356 -130035 -25280 -129121
rect -24748 -130035 -24672 -129121
rect -24140 -130035 -24064 -129121
rect -23532 -130035 -23456 -129121
rect -22924 -130035 -22848 -129121
rect -22316 -130035 -22240 -129121
rect -21708 -130035 -21632 -129121
rect -21100 -130035 -21024 -129121
rect -20492 -130035 -20416 -129121
rect -19884 -130035 -19808 -129121
rect -19276 -130035 -19200 -129121
rect -18668 -130035 -18592 -129121
rect -18060 -130035 -17984 -129121
rect -17452 -130035 -17376 -129121
rect -16844 -130035 -16768 -129121
rect -16236 -130035 -16160 -129121
rect -15628 -130035 -15552 -129121
rect -15020 -130035 -14944 -129121
rect -12812 -130035 -12736 -129121
rect -12204 -130035 -12128 -129121
rect -11596 -130035 -11520 -129121
rect -10988 -130035 -10912 -129121
rect -10380 -130035 -10304 -129121
rect -9772 -130035 -9696 -129121
rect -9164 -130035 -9088 -129121
rect -8556 -130035 -8480 -129121
rect -7948 -130035 -7872 -129121
rect -7340 -130035 -7264 -129121
rect -6732 -130035 -6656 -129121
rect -6124 -130035 -6048 -129121
rect -5516 -130035 -5440 -129121
rect -4908 -130035 -4832 -129121
rect -4300 -130035 -4224 -129121
rect -3692 -130035 -3616 -129121
rect -3084 -130035 -3008 -129121
rect -2476 -130035 -2400 -129121
rect -1868 -130035 -1792 -129121
rect -1260 -130035 -1184 -129121
rect -652 -130035 -576 -129121
rect -44 -130035 32 -129121
rect 564 -130035 640 -129121
rect 1172 -130035 1248 -129121
rect 1780 -130035 1856 -129121
rect 2388 -130035 2464 -129121
rect 2996 -130035 3072 -129121
rect 3604 -130035 3680 -129121
rect 4212 -130035 4288 -129121
rect 4820 -130035 4896 -129121
rect 5428 -130035 5504 -129121
rect 6036 -130035 6112 -129121
rect 6644 -130035 6720 -129121
rect 7252 -130035 7328 -129121
rect 7860 -130035 7936 -129121
rect 8468 -130035 8544 -129121
rect 9076 -130035 9152 -129121
rect 9684 -130035 9760 -129121
rect 10292 -130035 10368 -129121
rect 10900 -130035 10976 -129121
rect 11508 -130035 11584 -129121
rect 12116 -130035 12192 -129121
rect 12724 -130035 12800 -129121
rect 13332 -130035 13408 -129121
rect 13940 -130035 14016 -129121
rect 14548 -130035 14624 -129121
rect 15156 -130035 15232 -129121
rect 15764 -130035 15840 -129121
rect 16372 -130035 16448 -129121
rect 16980 -130035 17056 -129121
rect 19188 -130035 19264 -129121
rect 19796 -130035 19872 -129121
rect 20404 -130035 20480 -129121
rect 21012 -130035 21088 -129121
rect 21620 -130035 21696 -129121
rect 22228 -130035 22304 -129121
rect 22836 -130035 22912 -129121
rect 23444 -130035 23520 -129121
rect 24052 -130035 24128 -129121
rect 24660 -130035 24736 -129121
rect 25268 -130035 25344 -129121
rect 25876 -130035 25952 -129121
rect 26484 -130035 26560 -129121
rect 27092 -130035 27168 -129121
rect 27700 -130035 27776 -129121
rect 28308 -130035 28384 -129121
rect 28916 -130035 28992 -129121
rect 29524 -130035 29600 -129121
rect 30132 -130035 30208 -129121
rect 30740 -130035 30816 -129121
rect 31348 -130035 31424 -129121
rect 31956 -130035 32032 -129121
rect 32564 -130035 32640 -129121
rect 33172 -130035 33248 -129121
rect 33780 -130035 33856 -129121
rect 34388 -130035 34464 -129121
rect 34996 -130035 35072 -129121
rect 35604 -130035 35680 -129121
rect 36212 -130035 36288 -129121
rect 36820 -130035 36896 -129121
rect 37428 -130035 37504 -129121
rect 38036 -130035 38112 -129121
rect 38644 -130035 38720 -129121
rect 39252 -130035 39328 -129121
rect 39860 -130035 39936 -129121
rect 40468 -130035 40544 -129121
rect 41076 -130035 41152 -129121
rect 41684 -130035 41760 -129121
rect 42292 -130035 42368 -129121
rect 42900 -130035 42976 -129121
rect 43508 -130035 43584 -129121
rect 44116 -130035 44192 -129121
rect 44724 -130035 44800 -129121
rect 45332 -130035 45408 -129121
rect 45940 -130035 46016 -129121
rect 46548 -130035 46624 -129121
rect 47156 -130035 47232 -129121
rect 47764 -130035 47840 -129121
rect 48372 -130035 48448 -129121
rect 48980 -130035 49056 -129121
rect 51188 -130035 51264 -129121
rect 51796 -130035 51872 -129121
rect 52404 -130035 52480 -129121
rect 53012 -130035 53088 -129121
rect 53620 -130035 53696 -129121
rect 54228 -130035 54304 -129121
rect 54836 -130035 54912 -129121
rect 55444 -130035 55520 -129121
rect 56052 -130035 56128 -129121
rect 56660 -130035 56736 -129121
rect 57268 -130035 57344 -129121
rect 57876 -130035 57952 -129121
rect 58484 -130035 58560 -129121
rect 59092 -130035 59168 -129121
rect 59700 -130035 59776 -129121
rect 60308 -130035 60384 -129121
rect 60916 -130035 60992 -129121
rect 61524 -130035 61600 -129121
rect 62132 -130035 62208 -129121
rect 62740 -130035 62816 -129121
rect 63348 -130035 63424 -129121
rect 63956 -130035 64032 -129121
rect 64564 -130035 64640 -129121
rect 65172 -130035 65248 -129121
rect 65780 -130035 65856 -129121
rect 66388 -130035 66464 -129121
rect 66996 -130035 67072 -129121
rect 67604 -130035 67680 -129121
rect 68212 -130035 68288 -129121
rect 68820 -130035 68896 -129121
rect 69428 -130035 69504 -129121
rect 70036 -130035 70112 -129121
rect 70644 -130035 70720 -129121
rect 71252 -130035 71328 -129121
rect 71860 -130035 71936 -129121
rect 72468 -130035 72544 -129121
rect 73076 -130035 73152 -129121
rect 73684 -130035 73760 -129121
rect 74292 -130035 74368 -129121
rect 74900 -130035 74976 -129121
rect 75508 -130035 75584 -129121
rect 76116 -130035 76192 -129121
rect 76724 -130035 76800 -129121
rect 77332 -130035 77408 -129121
rect 77940 -130035 78016 -129121
rect 78548 -130035 78624 -129121
rect 79156 -130035 79232 -129121
rect 79764 -130035 79840 -129121
rect 80372 -130035 80448 -129121
rect 80980 -130035 81056 -129121
rect 83188 -130035 83264 -129121
rect 83796 -130035 83872 -129121
rect 84404 -130035 84480 -129121
rect 85012 -130035 85088 -129121
rect 85620 -130035 85696 -129121
rect 86228 -130035 86304 -129121
rect 86836 -130035 86912 -129121
rect 87444 -130035 87520 -129121
rect 88052 -130035 88128 -129121
rect 88660 -130035 88736 -129121
rect 89268 -130035 89344 -129121
rect 89876 -130035 89952 -129121
rect 90484 -130035 90560 -129121
rect 91092 -130035 91168 -129121
rect 91700 -130035 91776 -129121
rect 92308 -130035 92384 -129121
rect 92916 -130035 92992 -129121
rect 93524 -130035 93600 -129121
rect 94132 -130035 94208 -129121
rect 94740 -130035 94816 -129121
rect 95348 -130035 95424 -129121
rect 95956 -130035 96032 -129121
rect 96564 -130035 96640 -129121
rect 97172 -130035 97248 -129121
rect 97780 -130035 97856 -129121
rect 98388 -130035 98464 -129121
rect 98996 -130035 99072 -129121
rect 99604 -130035 99680 -129121
rect 100212 -130035 100288 -129121
rect 100820 -130035 100896 -129121
rect 101428 -130035 101504 -129121
rect 102036 -130035 102112 -129121
rect 102644 -130035 102720 -129121
rect 103252 -130035 103328 -129121
rect 103860 -130035 103936 -129121
rect 104468 -130035 104544 -129121
rect 105076 -130035 105152 -129121
rect 105684 -130035 105760 -129121
rect 106292 -130035 106368 -129121
rect 106900 -130035 106976 -129121
rect 107508 -130035 107584 -129121
rect 108116 -130035 108192 -129121
rect 108724 -130035 108800 -129121
rect 109332 -130035 109408 -129121
rect 109940 -130035 110016 -129121
rect 110548 -130035 110624 -129121
rect 111156 -130035 111232 -129121
rect 111764 -130035 111840 -129121
rect 112372 -130035 112448 -129121
rect 112980 -130035 113056 -129121
rect 115188 -130035 115264 -129121
rect 115796 -130035 115872 -129121
rect 116404 -130035 116480 -129121
rect 117012 -130035 117088 -129121
rect 117620 -130035 117696 -129121
rect 118228 -130035 118304 -129121
rect 118836 -130035 118912 -129121
rect 119444 -130035 119520 -129121
rect 120052 -130035 120128 -129121
rect 120660 -130035 120736 -129121
rect 121268 -130035 121344 -129121
rect 121876 -130035 121952 -129121
rect 122484 -130035 122560 -129121
rect 123092 -130035 123168 -129121
rect 123700 -130035 123776 -129121
rect 124308 -130035 124384 -129121
rect 124916 -130035 124992 -129121
rect 125524 -130035 125600 -129121
rect 126132 -130035 126208 -129121
rect 126740 -130035 126816 -129121
rect 127348 -130035 127424 -129121
rect 127956 -130035 128032 -129121
rect 128564 -130035 128640 -129121
rect 129172 -130035 129248 -129121
rect 129780 -130035 129856 -129121
rect 130388 -130035 130464 -129121
rect 130996 -130035 131072 -129121
rect 131604 -130035 131680 -129121
rect 132212 -130035 132288 -129121
rect 132820 -130035 132896 -129121
rect 133428 -130035 133504 -129121
rect 134036 -130035 134112 -129121
rect 134644 -130035 134720 -129121
rect 135252 -130035 135328 -129121
rect 135860 -130035 135936 -129121
rect 136468 -130035 136544 -129121
rect 137076 -130035 137152 -129121
rect 137684 -130035 137760 -129121
rect 138292 -130035 138368 -129121
rect 138900 -130035 138976 -129121
rect 139508 -130035 139584 -129121
rect 140116 -130035 140192 -129121
rect 140724 -130035 140800 -129121
rect 141332 -130035 141408 -129121
rect 141940 -130035 142016 -129121
rect 142548 -130035 142624 -129121
rect 143156 -130035 143232 -129121
rect 143764 -130035 143840 -129121
rect 144372 -130035 144448 -129121
rect 144980 -130035 145056 -129121
rect 147188 -130035 147264 -129121
rect 147796 -130035 147872 -129121
rect 148404 -130035 148480 -129121
rect 149012 -130035 149088 -129121
rect 149620 -130035 149696 -129121
rect 150228 -130035 150304 -129121
rect 150836 -130035 150912 -129121
rect 151444 -130035 151520 -129121
rect 152052 -130035 152128 -129121
rect 152660 -130035 152736 -129121
rect 153268 -130035 153344 -129121
rect 153876 -130035 153952 -129121
rect 154484 -130035 154560 -129121
rect 155092 -130035 155168 -129121
rect 155700 -130035 155776 -129121
rect 156308 -130035 156384 -129121
rect 156916 -130035 156992 -129121
rect 157524 -130035 157600 -129121
rect 158132 -130035 158208 -129121
rect 158740 -130035 158816 -129121
rect 159348 -130035 159424 -129121
rect 159956 -130035 160032 -129121
rect 160564 -130035 160640 -129121
rect 161172 -130035 161248 -129121
rect 161780 -130035 161856 -129121
rect 162388 -130035 162464 -129121
rect 162996 -130035 163072 -129121
rect 163604 -130035 163680 -129121
rect 164212 -130035 164288 -129121
rect 164820 -130035 164896 -129121
rect 165428 -130035 165504 -129121
rect 166036 -130035 166112 -129121
rect 166644 -130035 166720 -129121
rect 167252 -130035 167328 -129121
rect 167860 -130035 167936 -129121
rect 168468 -130035 168544 -129121
rect 169076 -130035 169152 -129121
rect 169684 -130035 169760 -129121
rect 170292 -130035 170368 -129121
rect 170900 -130035 170976 -129121
rect 171508 -130035 171584 -129121
rect 172116 -130035 172192 -129121
rect 172724 -130035 172800 -129121
rect 173332 -130035 173408 -129121
rect 173940 -130035 174016 -129121
rect 174548 -130035 174624 -129121
rect 175156 -130035 175232 -129121
rect 175764 -130035 175840 -129121
rect 176372 -130035 176448 -129121
rect 176980 -130035 177056 -129121
rect 177664 -130035 178308 -104602
rect -108812 -130602 178308 -130035
rect -108812 -131251 177664 -130602
rect -108812 -131295 -13354 -131251
rect -13310 -131295 -13254 -131251
rect -13210 -131295 -13154 -131251
rect -13110 -131295 -13054 -131251
rect -13010 -131295 -12954 -131251
rect -12910 -131295 -12854 -131251
rect -12810 -131295 -12754 -131251
rect -12710 -131295 -12654 -131251
rect -12610 -131295 -12554 -131251
rect -12510 -131295 -12454 -131251
rect -12410 -131295 -12354 -131251
rect -12310 -131295 -12254 -131251
rect -12210 -131295 -12154 -131251
rect -12110 -131295 -12054 -131251
rect -12010 -131295 -11954 -131251
rect -11910 -131295 -11854 -131251
rect -11810 -131295 -11354 -131251
rect -11310 -131295 -11254 -131251
rect -11210 -131295 -11154 -131251
rect -11110 -131295 -11054 -131251
rect -11010 -131295 -10954 -131251
rect -10910 -131295 -10854 -131251
rect -10810 -131295 -10754 -131251
rect -10710 -131295 -10654 -131251
rect -10610 -131295 -10554 -131251
rect -10510 -131295 -10454 -131251
rect -10410 -131295 -10354 -131251
rect -10310 -131295 -10254 -131251
rect -10210 -131295 -10154 -131251
rect -10110 -131295 -10054 -131251
rect -10010 -131295 -9954 -131251
rect -9910 -131295 -9854 -131251
rect -9810 -131295 -9354 -131251
rect -9310 -131295 -9254 -131251
rect -9210 -131295 -9154 -131251
rect -9110 -131295 -9054 -131251
rect -9010 -131295 -8954 -131251
rect -8910 -131295 -8854 -131251
rect -8810 -131295 -8754 -131251
rect -8710 -131295 -8654 -131251
rect -8610 -131295 -8554 -131251
rect -8510 -131295 -8454 -131251
rect -8410 -131295 -8354 -131251
rect -8310 -131295 -8254 -131251
rect -8210 -131295 -8154 -131251
rect -8110 -131295 -8054 -131251
rect -8010 -131295 -7954 -131251
rect -7910 -131295 -7854 -131251
rect -7810 -131295 -7354 -131251
rect -7310 -131295 -7254 -131251
rect -7210 -131295 -7154 -131251
rect -7110 -131295 -7054 -131251
rect -7010 -131295 -6954 -131251
rect -6910 -131295 -6854 -131251
rect -6810 -131295 -6754 -131251
rect -6710 -131295 -6654 -131251
rect -6610 -131295 -6554 -131251
rect -6510 -131295 -6454 -131251
rect -6410 -131295 -6354 -131251
rect -6310 -131295 -6254 -131251
rect -6210 -131295 -6154 -131251
rect -6110 -131295 -6054 -131251
rect -6010 -131295 -5954 -131251
rect -5910 -131295 -5854 -131251
rect -5810 -131295 177664 -131251
rect -108812 -131351 177664 -131295
rect -108812 -131395 -13354 -131351
rect -13310 -131395 -13254 -131351
rect -13210 -131395 -13154 -131351
rect -13110 -131395 -13054 -131351
rect -13010 -131395 -12954 -131351
rect -12910 -131395 -12854 -131351
rect -12810 -131395 -12754 -131351
rect -12710 -131395 -12654 -131351
rect -12610 -131395 -12554 -131351
rect -12510 -131395 -12454 -131351
rect -12410 -131395 -12354 -131351
rect -12310 -131395 -12254 -131351
rect -12210 -131395 -12154 -131351
rect -12110 -131395 -12054 -131351
rect -12010 -131395 -11954 -131351
rect -11910 -131395 -11854 -131351
rect -11810 -131395 -11354 -131351
rect -11310 -131395 -11254 -131351
rect -11210 -131395 -11154 -131351
rect -11110 -131395 -11054 -131351
rect -11010 -131395 -10954 -131351
rect -10910 -131395 -10854 -131351
rect -10810 -131395 -10754 -131351
rect -10710 -131395 -10654 -131351
rect -10610 -131395 -10554 -131351
rect -10510 -131395 -10454 -131351
rect -10410 -131395 -10354 -131351
rect -10310 -131395 -10254 -131351
rect -10210 -131395 -10154 -131351
rect -10110 -131395 -10054 -131351
rect -10010 -131395 -9954 -131351
rect -9910 -131395 -9854 -131351
rect -9810 -131395 -9354 -131351
rect -9310 -131395 -9254 -131351
rect -9210 -131395 -9154 -131351
rect -9110 -131395 -9054 -131351
rect -9010 -131395 -8954 -131351
rect -8910 -131395 -8854 -131351
rect -8810 -131395 -8754 -131351
rect -8710 -131395 -8654 -131351
rect -8610 -131395 -8554 -131351
rect -8510 -131395 -8454 -131351
rect -8410 -131395 -8354 -131351
rect -8310 -131395 -8254 -131351
rect -8210 -131395 -8154 -131351
rect -8110 -131395 -8054 -131351
rect -8010 -131395 -7954 -131351
rect -7910 -131395 -7854 -131351
rect -7810 -131395 -7354 -131351
rect -7310 -131395 -7254 -131351
rect -7210 -131395 -7154 -131351
rect -7110 -131395 -7054 -131351
rect -7010 -131395 -6954 -131351
rect -6910 -131395 -6854 -131351
rect -6810 -131395 -6754 -131351
rect -6710 -131395 -6654 -131351
rect -6610 -131395 -6554 -131351
rect -6510 -131395 -6454 -131351
rect -6410 -131395 -6354 -131351
rect -6310 -131395 -6254 -131351
rect -6210 -131395 -6154 -131351
rect -6110 -131395 -6054 -131351
rect -6010 -131395 -5954 -131351
rect -5910 -131395 -5854 -131351
rect -5810 -131385 177664 -131351
rect -5810 -131395 37387 -131385
rect -108812 -131429 37387 -131395
rect 37431 -131429 37487 -131385
rect 37531 -131429 37587 -131385
rect 37631 -131429 37687 -131385
rect 37731 -131429 37787 -131385
rect 37831 -131429 37887 -131385
rect 37931 -131429 37987 -131385
rect 38031 -131429 38087 -131385
rect 38131 -131429 38187 -131385
rect 38231 -131429 38287 -131385
rect 38331 -131429 38387 -131385
rect 38431 -131429 38487 -131385
rect 38531 -131429 38587 -131385
rect 38631 -131429 38687 -131385
rect 38731 -131429 38787 -131385
rect 38831 -131429 38887 -131385
rect 38931 -131429 39387 -131385
rect 39431 -131429 39487 -131385
rect 39531 -131429 39587 -131385
rect 39631 -131429 39687 -131385
rect 39731 -131429 39787 -131385
rect 39831 -131429 39887 -131385
rect 39931 -131429 39987 -131385
rect 40031 -131429 40087 -131385
rect 40131 -131429 40187 -131385
rect 40231 -131429 40287 -131385
rect 40331 -131429 40387 -131385
rect 40431 -131429 40487 -131385
rect 40531 -131429 40587 -131385
rect 40631 -131429 40687 -131385
rect 40731 -131429 40787 -131385
rect 40831 -131429 40887 -131385
rect 40931 -131429 41387 -131385
rect 41431 -131429 41487 -131385
rect 41531 -131429 41587 -131385
rect 41631 -131429 41687 -131385
rect 41731 -131429 41787 -131385
rect 41831 -131429 41887 -131385
rect 41931 -131429 41987 -131385
rect 42031 -131429 42087 -131385
rect 42131 -131429 42187 -131385
rect 42231 -131429 42287 -131385
rect 42331 -131429 42387 -131385
rect 42431 -131429 42487 -131385
rect 42531 -131429 42587 -131385
rect 42631 -131429 42687 -131385
rect 42731 -131429 42787 -131385
rect 42831 -131429 42887 -131385
rect 42931 -131429 43387 -131385
rect 43431 -131429 43487 -131385
rect 43531 -131429 43587 -131385
rect 43631 -131429 43687 -131385
rect 43731 -131429 43787 -131385
rect 43831 -131429 43887 -131385
rect 43931 -131429 43987 -131385
rect 44031 -131429 44087 -131385
rect 44131 -131429 44187 -131385
rect 44231 -131429 44287 -131385
rect 44331 -131429 44387 -131385
rect 44431 -131429 44487 -131385
rect 44531 -131429 44587 -131385
rect 44631 -131429 44687 -131385
rect 44731 -131429 44787 -131385
rect 44831 -131429 44887 -131385
rect 44931 -131429 177664 -131385
rect -108812 -131451 177664 -131429
rect -108812 -131495 -13354 -131451
rect -13310 -131495 -13254 -131451
rect -13210 -131495 -13154 -131451
rect -13110 -131495 -13054 -131451
rect -13010 -131495 -12954 -131451
rect -12910 -131495 -12854 -131451
rect -12810 -131495 -12754 -131451
rect -12710 -131495 -12654 -131451
rect -12610 -131495 -12554 -131451
rect -12510 -131495 -12454 -131451
rect -12410 -131495 -12354 -131451
rect -12310 -131495 -12254 -131451
rect -12210 -131495 -12154 -131451
rect -12110 -131495 -12054 -131451
rect -12010 -131495 -11954 -131451
rect -11910 -131495 -11854 -131451
rect -11810 -131495 -11354 -131451
rect -11310 -131495 -11254 -131451
rect -11210 -131495 -11154 -131451
rect -11110 -131495 -11054 -131451
rect -11010 -131495 -10954 -131451
rect -10910 -131495 -10854 -131451
rect -10810 -131495 -10754 -131451
rect -10710 -131495 -10654 -131451
rect -10610 -131495 -10554 -131451
rect -10510 -131495 -10454 -131451
rect -10410 -131495 -10354 -131451
rect -10310 -131495 -10254 -131451
rect -10210 -131495 -10154 -131451
rect -10110 -131495 -10054 -131451
rect -10010 -131495 -9954 -131451
rect -9910 -131495 -9854 -131451
rect -9810 -131495 -9354 -131451
rect -9310 -131495 -9254 -131451
rect -9210 -131495 -9154 -131451
rect -9110 -131495 -9054 -131451
rect -9010 -131495 -8954 -131451
rect -8910 -131495 -8854 -131451
rect -8810 -131495 -8754 -131451
rect -8710 -131495 -8654 -131451
rect -8610 -131495 -8554 -131451
rect -8510 -131495 -8454 -131451
rect -8410 -131495 -8354 -131451
rect -8310 -131495 -8254 -131451
rect -8210 -131495 -8154 -131451
rect -8110 -131495 -8054 -131451
rect -8010 -131495 -7954 -131451
rect -7910 -131495 -7854 -131451
rect -7810 -131495 -7354 -131451
rect -7310 -131495 -7254 -131451
rect -7210 -131495 -7154 -131451
rect -7110 -131495 -7054 -131451
rect -7010 -131495 -6954 -131451
rect -6910 -131495 -6854 -131451
rect -6810 -131495 -6754 -131451
rect -6710 -131495 -6654 -131451
rect -6610 -131495 -6554 -131451
rect -6510 -131495 -6454 -131451
rect -6410 -131495 -6354 -131451
rect -6310 -131495 -6254 -131451
rect -6210 -131495 -6154 -131451
rect -6110 -131495 -6054 -131451
rect -6010 -131495 -5954 -131451
rect -5910 -131495 -5854 -131451
rect -5810 -131485 177664 -131451
rect -5810 -131495 37387 -131485
rect -108812 -131529 37387 -131495
rect 37431 -131529 37487 -131485
rect 37531 -131529 37587 -131485
rect 37631 -131529 37687 -131485
rect 37731 -131529 37787 -131485
rect 37831 -131529 37887 -131485
rect 37931 -131529 37987 -131485
rect 38031 -131529 38087 -131485
rect 38131 -131529 38187 -131485
rect 38231 -131529 38287 -131485
rect 38331 -131529 38387 -131485
rect 38431 -131529 38487 -131485
rect 38531 -131529 38587 -131485
rect 38631 -131529 38687 -131485
rect 38731 -131529 38787 -131485
rect 38831 -131529 38887 -131485
rect 38931 -131529 39387 -131485
rect 39431 -131529 39487 -131485
rect 39531 -131529 39587 -131485
rect 39631 -131529 39687 -131485
rect 39731 -131529 39787 -131485
rect 39831 -131529 39887 -131485
rect 39931 -131529 39987 -131485
rect 40031 -131529 40087 -131485
rect 40131 -131529 40187 -131485
rect 40231 -131529 40287 -131485
rect 40331 -131529 40387 -131485
rect 40431 -131529 40487 -131485
rect 40531 -131529 40587 -131485
rect 40631 -131529 40687 -131485
rect 40731 -131529 40787 -131485
rect 40831 -131529 40887 -131485
rect 40931 -131529 41387 -131485
rect 41431 -131529 41487 -131485
rect 41531 -131529 41587 -131485
rect 41631 -131529 41687 -131485
rect 41731 -131529 41787 -131485
rect 41831 -131529 41887 -131485
rect 41931 -131529 41987 -131485
rect 42031 -131529 42087 -131485
rect 42131 -131529 42187 -131485
rect 42231 -131529 42287 -131485
rect 42331 -131529 42387 -131485
rect 42431 -131529 42487 -131485
rect 42531 -131529 42587 -131485
rect 42631 -131529 42687 -131485
rect 42731 -131529 42787 -131485
rect 42831 -131529 42887 -131485
rect 42931 -131529 43387 -131485
rect 43431 -131529 43487 -131485
rect 43531 -131529 43587 -131485
rect 43631 -131529 43687 -131485
rect 43731 -131529 43787 -131485
rect 43831 -131529 43887 -131485
rect 43931 -131529 43987 -131485
rect 44031 -131529 44087 -131485
rect 44131 -131529 44187 -131485
rect 44231 -131529 44287 -131485
rect 44331 -131529 44387 -131485
rect 44431 -131529 44487 -131485
rect 44531 -131529 44587 -131485
rect 44631 -131529 44687 -131485
rect 44731 -131529 44787 -131485
rect 44831 -131529 44887 -131485
rect 44931 -131529 177664 -131485
rect -108812 -131551 177664 -131529
rect -108812 -131595 -13354 -131551
rect -13310 -131595 -13254 -131551
rect -13210 -131595 -13154 -131551
rect -13110 -131595 -13054 -131551
rect -13010 -131595 -12954 -131551
rect -12910 -131595 -12854 -131551
rect -12810 -131595 -12754 -131551
rect -12710 -131595 -12654 -131551
rect -12610 -131595 -12554 -131551
rect -12510 -131595 -12454 -131551
rect -12410 -131595 -12354 -131551
rect -12310 -131595 -12254 -131551
rect -12210 -131595 -12154 -131551
rect -12110 -131595 -12054 -131551
rect -12010 -131595 -11954 -131551
rect -11910 -131595 -11854 -131551
rect -11810 -131595 -11354 -131551
rect -11310 -131595 -11254 -131551
rect -11210 -131595 -11154 -131551
rect -11110 -131595 -11054 -131551
rect -11010 -131595 -10954 -131551
rect -10910 -131595 -10854 -131551
rect -10810 -131595 -10754 -131551
rect -10710 -131595 -10654 -131551
rect -10610 -131595 -10554 -131551
rect -10510 -131595 -10454 -131551
rect -10410 -131595 -10354 -131551
rect -10310 -131595 -10254 -131551
rect -10210 -131595 -10154 -131551
rect -10110 -131595 -10054 -131551
rect -10010 -131595 -9954 -131551
rect -9910 -131595 -9854 -131551
rect -9810 -131595 -9354 -131551
rect -9310 -131595 -9254 -131551
rect -9210 -131595 -9154 -131551
rect -9110 -131595 -9054 -131551
rect -9010 -131595 -8954 -131551
rect -8910 -131595 -8854 -131551
rect -8810 -131595 -8754 -131551
rect -8710 -131595 -8654 -131551
rect -8610 -131595 -8554 -131551
rect -8510 -131595 -8454 -131551
rect -8410 -131595 -8354 -131551
rect -8310 -131595 -8254 -131551
rect -8210 -131595 -8154 -131551
rect -8110 -131595 -8054 -131551
rect -8010 -131595 -7954 -131551
rect -7910 -131595 -7854 -131551
rect -7810 -131595 -7354 -131551
rect -7310 -131595 -7254 -131551
rect -7210 -131595 -7154 -131551
rect -7110 -131595 -7054 -131551
rect -7010 -131595 -6954 -131551
rect -6910 -131595 -6854 -131551
rect -6810 -131595 -6754 -131551
rect -6710 -131595 -6654 -131551
rect -6610 -131595 -6554 -131551
rect -6510 -131595 -6454 -131551
rect -6410 -131595 -6354 -131551
rect -6310 -131595 -6254 -131551
rect -6210 -131595 -6154 -131551
rect -6110 -131595 -6054 -131551
rect -6010 -131595 -5954 -131551
rect -5910 -131595 -5854 -131551
rect -5810 -131585 177664 -131551
rect -5810 -131595 37387 -131585
rect -108812 -131629 37387 -131595
rect 37431 -131629 37487 -131585
rect 37531 -131629 37587 -131585
rect 37631 -131629 37687 -131585
rect 37731 -131629 37787 -131585
rect 37831 -131629 37887 -131585
rect 37931 -131629 37987 -131585
rect 38031 -131629 38087 -131585
rect 38131 -131629 38187 -131585
rect 38231 -131629 38287 -131585
rect 38331 -131629 38387 -131585
rect 38431 -131629 38487 -131585
rect 38531 -131629 38587 -131585
rect 38631 -131629 38687 -131585
rect 38731 -131629 38787 -131585
rect 38831 -131629 38887 -131585
rect 38931 -131629 39387 -131585
rect 39431 -131629 39487 -131585
rect 39531 -131629 39587 -131585
rect 39631 -131629 39687 -131585
rect 39731 -131629 39787 -131585
rect 39831 -131629 39887 -131585
rect 39931 -131629 39987 -131585
rect 40031 -131629 40087 -131585
rect 40131 -131629 40187 -131585
rect 40231 -131629 40287 -131585
rect 40331 -131629 40387 -131585
rect 40431 -131629 40487 -131585
rect 40531 -131629 40587 -131585
rect 40631 -131629 40687 -131585
rect 40731 -131629 40787 -131585
rect 40831 -131629 40887 -131585
rect 40931 -131629 41387 -131585
rect 41431 -131629 41487 -131585
rect 41531 -131629 41587 -131585
rect 41631 -131629 41687 -131585
rect 41731 -131629 41787 -131585
rect 41831 -131629 41887 -131585
rect 41931 -131629 41987 -131585
rect 42031 -131629 42087 -131585
rect 42131 -131629 42187 -131585
rect 42231 -131629 42287 -131585
rect 42331 -131629 42387 -131585
rect 42431 -131629 42487 -131585
rect 42531 -131629 42587 -131585
rect 42631 -131629 42687 -131585
rect 42731 -131629 42787 -131585
rect 42831 -131629 42887 -131585
rect 42931 -131629 43387 -131585
rect 43431 -131629 43487 -131585
rect 43531 -131629 43587 -131585
rect 43631 -131629 43687 -131585
rect 43731 -131629 43787 -131585
rect 43831 -131629 43887 -131585
rect 43931 -131629 43987 -131585
rect 44031 -131629 44087 -131585
rect 44131 -131629 44187 -131585
rect 44231 -131629 44287 -131585
rect 44331 -131629 44387 -131585
rect 44431 -131629 44487 -131585
rect 44531 -131629 44587 -131585
rect 44631 -131629 44687 -131585
rect 44731 -131629 44787 -131585
rect 44831 -131629 44887 -131585
rect 44931 -131629 177664 -131585
rect -108812 -131651 177664 -131629
rect -108812 -131695 -13354 -131651
rect -13310 -131695 -13254 -131651
rect -13210 -131695 -13154 -131651
rect -13110 -131695 -13054 -131651
rect -13010 -131695 -12954 -131651
rect -12910 -131695 -12854 -131651
rect -12810 -131695 -12754 -131651
rect -12710 -131695 -12654 -131651
rect -12610 -131695 -12554 -131651
rect -12510 -131695 -12454 -131651
rect -12410 -131695 -12354 -131651
rect -12310 -131695 -12254 -131651
rect -12210 -131695 -12154 -131651
rect -12110 -131695 -12054 -131651
rect -12010 -131695 -11954 -131651
rect -11910 -131695 -11854 -131651
rect -11810 -131695 -11354 -131651
rect -11310 -131695 -11254 -131651
rect -11210 -131695 -11154 -131651
rect -11110 -131695 -11054 -131651
rect -11010 -131695 -10954 -131651
rect -10910 -131695 -10854 -131651
rect -10810 -131695 -10754 -131651
rect -10710 -131695 -10654 -131651
rect -10610 -131695 -10554 -131651
rect -10510 -131695 -10454 -131651
rect -10410 -131695 -10354 -131651
rect -10310 -131695 -10254 -131651
rect -10210 -131695 -10154 -131651
rect -10110 -131695 -10054 -131651
rect -10010 -131695 -9954 -131651
rect -9910 -131695 -9854 -131651
rect -9810 -131695 -9354 -131651
rect -9310 -131695 -9254 -131651
rect -9210 -131695 -9154 -131651
rect -9110 -131695 -9054 -131651
rect -9010 -131695 -8954 -131651
rect -8910 -131695 -8854 -131651
rect -8810 -131695 -8754 -131651
rect -8710 -131695 -8654 -131651
rect -8610 -131695 -8554 -131651
rect -8510 -131695 -8454 -131651
rect -8410 -131695 -8354 -131651
rect -8310 -131695 -8254 -131651
rect -8210 -131695 -8154 -131651
rect -8110 -131695 -8054 -131651
rect -8010 -131695 -7954 -131651
rect -7910 -131695 -7854 -131651
rect -7810 -131695 -7354 -131651
rect -7310 -131695 -7254 -131651
rect -7210 -131695 -7154 -131651
rect -7110 -131695 -7054 -131651
rect -7010 -131695 -6954 -131651
rect -6910 -131695 -6854 -131651
rect -6810 -131695 -6754 -131651
rect -6710 -131695 -6654 -131651
rect -6610 -131695 -6554 -131651
rect -6510 -131695 -6454 -131651
rect -6410 -131695 -6354 -131651
rect -6310 -131695 -6254 -131651
rect -6210 -131695 -6154 -131651
rect -6110 -131695 -6054 -131651
rect -6010 -131695 -5954 -131651
rect -5910 -131695 -5854 -131651
rect -5810 -131685 177664 -131651
rect -5810 -131695 37387 -131685
rect -108812 -131729 37387 -131695
rect 37431 -131729 37487 -131685
rect 37531 -131729 37587 -131685
rect 37631 -131729 37687 -131685
rect 37731 -131729 37787 -131685
rect 37831 -131729 37887 -131685
rect 37931 -131729 37987 -131685
rect 38031 -131729 38087 -131685
rect 38131 -131729 38187 -131685
rect 38231 -131729 38287 -131685
rect 38331 -131729 38387 -131685
rect 38431 -131729 38487 -131685
rect 38531 -131729 38587 -131685
rect 38631 -131729 38687 -131685
rect 38731 -131729 38787 -131685
rect 38831 -131729 38887 -131685
rect 38931 -131729 39387 -131685
rect 39431 -131729 39487 -131685
rect 39531 -131729 39587 -131685
rect 39631 -131729 39687 -131685
rect 39731 -131729 39787 -131685
rect 39831 -131729 39887 -131685
rect 39931 -131729 39987 -131685
rect 40031 -131729 40087 -131685
rect 40131 -131729 40187 -131685
rect 40231 -131729 40287 -131685
rect 40331 -131729 40387 -131685
rect 40431 -131729 40487 -131685
rect 40531 -131729 40587 -131685
rect 40631 -131729 40687 -131685
rect 40731 -131729 40787 -131685
rect 40831 -131729 40887 -131685
rect 40931 -131729 41387 -131685
rect 41431 -131729 41487 -131685
rect 41531 -131729 41587 -131685
rect 41631 -131729 41687 -131685
rect 41731 -131729 41787 -131685
rect 41831 -131729 41887 -131685
rect 41931 -131729 41987 -131685
rect 42031 -131729 42087 -131685
rect 42131 -131729 42187 -131685
rect 42231 -131729 42287 -131685
rect 42331 -131729 42387 -131685
rect 42431 -131729 42487 -131685
rect 42531 -131729 42587 -131685
rect 42631 -131729 42687 -131685
rect 42731 -131729 42787 -131685
rect 42831 -131729 42887 -131685
rect 42931 -131729 43387 -131685
rect 43431 -131729 43487 -131685
rect 43531 -131729 43587 -131685
rect 43631 -131729 43687 -131685
rect 43731 -131729 43787 -131685
rect 43831 -131729 43887 -131685
rect 43931 -131729 43987 -131685
rect 44031 -131729 44087 -131685
rect 44131 -131729 44187 -131685
rect 44231 -131729 44287 -131685
rect 44331 -131729 44387 -131685
rect 44431 -131729 44487 -131685
rect 44531 -131729 44587 -131685
rect 44631 -131729 44687 -131685
rect 44731 -131729 44787 -131685
rect 44831 -131729 44887 -131685
rect 44931 -131729 177664 -131685
rect -108812 -131751 177664 -131729
rect -108812 -131795 -13354 -131751
rect -13310 -131795 -13254 -131751
rect -13210 -131795 -13154 -131751
rect -13110 -131795 -13054 -131751
rect -13010 -131795 -12954 -131751
rect -12910 -131795 -12854 -131751
rect -12810 -131795 -12754 -131751
rect -12710 -131795 -12654 -131751
rect -12610 -131795 -12554 -131751
rect -12510 -131795 -12454 -131751
rect -12410 -131795 -12354 -131751
rect -12310 -131795 -12254 -131751
rect -12210 -131795 -12154 -131751
rect -12110 -131795 -12054 -131751
rect -12010 -131795 -11954 -131751
rect -11910 -131795 -11854 -131751
rect -11810 -131795 -11354 -131751
rect -11310 -131795 -11254 -131751
rect -11210 -131795 -11154 -131751
rect -11110 -131795 -11054 -131751
rect -11010 -131795 -10954 -131751
rect -10910 -131795 -10854 -131751
rect -10810 -131795 -10754 -131751
rect -10710 -131795 -10654 -131751
rect -10610 -131795 -10554 -131751
rect -10510 -131795 -10454 -131751
rect -10410 -131795 -10354 -131751
rect -10310 -131795 -10254 -131751
rect -10210 -131795 -10154 -131751
rect -10110 -131795 -10054 -131751
rect -10010 -131795 -9954 -131751
rect -9910 -131795 -9854 -131751
rect -9810 -131795 -9354 -131751
rect -9310 -131795 -9254 -131751
rect -9210 -131795 -9154 -131751
rect -9110 -131795 -9054 -131751
rect -9010 -131795 -8954 -131751
rect -8910 -131795 -8854 -131751
rect -8810 -131795 -8754 -131751
rect -8710 -131795 -8654 -131751
rect -8610 -131795 -8554 -131751
rect -8510 -131795 -8454 -131751
rect -8410 -131795 -8354 -131751
rect -8310 -131795 -8254 -131751
rect -8210 -131795 -8154 -131751
rect -8110 -131795 -8054 -131751
rect -8010 -131795 -7954 -131751
rect -7910 -131795 -7854 -131751
rect -7810 -131795 -7354 -131751
rect -7310 -131795 -7254 -131751
rect -7210 -131795 -7154 -131751
rect -7110 -131795 -7054 -131751
rect -7010 -131795 -6954 -131751
rect -6910 -131795 -6854 -131751
rect -6810 -131795 -6754 -131751
rect -6710 -131795 -6654 -131751
rect -6610 -131795 -6554 -131751
rect -6510 -131795 -6454 -131751
rect -6410 -131795 -6354 -131751
rect -6310 -131795 -6254 -131751
rect -6210 -131795 -6154 -131751
rect -6110 -131795 -6054 -131751
rect -6010 -131795 -5954 -131751
rect -5910 -131795 -5854 -131751
rect -5810 -131785 177664 -131751
rect -5810 -131795 37387 -131785
rect -108812 -131829 37387 -131795
rect 37431 -131829 37487 -131785
rect 37531 -131829 37587 -131785
rect 37631 -131829 37687 -131785
rect 37731 -131829 37787 -131785
rect 37831 -131829 37887 -131785
rect 37931 -131829 37987 -131785
rect 38031 -131829 38087 -131785
rect 38131 -131829 38187 -131785
rect 38231 -131829 38287 -131785
rect 38331 -131829 38387 -131785
rect 38431 -131829 38487 -131785
rect 38531 -131829 38587 -131785
rect 38631 -131829 38687 -131785
rect 38731 -131829 38787 -131785
rect 38831 -131829 38887 -131785
rect 38931 -131829 39387 -131785
rect 39431 -131829 39487 -131785
rect 39531 -131829 39587 -131785
rect 39631 -131829 39687 -131785
rect 39731 -131829 39787 -131785
rect 39831 -131829 39887 -131785
rect 39931 -131829 39987 -131785
rect 40031 -131829 40087 -131785
rect 40131 -131829 40187 -131785
rect 40231 -131829 40287 -131785
rect 40331 -131829 40387 -131785
rect 40431 -131829 40487 -131785
rect 40531 -131829 40587 -131785
rect 40631 -131829 40687 -131785
rect 40731 -131829 40787 -131785
rect 40831 -131829 40887 -131785
rect 40931 -131829 41387 -131785
rect 41431 -131829 41487 -131785
rect 41531 -131829 41587 -131785
rect 41631 -131829 41687 -131785
rect 41731 -131829 41787 -131785
rect 41831 -131829 41887 -131785
rect 41931 -131829 41987 -131785
rect 42031 -131829 42087 -131785
rect 42131 -131829 42187 -131785
rect 42231 -131829 42287 -131785
rect 42331 -131829 42387 -131785
rect 42431 -131829 42487 -131785
rect 42531 -131829 42587 -131785
rect 42631 -131829 42687 -131785
rect 42731 -131829 42787 -131785
rect 42831 -131829 42887 -131785
rect 42931 -131829 43387 -131785
rect 43431 -131829 43487 -131785
rect 43531 -131829 43587 -131785
rect 43631 -131829 43687 -131785
rect 43731 -131829 43787 -131785
rect 43831 -131829 43887 -131785
rect 43931 -131829 43987 -131785
rect 44031 -131829 44087 -131785
rect 44131 -131829 44187 -131785
rect 44231 -131829 44287 -131785
rect 44331 -131829 44387 -131785
rect 44431 -131829 44487 -131785
rect 44531 -131829 44587 -131785
rect 44631 -131829 44687 -131785
rect 44731 -131829 44787 -131785
rect 44831 -131829 44887 -131785
rect 44931 -131829 177664 -131785
rect -108812 -131851 177664 -131829
rect -108812 -131895 -13354 -131851
rect -13310 -131895 -13254 -131851
rect -13210 -131895 -13154 -131851
rect -13110 -131895 -13054 -131851
rect -13010 -131895 -12954 -131851
rect -12910 -131895 -12854 -131851
rect -12810 -131895 -12754 -131851
rect -12710 -131895 -12654 -131851
rect -12610 -131895 -12554 -131851
rect -12510 -131895 -12454 -131851
rect -12410 -131895 -12354 -131851
rect -12310 -131895 -12254 -131851
rect -12210 -131895 -12154 -131851
rect -12110 -131895 -12054 -131851
rect -12010 -131895 -11954 -131851
rect -11910 -131895 -11854 -131851
rect -11810 -131895 -11354 -131851
rect -11310 -131895 -11254 -131851
rect -11210 -131895 -11154 -131851
rect -11110 -131895 -11054 -131851
rect -11010 -131895 -10954 -131851
rect -10910 -131895 -10854 -131851
rect -10810 -131895 -10754 -131851
rect -10710 -131895 -10654 -131851
rect -10610 -131895 -10554 -131851
rect -10510 -131895 -10454 -131851
rect -10410 -131895 -10354 -131851
rect -10310 -131895 -10254 -131851
rect -10210 -131895 -10154 -131851
rect -10110 -131895 -10054 -131851
rect -10010 -131895 -9954 -131851
rect -9910 -131895 -9854 -131851
rect -9810 -131895 -9354 -131851
rect -9310 -131895 -9254 -131851
rect -9210 -131895 -9154 -131851
rect -9110 -131895 -9054 -131851
rect -9010 -131895 -8954 -131851
rect -8910 -131895 -8854 -131851
rect -8810 -131895 -8754 -131851
rect -8710 -131895 -8654 -131851
rect -8610 -131895 -8554 -131851
rect -8510 -131895 -8454 -131851
rect -8410 -131895 -8354 -131851
rect -8310 -131895 -8254 -131851
rect -8210 -131895 -8154 -131851
rect -8110 -131895 -8054 -131851
rect -8010 -131895 -7954 -131851
rect -7910 -131895 -7854 -131851
rect -7810 -131895 -7354 -131851
rect -7310 -131895 -7254 -131851
rect -7210 -131895 -7154 -131851
rect -7110 -131895 -7054 -131851
rect -7010 -131895 -6954 -131851
rect -6910 -131895 -6854 -131851
rect -6810 -131895 -6754 -131851
rect -6710 -131895 -6654 -131851
rect -6610 -131895 -6554 -131851
rect -6510 -131895 -6454 -131851
rect -6410 -131895 -6354 -131851
rect -6310 -131895 -6254 -131851
rect -6210 -131895 -6154 -131851
rect -6110 -131895 -6054 -131851
rect -6010 -131895 -5954 -131851
rect -5910 -131895 -5854 -131851
rect -5810 -131885 177664 -131851
rect -5810 -131895 37387 -131885
rect -108812 -131929 37387 -131895
rect 37431 -131929 37487 -131885
rect 37531 -131929 37587 -131885
rect 37631 -131929 37687 -131885
rect 37731 -131929 37787 -131885
rect 37831 -131929 37887 -131885
rect 37931 -131929 37987 -131885
rect 38031 -131929 38087 -131885
rect 38131 -131929 38187 -131885
rect 38231 -131929 38287 -131885
rect 38331 -131929 38387 -131885
rect 38431 -131929 38487 -131885
rect 38531 -131929 38587 -131885
rect 38631 -131929 38687 -131885
rect 38731 -131929 38787 -131885
rect 38831 -131929 38887 -131885
rect 38931 -131929 39387 -131885
rect 39431 -131929 39487 -131885
rect 39531 -131929 39587 -131885
rect 39631 -131929 39687 -131885
rect 39731 -131929 39787 -131885
rect 39831 -131929 39887 -131885
rect 39931 -131929 39987 -131885
rect 40031 -131929 40087 -131885
rect 40131 -131929 40187 -131885
rect 40231 -131929 40287 -131885
rect 40331 -131929 40387 -131885
rect 40431 -131929 40487 -131885
rect 40531 -131929 40587 -131885
rect 40631 -131929 40687 -131885
rect 40731 -131929 40787 -131885
rect 40831 -131929 40887 -131885
rect 40931 -131929 41387 -131885
rect 41431 -131929 41487 -131885
rect 41531 -131929 41587 -131885
rect 41631 -131929 41687 -131885
rect 41731 -131929 41787 -131885
rect 41831 -131929 41887 -131885
rect 41931 -131929 41987 -131885
rect 42031 -131929 42087 -131885
rect 42131 -131929 42187 -131885
rect 42231 -131929 42287 -131885
rect 42331 -131929 42387 -131885
rect 42431 -131929 42487 -131885
rect 42531 -131929 42587 -131885
rect 42631 -131929 42687 -131885
rect 42731 -131929 42787 -131885
rect 42831 -131929 42887 -131885
rect 42931 -131929 43387 -131885
rect 43431 -131929 43487 -131885
rect 43531 -131929 43587 -131885
rect 43631 -131929 43687 -131885
rect 43731 -131929 43787 -131885
rect 43831 -131929 43887 -131885
rect 43931 -131929 43987 -131885
rect 44031 -131929 44087 -131885
rect 44131 -131929 44187 -131885
rect 44231 -131929 44287 -131885
rect 44331 -131929 44387 -131885
rect 44431 -131929 44487 -131885
rect 44531 -131929 44587 -131885
rect 44631 -131929 44687 -131885
rect 44731 -131929 44787 -131885
rect 44831 -131929 44887 -131885
rect 44931 -131929 177664 -131885
rect -108812 -131951 177664 -131929
rect -108812 -131995 -13354 -131951
rect -13310 -131995 -13254 -131951
rect -13210 -131995 -13154 -131951
rect -13110 -131995 -13054 -131951
rect -13010 -131995 -12954 -131951
rect -12910 -131995 -12854 -131951
rect -12810 -131995 -12754 -131951
rect -12710 -131995 -12654 -131951
rect -12610 -131995 -12554 -131951
rect -12510 -131995 -12454 -131951
rect -12410 -131995 -12354 -131951
rect -12310 -131995 -12254 -131951
rect -12210 -131995 -12154 -131951
rect -12110 -131995 -12054 -131951
rect -12010 -131995 -11954 -131951
rect -11910 -131995 -11854 -131951
rect -11810 -131995 -11354 -131951
rect -11310 -131995 -11254 -131951
rect -11210 -131995 -11154 -131951
rect -11110 -131995 -11054 -131951
rect -11010 -131995 -10954 -131951
rect -10910 -131995 -10854 -131951
rect -10810 -131995 -10754 -131951
rect -10710 -131995 -10654 -131951
rect -10610 -131995 -10554 -131951
rect -10510 -131995 -10454 -131951
rect -10410 -131995 -10354 -131951
rect -10310 -131995 -10254 -131951
rect -10210 -131995 -10154 -131951
rect -10110 -131995 -10054 -131951
rect -10010 -131995 -9954 -131951
rect -9910 -131995 -9854 -131951
rect -9810 -131995 -9354 -131951
rect -9310 -131995 -9254 -131951
rect -9210 -131995 -9154 -131951
rect -9110 -131995 -9054 -131951
rect -9010 -131995 -8954 -131951
rect -8910 -131995 -8854 -131951
rect -8810 -131995 -8754 -131951
rect -8710 -131995 -8654 -131951
rect -8610 -131995 -8554 -131951
rect -8510 -131995 -8454 -131951
rect -8410 -131995 -8354 -131951
rect -8310 -131995 -8254 -131951
rect -8210 -131995 -8154 -131951
rect -8110 -131995 -8054 -131951
rect -8010 -131995 -7954 -131951
rect -7910 -131995 -7854 -131951
rect -7810 -131995 -7354 -131951
rect -7310 -131995 -7254 -131951
rect -7210 -131995 -7154 -131951
rect -7110 -131995 -7054 -131951
rect -7010 -131995 -6954 -131951
rect -6910 -131995 -6854 -131951
rect -6810 -131995 -6754 -131951
rect -6710 -131995 -6654 -131951
rect -6610 -131995 -6554 -131951
rect -6510 -131995 -6454 -131951
rect -6410 -131995 -6354 -131951
rect -6310 -131995 -6254 -131951
rect -6210 -131995 -6154 -131951
rect -6110 -131995 -6054 -131951
rect -6010 -131995 -5954 -131951
rect -5910 -131995 -5854 -131951
rect -5810 -131985 177664 -131951
rect -5810 -131995 37387 -131985
rect -108812 -132029 37387 -131995
rect 37431 -132029 37487 -131985
rect 37531 -132029 37587 -131985
rect 37631 -132029 37687 -131985
rect 37731 -132029 37787 -131985
rect 37831 -132029 37887 -131985
rect 37931 -132029 37987 -131985
rect 38031 -132029 38087 -131985
rect 38131 -132029 38187 -131985
rect 38231 -132029 38287 -131985
rect 38331 -132029 38387 -131985
rect 38431 -132029 38487 -131985
rect 38531 -132029 38587 -131985
rect 38631 -132029 38687 -131985
rect 38731 -132029 38787 -131985
rect 38831 -132029 38887 -131985
rect 38931 -132029 39387 -131985
rect 39431 -132029 39487 -131985
rect 39531 -132029 39587 -131985
rect 39631 -132029 39687 -131985
rect 39731 -132029 39787 -131985
rect 39831 -132029 39887 -131985
rect 39931 -132029 39987 -131985
rect 40031 -132029 40087 -131985
rect 40131 -132029 40187 -131985
rect 40231 -132029 40287 -131985
rect 40331 -132029 40387 -131985
rect 40431 -132029 40487 -131985
rect 40531 -132029 40587 -131985
rect 40631 -132029 40687 -131985
rect 40731 -132029 40787 -131985
rect 40831 -132029 40887 -131985
rect 40931 -132029 41387 -131985
rect 41431 -132029 41487 -131985
rect 41531 -132029 41587 -131985
rect 41631 -132029 41687 -131985
rect 41731 -132029 41787 -131985
rect 41831 -132029 41887 -131985
rect 41931 -132029 41987 -131985
rect 42031 -132029 42087 -131985
rect 42131 -132029 42187 -131985
rect 42231 -132029 42287 -131985
rect 42331 -132029 42387 -131985
rect 42431 -132029 42487 -131985
rect 42531 -132029 42587 -131985
rect 42631 -132029 42687 -131985
rect 42731 -132029 42787 -131985
rect 42831 -132029 42887 -131985
rect 42931 -132029 43387 -131985
rect 43431 -132029 43487 -131985
rect 43531 -132029 43587 -131985
rect 43631 -132029 43687 -131985
rect 43731 -132029 43787 -131985
rect 43831 -132029 43887 -131985
rect 43931 -132029 43987 -131985
rect 44031 -132029 44087 -131985
rect 44131 -132029 44187 -131985
rect 44231 -132029 44287 -131985
rect 44331 -132029 44387 -131985
rect 44431 -132029 44487 -131985
rect 44531 -132029 44587 -131985
rect 44631 -132029 44687 -131985
rect 44731 -132029 44787 -131985
rect 44831 -132029 44887 -131985
rect 44931 -132029 177664 -131985
rect -108812 -132051 177664 -132029
rect -108812 -132095 -13354 -132051
rect -13310 -132095 -13254 -132051
rect -13210 -132095 -13154 -132051
rect -13110 -132095 -13054 -132051
rect -13010 -132095 -12954 -132051
rect -12910 -132095 -12854 -132051
rect -12810 -132095 -12754 -132051
rect -12710 -132095 -12654 -132051
rect -12610 -132095 -12554 -132051
rect -12510 -132095 -12454 -132051
rect -12410 -132095 -12354 -132051
rect -12310 -132095 -12254 -132051
rect -12210 -132095 -12154 -132051
rect -12110 -132095 -12054 -132051
rect -12010 -132095 -11954 -132051
rect -11910 -132095 -11854 -132051
rect -11810 -132095 -11354 -132051
rect -11310 -132095 -11254 -132051
rect -11210 -132095 -11154 -132051
rect -11110 -132095 -11054 -132051
rect -11010 -132095 -10954 -132051
rect -10910 -132095 -10854 -132051
rect -10810 -132095 -10754 -132051
rect -10710 -132095 -10654 -132051
rect -10610 -132095 -10554 -132051
rect -10510 -132095 -10454 -132051
rect -10410 -132095 -10354 -132051
rect -10310 -132095 -10254 -132051
rect -10210 -132095 -10154 -132051
rect -10110 -132095 -10054 -132051
rect -10010 -132095 -9954 -132051
rect -9910 -132095 -9854 -132051
rect -9810 -132095 -9354 -132051
rect -9310 -132095 -9254 -132051
rect -9210 -132095 -9154 -132051
rect -9110 -132095 -9054 -132051
rect -9010 -132095 -8954 -132051
rect -8910 -132095 -8854 -132051
rect -8810 -132095 -8754 -132051
rect -8710 -132095 -8654 -132051
rect -8610 -132095 -8554 -132051
rect -8510 -132095 -8454 -132051
rect -8410 -132095 -8354 -132051
rect -8310 -132095 -8254 -132051
rect -8210 -132095 -8154 -132051
rect -8110 -132095 -8054 -132051
rect -8010 -132095 -7954 -132051
rect -7910 -132095 -7854 -132051
rect -7810 -132095 -7354 -132051
rect -7310 -132095 -7254 -132051
rect -7210 -132095 -7154 -132051
rect -7110 -132095 -7054 -132051
rect -7010 -132095 -6954 -132051
rect -6910 -132095 -6854 -132051
rect -6810 -132095 -6754 -132051
rect -6710 -132095 -6654 -132051
rect -6610 -132095 -6554 -132051
rect -6510 -132095 -6454 -132051
rect -6410 -132095 -6354 -132051
rect -6310 -132095 -6254 -132051
rect -6210 -132095 -6154 -132051
rect -6110 -132095 -6054 -132051
rect -6010 -132095 -5954 -132051
rect -5910 -132095 -5854 -132051
rect -5810 -132085 177664 -132051
rect -5810 -132095 37387 -132085
rect -108812 -132129 37387 -132095
rect 37431 -132129 37487 -132085
rect 37531 -132129 37587 -132085
rect 37631 -132129 37687 -132085
rect 37731 -132129 37787 -132085
rect 37831 -132129 37887 -132085
rect 37931 -132129 37987 -132085
rect 38031 -132129 38087 -132085
rect 38131 -132129 38187 -132085
rect 38231 -132129 38287 -132085
rect 38331 -132129 38387 -132085
rect 38431 -132129 38487 -132085
rect 38531 -132129 38587 -132085
rect 38631 -132129 38687 -132085
rect 38731 -132129 38787 -132085
rect 38831 -132129 38887 -132085
rect 38931 -132129 39387 -132085
rect 39431 -132129 39487 -132085
rect 39531 -132129 39587 -132085
rect 39631 -132129 39687 -132085
rect 39731 -132129 39787 -132085
rect 39831 -132129 39887 -132085
rect 39931 -132129 39987 -132085
rect 40031 -132129 40087 -132085
rect 40131 -132129 40187 -132085
rect 40231 -132129 40287 -132085
rect 40331 -132129 40387 -132085
rect 40431 -132129 40487 -132085
rect 40531 -132129 40587 -132085
rect 40631 -132129 40687 -132085
rect 40731 -132129 40787 -132085
rect 40831 -132129 40887 -132085
rect 40931 -132129 41387 -132085
rect 41431 -132129 41487 -132085
rect 41531 -132129 41587 -132085
rect 41631 -132129 41687 -132085
rect 41731 -132129 41787 -132085
rect 41831 -132129 41887 -132085
rect 41931 -132129 41987 -132085
rect 42031 -132129 42087 -132085
rect 42131 -132129 42187 -132085
rect 42231 -132129 42287 -132085
rect 42331 -132129 42387 -132085
rect 42431 -132129 42487 -132085
rect 42531 -132129 42587 -132085
rect 42631 -132129 42687 -132085
rect 42731 -132129 42787 -132085
rect 42831 -132129 42887 -132085
rect 42931 -132129 43387 -132085
rect 43431 -132129 43487 -132085
rect 43531 -132129 43587 -132085
rect 43631 -132129 43687 -132085
rect 43731 -132129 43787 -132085
rect 43831 -132129 43887 -132085
rect 43931 -132129 43987 -132085
rect 44031 -132129 44087 -132085
rect 44131 -132129 44187 -132085
rect 44231 -132129 44287 -132085
rect 44331 -132129 44387 -132085
rect 44431 -132129 44487 -132085
rect 44531 -132129 44587 -132085
rect 44631 -132129 44687 -132085
rect 44731 -132129 44787 -132085
rect 44831 -132129 44887 -132085
rect 44931 -132129 177664 -132085
rect -108812 -132151 177664 -132129
rect -108812 -132195 -13354 -132151
rect -13310 -132195 -13254 -132151
rect -13210 -132195 -13154 -132151
rect -13110 -132195 -13054 -132151
rect -13010 -132195 -12954 -132151
rect -12910 -132195 -12854 -132151
rect -12810 -132195 -12754 -132151
rect -12710 -132195 -12654 -132151
rect -12610 -132195 -12554 -132151
rect -12510 -132195 -12454 -132151
rect -12410 -132195 -12354 -132151
rect -12310 -132195 -12254 -132151
rect -12210 -132195 -12154 -132151
rect -12110 -132195 -12054 -132151
rect -12010 -132195 -11954 -132151
rect -11910 -132195 -11854 -132151
rect -11810 -132195 -11354 -132151
rect -11310 -132195 -11254 -132151
rect -11210 -132195 -11154 -132151
rect -11110 -132195 -11054 -132151
rect -11010 -132195 -10954 -132151
rect -10910 -132195 -10854 -132151
rect -10810 -132195 -10754 -132151
rect -10710 -132195 -10654 -132151
rect -10610 -132195 -10554 -132151
rect -10510 -132195 -10454 -132151
rect -10410 -132195 -10354 -132151
rect -10310 -132195 -10254 -132151
rect -10210 -132195 -10154 -132151
rect -10110 -132195 -10054 -132151
rect -10010 -132195 -9954 -132151
rect -9910 -132195 -9854 -132151
rect -9810 -132195 -9354 -132151
rect -9310 -132195 -9254 -132151
rect -9210 -132195 -9154 -132151
rect -9110 -132195 -9054 -132151
rect -9010 -132195 -8954 -132151
rect -8910 -132195 -8854 -132151
rect -8810 -132195 -8754 -132151
rect -8710 -132195 -8654 -132151
rect -8610 -132195 -8554 -132151
rect -8510 -132195 -8454 -132151
rect -8410 -132195 -8354 -132151
rect -8310 -132195 -8254 -132151
rect -8210 -132195 -8154 -132151
rect -8110 -132195 -8054 -132151
rect -8010 -132195 -7954 -132151
rect -7910 -132195 -7854 -132151
rect -7810 -132195 -7354 -132151
rect -7310 -132195 -7254 -132151
rect -7210 -132195 -7154 -132151
rect -7110 -132195 -7054 -132151
rect -7010 -132195 -6954 -132151
rect -6910 -132195 -6854 -132151
rect -6810 -132195 -6754 -132151
rect -6710 -132195 -6654 -132151
rect -6610 -132195 -6554 -132151
rect -6510 -132195 -6454 -132151
rect -6410 -132195 -6354 -132151
rect -6310 -132195 -6254 -132151
rect -6210 -132195 -6154 -132151
rect -6110 -132195 -6054 -132151
rect -6010 -132195 -5954 -132151
rect -5910 -132195 -5854 -132151
rect -5810 -132185 177664 -132151
rect -5810 -132195 37387 -132185
rect -108812 -132229 37387 -132195
rect 37431 -132229 37487 -132185
rect 37531 -132229 37587 -132185
rect 37631 -132229 37687 -132185
rect 37731 -132229 37787 -132185
rect 37831 -132229 37887 -132185
rect 37931 -132229 37987 -132185
rect 38031 -132229 38087 -132185
rect 38131 -132229 38187 -132185
rect 38231 -132229 38287 -132185
rect 38331 -132229 38387 -132185
rect 38431 -132229 38487 -132185
rect 38531 -132229 38587 -132185
rect 38631 -132229 38687 -132185
rect 38731 -132229 38787 -132185
rect 38831 -132229 38887 -132185
rect 38931 -132229 39387 -132185
rect 39431 -132229 39487 -132185
rect 39531 -132229 39587 -132185
rect 39631 -132229 39687 -132185
rect 39731 -132229 39787 -132185
rect 39831 -132229 39887 -132185
rect 39931 -132229 39987 -132185
rect 40031 -132229 40087 -132185
rect 40131 -132229 40187 -132185
rect 40231 -132229 40287 -132185
rect 40331 -132229 40387 -132185
rect 40431 -132229 40487 -132185
rect 40531 -132229 40587 -132185
rect 40631 -132229 40687 -132185
rect 40731 -132229 40787 -132185
rect 40831 -132229 40887 -132185
rect 40931 -132229 41387 -132185
rect 41431 -132229 41487 -132185
rect 41531 -132229 41587 -132185
rect 41631 -132229 41687 -132185
rect 41731 -132229 41787 -132185
rect 41831 -132229 41887 -132185
rect 41931 -132229 41987 -132185
rect 42031 -132229 42087 -132185
rect 42131 -132229 42187 -132185
rect 42231 -132229 42287 -132185
rect 42331 -132229 42387 -132185
rect 42431 -132229 42487 -132185
rect 42531 -132229 42587 -132185
rect 42631 -132229 42687 -132185
rect 42731 -132229 42787 -132185
rect 42831 -132229 42887 -132185
rect 42931 -132229 43387 -132185
rect 43431 -132229 43487 -132185
rect 43531 -132229 43587 -132185
rect 43631 -132229 43687 -132185
rect 43731 -132229 43787 -132185
rect 43831 -132229 43887 -132185
rect 43931 -132229 43987 -132185
rect 44031 -132229 44087 -132185
rect 44131 -132229 44187 -132185
rect 44231 -132229 44287 -132185
rect 44331 -132229 44387 -132185
rect 44431 -132229 44487 -132185
rect 44531 -132229 44587 -132185
rect 44631 -132229 44687 -132185
rect 44731 -132229 44787 -132185
rect 44831 -132229 44887 -132185
rect 44931 -132229 177664 -132185
rect -108812 -132251 177664 -132229
rect -108812 -132295 -13354 -132251
rect -13310 -132295 -13254 -132251
rect -13210 -132295 -13154 -132251
rect -13110 -132295 -13054 -132251
rect -13010 -132295 -12954 -132251
rect -12910 -132295 -12854 -132251
rect -12810 -132295 -12754 -132251
rect -12710 -132295 -12654 -132251
rect -12610 -132295 -12554 -132251
rect -12510 -132295 -12454 -132251
rect -12410 -132295 -12354 -132251
rect -12310 -132295 -12254 -132251
rect -12210 -132295 -12154 -132251
rect -12110 -132295 -12054 -132251
rect -12010 -132295 -11954 -132251
rect -11910 -132295 -11854 -132251
rect -11810 -132295 -11354 -132251
rect -11310 -132295 -11254 -132251
rect -11210 -132295 -11154 -132251
rect -11110 -132295 -11054 -132251
rect -11010 -132295 -10954 -132251
rect -10910 -132295 -10854 -132251
rect -10810 -132295 -10754 -132251
rect -10710 -132295 -10654 -132251
rect -10610 -132295 -10554 -132251
rect -10510 -132295 -10454 -132251
rect -10410 -132295 -10354 -132251
rect -10310 -132295 -10254 -132251
rect -10210 -132295 -10154 -132251
rect -10110 -132295 -10054 -132251
rect -10010 -132295 -9954 -132251
rect -9910 -132295 -9854 -132251
rect -9810 -132295 -9354 -132251
rect -9310 -132295 -9254 -132251
rect -9210 -132295 -9154 -132251
rect -9110 -132295 -9054 -132251
rect -9010 -132295 -8954 -132251
rect -8910 -132295 -8854 -132251
rect -8810 -132295 -8754 -132251
rect -8710 -132295 -8654 -132251
rect -8610 -132295 -8554 -132251
rect -8510 -132295 -8454 -132251
rect -8410 -132295 -8354 -132251
rect -8310 -132295 -8254 -132251
rect -8210 -132295 -8154 -132251
rect -8110 -132295 -8054 -132251
rect -8010 -132295 -7954 -132251
rect -7910 -132295 -7854 -132251
rect -7810 -132295 -7354 -132251
rect -7310 -132295 -7254 -132251
rect -7210 -132295 -7154 -132251
rect -7110 -132295 -7054 -132251
rect -7010 -132295 -6954 -132251
rect -6910 -132295 -6854 -132251
rect -6810 -132295 -6754 -132251
rect -6710 -132295 -6654 -132251
rect -6610 -132295 -6554 -132251
rect -6510 -132295 -6454 -132251
rect -6410 -132295 -6354 -132251
rect -6310 -132295 -6254 -132251
rect -6210 -132295 -6154 -132251
rect -6110 -132295 -6054 -132251
rect -6010 -132295 -5954 -132251
rect -5910 -132295 -5854 -132251
rect -5810 -132285 177664 -132251
rect -5810 -132295 37387 -132285
rect -108812 -132329 37387 -132295
rect 37431 -132329 37487 -132285
rect 37531 -132329 37587 -132285
rect 37631 -132329 37687 -132285
rect 37731 -132329 37787 -132285
rect 37831 -132329 37887 -132285
rect 37931 -132329 37987 -132285
rect 38031 -132329 38087 -132285
rect 38131 -132329 38187 -132285
rect 38231 -132329 38287 -132285
rect 38331 -132329 38387 -132285
rect 38431 -132329 38487 -132285
rect 38531 -132329 38587 -132285
rect 38631 -132329 38687 -132285
rect 38731 -132329 38787 -132285
rect 38831 -132329 38887 -132285
rect 38931 -132329 39387 -132285
rect 39431 -132329 39487 -132285
rect 39531 -132329 39587 -132285
rect 39631 -132329 39687 -132285
rect 39731 -132329 39787 -132285
rect 39831 -132329 39887 -132285
rect 39931 -132329 39987 -132285
rect 40031 -132329 40087 -132285
rect 40131 -132329 40187 -132285
rect 40231 -132329 40287 -132285
rect 40331 -132329 40387 -132285
rect 40431 -132329 40487 -132285
rect 40531 -132329 40587 -132285
rect 40631 -132329 40687 -132285
rect 40731 -132329 40787 -132285
rect 40831 -132329 40887 -132285
rect 40931 -132329 41387 -132285
rect 41431 -132329 41487 -132285
rect 41531 -132329 41587 -132285
rect 41631 -132329 41687 -132285
rect 41731 -132329 41787 -132285
rect 41831 -132329 41887 -132285
rect 41931 -132329 41987 -132285
rect 42031 -132329 42087 -132285
rect 42131 -132329 42187 -132285
rect 42231 -132329 42287 -132285
rect 42331 -132329 42387 -132285
rect 42431 -132329 42487 -132285
rect 42531 -132329 42587 -132285
rect 42631 -132329 42687 -132285
rect 42731 -132329 42787 -132285
rect 42831 -132329 42887 -132285
rect 42931 -132329 43387 -132285
rect 43431 -132329 43487 -132285
rect 43531 -132329 43587 -132285
rect 43631 -132329 43687 -132285
rect 43731 -132329 43787 -132285
rect 43831 -132329 43887 -132285
rect 43931 -132329 43987 -132285
rect 44031 -132329 44087 -132285
rect 44131 -132329 44187 -132285
rect 44231 -132329 44287 -132285
rect 44331 -132329 44387 -132285
rect 44431 -132329 44487 -132285
rect 44531 -132329 44587 -132285
rect 44631 -132329 44687 -132285
rect 44731 -132329 44787 -132285
rect 44831 -132329 44887 -132285
rect 44931 -132329 177664 -132285
rect -108812 -132351 177664 -132329
rect -108812 -132395 -13354 -132351
rect -13310 -132395 -13254 -132351
rect -13210 -132395 -13154 -132351
rect -13110 -132395 -13054 -132351
rect -13010 -132395 -12954 -132351
rect -12910 -132395 -12854 -132351
rect -12810 -132395 -12754 -132351
rect -12710 -132395 -12654 -132351
rect -12610 -132395 -12554 -132351
rect -12510 -132395 -12454 -132351
rect -12410 -132395 -12354 -132351
rect -12310 -132395 -12254 -132351
rect -12210 -132395 -12154 -132351
rect -12110 -132395 -12054 -132351
rect -12010 -132395 -11954 -132351
rect -11910 -132395 -11854 -132351
rect -11810 -132395 -11354 -132351
rect -11310 -132395 -11254 -132351
rect -11210 -132395 -11154 -132351
rect -11110 -132395 -11054 -132351
rect -11010 -132395 -10954 -132351
rect -10910 -132395 -10854 -132351
rect -10810 -132395 -10754 -132351
rect -10710 -132395 -10654 -132351
rect -10610 -132395 -10554 -132351
rect -10510 -132395 -10454 -132351
rect -10410 -132395 -10354 -132351
rect -10310 -132395 -10254 -132351
rect -10210 -132395 -10154 -132351
rect -10110 -132395 -10054 -132351
rect -10010 -132395 -9954 -132351
rect -9910 -132395 -9854 -132351
rect -9810 -132395 -9354 -132351
rect -9310 -132395 -9254 -132351
rect -9210 -132395 -9154 -132351
rect -9110 -132395 -9054 -132351
rect -9010 -132395 -8954 -132351
rect -8910 -132395 -8854 -132351
rect -8810 -132395 -8754 -132351
rect -8710 -132395 -8654 -132351
rect -8610 -132395 -8554 -132351
rect -8510 -132395 -8454 -132351
rect -8410 -132395 -8354 -132351
rect -8310 -132395 -8254 -132351
rect -8210 -132395 -8154 -132351
rect -8110 -132395 -8054 -132351
rect -8010 -132395 -7954 -132351
rect -7910 -132395 -7854 -132351
rect -7810 -132395 -7354 -132351
rect -7310 -132395 -7254 -132351
rect -7210 -132395 -7154 -132351
rect -7110 -132395 -7054 -132351
rect -7010 -132395 -6954 -132351
rect -6910 -132395 -6854 -132351
rect -6810 -132395 -6754 -132351
rect -6710 -132395 -6654 -132351
rect -6610 -132395 -6554 -132351
rect -6510 -132395 -6454 -132351
rect -6410 -132395 -6354 -132351
rect -6310 -132395 -6254 -132351
rect -6210 -132395 -6154 -132351
rect -6110 -132395 -6054 -132351
rect -6010 -132395 -5954 -132351
rect -5910 -132395 -5854 -132351
rect -5810 -132385 177664 -132351
rect -5810 -132395 37387 -132385
rect -108812 -132429 37387 -132395
rect 37431 -132429 37487 -132385
rect 37531 -132429 37587 -132385
rect 37631 -132429 37687 -132385
rect 37731 -132429 37787 -132385
rect 37831 -132429 37887 -132385
rect 37931 -132429 37987 -132385
rect 38031 -132429 38087 -132385
rect 38131 -132429 38187 -132385
rect 38231 -132429 38287 -132385
rect 38331 -132429 38387 -132385
rect 38431 -132429 38487 -132385
rect 38531 -132429 38587 -132385
rect 38631 -132429 38687 -132385
rect 38731 -132429 38787 -132385
rect 38831 -132429 38887 -132385
rect 38931 -132429 39387 -132385
rect 39431 -132429 39487 -132385
rect 39531 -132429 39587 -132385
rect 39631 -132429 39687 -132385
rect 39731 -132429 39787 -132385
rect 39831 -132429 39887 -132385
rect 39931 -132429 39987 -132385
rect 40031 -132429 40087 -132385
rect 40131 -132429 40187 -132385
rect 40231 -132429 40287 -132385
rect 40331 -132429 40387 -132385
rect 40431 -132429 40487 -132385
rect 40531 -132429 40587 -132385
rect 40631 -132429 40687 -132385
rect 40731 -132429 40787 -132385
rect 40831 -132429 40887 -132385
rect 40931 -132429 41387 -132385
rect 41431 -132429 41487 -132385
rect 41531 -132429 41587 -132385
rect 41631 -132429 41687 -132385
rect 41731 -132429 41787 -132385
rect 41831 -132429 41887 -132385
rect 41931 -132429 41987 -132385
rect 42031 -132429 42087 -132385
rect 42131 -132429 42187 -132385
rect 42231 -132429 42287 -132385
rect 42331 -132429 42387 -132385
rect 42431 -132429 42487 -132385
rect 42531 -132429 42587 -132385
rect 42631 -132429 42687 -132385
rect 42731 -132429 42787 -132385
rect 42831 -132429 42887 -132385
rect 42931 -132429 43387 -132385
rect 43431 -132429 43487 -132385
rect 43531 -132429 43587 -132385
rect 43631 -132429 43687 -132385
rect 43731 -132429 43787 -132385
rect 43831 -132429 43887 -132385
rect 43931 -132429 43987 -132385
rect 44031 -132429 44087 -132385
rect 44131 -132429 44187 -132385
rect 44231 -132429 44287 -132385
rect 44331 -132429 44387 -132385
rect 44431 -132429 44487 -132385
rect 44531 -132429 44587 -132385
rect 44631 -132429 44687 -132385
rect 44731 -132429 44787 -132385
rect 44831 -132429 44887 -132385
rect 44931 -132429 177664 -132385
rect -108812 -132451 177664 -132429
rect -108812 -132495 -13354 -132451
rect -13310 -132495 -13254 -132451
rect -13210 -132495 -13154 -132451
rect -13110 -132495 -13054 -132451
rect -13010 -132495 -12954 -132451
rect -12910 -132495 -12854 -132451
rect -12810 -132495 -12754 -132451
rect -12710 -132495 -12654 -132451
rect -12610 -132495 -12554 -132451
rect -12510 -132495 -12454 -132451
rect -12410 -132495 -12354 -132451
rect -12310 -132495 -12254 -132451
rect -12210 -132495 -12154 -132451
rect -12110 -132495 -12054 -132451
rect -12010 -132495 -11954 -132451
rect -11910 -132495 -11854 -132451
rect -11810 -132495 -11354 -132451
rect -11310 -132495 -11254 -132451
rect -11210 -132495 -11154 -132451
rect -11110 -132495 -11054 -132451
rect -11010 -132495 -10954 -132451
rect -10910 -132495 -10854 -132451
rect -10810 -132495 -10754 -132451
rect -10710 -132495 -10654 -132451
rect -10610 -132495 -10554 -132451
rect -10510 -132495 -10454 -132451
rect -10410 -132495 -10354 -132451
rect -10310 -132495 -10254 -132451
rect -10210 -132495 -10154 -132451
rect -10110 -132495 -10054 -132451
rect -10010 -132495 -9954 -132451
rect -9910 -132495 -9854 -132451
rect -9810 -132495 -9354 -132451
rect -9310 -132495 -9254 -132451
rect -9210 -132495 -9154 -132451
rect -9110 -132495 -9054 -132451
rect -9010 -132495 -8954 -132451
rect -8910 -132495 -8854 -132451
rect -8810 -132495 -8754 -132451
rect -8710 -132495 -8654 -132451
rect -8610 -132495 -8554 -132451
rect -8510 -132495 -8454 -132451
rect -8410 -132495 -8354 -132451
rect -8310 -132495 -8254 -132451
rect -8210 -132495 -8154 -132451
rect -8110 -132495 -8054 -132451
rect -8010 -132495 -7954 -132451
rect -7910 -132495 -7854 -132451
rect -7810 -132495 -7354 -132451
rect -7310 -132495 -7254 -132451
rect -7210 -132495 -7154 -132451
rect -7110 -132495 -7054 -132451
rect -7010 -132495 -6954 -132451
rect -6910 -132495 -6854 -132451
rect -6810 -132495 -6754 -132451
rect -6710 -132495 -6654 -132451
rect -6610 -132495 -6554 -132451
rect -6510 -132495 -6454 -132451
rect -6410 -132495 -6354 -132451
rect -6310 -132495 -6254 -132451
rect -6210 -132495 -6154 -132451
rect -6110 -132495 -6054 -132451
rect -6010 -132495 -5954 -132451
rect -5910 -132495 -5854 -132451
rect -5810 -132485 177664 -132451
rect -5810 -132495 37387 -132485
rect -108812 -132529 37387 -132495
rect 37431 -132529 37487 -132485
rect 37531 -132529 37587 -132485
rect 37631 -132529 37687 -132485
rect 37731 -132529 37787 -132485
rect 37831 -132529 37887 -132485
rect 37931 -132529 37987 -132485
rect 38031 -132529 38087 -132485
rect 38131 -132529 38187 -132485
rect 38231 -132529 38287 -132485
rect 38331 -132529 38387 -132485
rect 38431 -132529 38487 -132485
rect 38531 -132529 38587 -132485
rect 38631 -132529 38687 -132485
rect 38731 -132529 38787 -132485
rect 38831 -132529 38887 -132485
rect 38931 -132529 39387 -132485
rect 39431 -132529 39487 -132485
rect 39531 -132529 39587 -132485
rect 39631 -132529 39687 -132485
rect 39731 -132529 39787 -132485
rect 39831 -132529 39887 -132485
rect 39931 -132529 39987 -132485
rect 40031 -132529 40087 -132485
rect 40131 -132529 40187 -132485
rect 40231 -132529 40287 -132485
rect 40331 -132529 40387 -132485
rect 40431 -132529 40487 -132485
rect 40531 -132529 40587 -132485
rect 40631 -132529 40687 -132485
rect 40731 -132529 40787 -132485
rect 40831 -132529 40887 -132485
rect 40931 -132529 41387 -132485
rect 41431 -132529 41487 -132485
rect 41531 -132529 41587 -132485
rect 41631 -132529 41687 -132485
rect 41731 -132529 41787 -132485
rect 41831 -132529 41887 -132485
rect 41931 -132529 41987 -132485
rect 42031 -132529 42087 -132485
rect 42131 -132529 42187 -132485
rect 42231 -132529 42287 -132485
rect 42331 -132529 42387 -132485
rect 42431 -132529 42487 -132485
rect 42531 -132529 42587 -132485
rect 42631 -132529 42687 -132485
rect 42731 -132529 42787 -132485
rect 42831 -132529 42887 -132485
rect 42931 -132529 43387 -132485
rect 43431 -132529 43487 -132485
rect 43531 -132529 43587 -132485
rect 43631 -132529 43687 -132485
rect 43731 -132529 43787 -132485
rect 43831 -132529 43887 -132485
rect 43931 -132529 43987 -132485
rect 44031 -132529 44087 -132485
rect 44131 -132529 44187 -132485
rect 44231 -132529 44287 -132485
rect 44331 -132529 44387 -132485
rect 44431 -132529 44487 -132485
rect 44531 -132529 44587 -132485
rect 44631 -132529 44687 -132485
rect 44731 -132529 44787 -132485
rect 44831 -132529 44887 -132485
rect 44931 -132529 177664 -132485
rect -108812 -132551 177664 -132529
rect -108812 -132595 -13354 -132551
rect -13310 -132595 -13254 -132551
rect -13210 -132595 -13154 -132551
rect -13110 -132595 -13054 -132551
rect -13010 -132595 -12954 -132551
rect -12910 -132595 -12854 -132551
rect -12810 -132595 -12754 -132551
rect -12710 -132595 -12654 -132551
rect -12610 -132595 -12554 -132551
rect -12510 -132595 -12454 -132551
rect -12410 -132595 -12354 -132551
rect -12310 -132595 -12254 -132551
rect -12210 -132595 -12154 -132551
rect -12110 -132595 -12054 -132551
rect -12010 -132595 -11954 -132551
rect -11910 -132595 -11854 -132551
rect -11810 -132595 -11354 -132551
rect -11310 -132595 -11254 -132551
rect -11210 -132595 -11154 -132551
rect -11110 -132595 -11054 -132551
rect -11010 -132595 -10954 -132551
rect -10910 -132595 -10854 -132551
rect -10810 -132595 -10754 -132551
rect -10710 -132595 -10654 -132551
rect -10610 -132595 -10554 -132551
rect -10510 -132595 -10454 -132551
rect -10410 -132595 -10354 -132551
rect -10310 -132595 -10254 -132551
rect -10210 -132595 -10154 -132551
rect -10110 -132595 -10054 -132551
rect -10010 -132595 -9954 -132551
rect -9910 -132595 -9854 -132551
rect -9810 -132595 -9354 -132551
rect -9310 -132595 -9254 -132551
rect -9210 -132595 -9154 -132551
rect -9110 -132595 -9054 -132551
rect -9010 -132595 -8954 -132551
rect -8910 -132595 -8854 -132551
rect -8810 -132595 -8754 -132551
rect -8710 -132595 -8654 -132551
rect -8610 -132595 -8554 -132551
rect -8510 -132595 -8454 -132551
rect -8410 -132595 -8354 -132551
rect -8310 -132595 -8254 -132551
rect -8210 -132595 -8154 -132551
rect -8110 -132595 -8054 -132551
rect -8010 -132595 -7954 -132551
rect -7910 -132595 -7854 -132551
rect -7810 -132595 -7354 -132551
rect -7310 -132595 -7254 -132551
rect -7210 -132595 -7154 -132551
rect -7110 -132595 -7054 -132551
rect -7010 -132595 -6954 -132551
rect -6910 -132595 -6854 -132551
rect -6810 -132595 -6754 -132551
rect -6710 -132595 -6654 -132551
rect -6610 -132595 -6554 -132551
rect -6510 -132595 -6454 -132551
rect -6410 -132595 -6354 -132551
rect -6310 -132595 -6254 -132551
rect -6210 -132595 -6154 -132551
rect -6110 -132595 -6054 -132551
rect -6010 -132595 -5954 -132551
rect -5910 -132595 -5854 -132551
rect -5810 -132585 177664 -132551
rect -5810 -132595 37387 -132585
rect -108812 -132629 37387 -132595
rect 37431 -132629 37487 -132585
rect 37531 -132629 37587 -132585
rect 37631 -132629 37687 -132585
rect 37731 -132629 37787 -132585
rect 37831 -132629 37887 -132585
rect 37931 -132629 37987 -132585
rect 38031 -132629 38087 -132585
rect 38131 -132629 38187 -132585
rect 38231 -132629 38287 -132585
rect 38331 -132629 38387 -132585
rect 38431 -132629 38487 -132585
rect 38531 -132629 38587 -132585
rect 38631 -132629 38687 -132585
rect 38731 -132629 38787 -132585
rect 38831 -132629 38887 -132585
rect 38931 -132629 39387 -132585
rect 39431 -132629 39487 -132585
rect 39531 -132629 39587 -132585
rect 39631 -132629 39687 -132585
rect 39731 -132629 39787 -132585
rect 39831 -132629 39887 -132585
rect 39931 -132629 39987 -132585
rect 40031 -132629 40087 -132585
rect 40131 -132629 40187 -132585
rect 40231 -132629 40287 -132585
rect 40331 -132629 40387 -132585
rect 40431 -132629 40487 -132585
rect 40531 -132629 40587 -132585
rect 40631 -132629 40687 -132585
rect 40731 -132629 40787 -132585
rect 40831 -132629 40887 -132585
rect 40931 -132629 41387 -132585
rect 41431 -132629 41487 -132585
rect 41531 -132629 41587 -132585
rect 41631 -132629 41687 -132585
rect 41731 -132629 41787 -132585
rect 41831 -132629 41887 -132585
rect 41931 -132629 41987 -132585
rect 42031 -132629 42087 -132585
rect 42131 -132629 42187 -132585
rect 42231 -132629 42287 -132585
rect 42331 -132629 42387 -132585
rect 42431 -132629 42487 -132585
rect 42531 -132629 42587 -132585
rect 42631 -132629 42687 -132585
rect 42731 -132629 42787 -132585
rect 42831 -132629 42887 -132585
rect 42931 -132629 43387 -132585
rect 43431 -132629 43487 -132585
rect 43531 -132629 43587 -132585
rect 43631 -132629 43687 -132585
rect 43731 -132629 43787 -132585
rect 43831 -132629 43887 -132585
rect 43931 -132629 43987 -132585
rect 44031 -132629 44087 -132585
rect 44131 -132629 44187 -132585
rect 44231 -132629 44287 -132585
rect 44331 -132629 44387 -132585
rect 44431 -132629 44487 -132585
rect 44531 -132629 44587 -132585
rect 44631 -132629 44687 -132585
rect 44731 -132629 44787 -132585
rect 44831 -132629 44887 -132585
rect 44931 -132629 177664 -132585
rect -108812 -132651 177664 -132629
rect -108812 -132695 -13354 -132651
rect -13310 -132695 -13254 -132651
rect -13210 -132695 -13154 -132651
rect -13110 -132695 -13054 -132651
rect -13010 -132695 -12954 -132651
rect -12910 -132695 -12854 -132651
rect -12810 -132695 -12754 -132651
rect -12710 -132695 -12654 -132651
rect -12610 -132695 -12554 -132651
rect -12510 -132695 -12454 -132651
rect -12410 -132695 -12354 -132651
rect -12310 -132695 -12254 -132651
rect -12210 -132695 -12154 -132651
rect -12110 -132695 -12054 -132651
rect -12010 -132695 -11954 -132651
rect -11910 -132695 -11854 -132651
rect -11810 -132695 -11354 -132651
rect -11310 -132695 -11254 -132651
rect -11210 -132695 -11154 -132651
rect -11110 -132695 -11054 -132651
rect -11010 -132695 -10954 -132651
rect -10910 -132695 -10854 -132651
rect -10810 -132695 -10754 -132651
rect -10710 -132695 -10654 -132651
rect -10610 -132695 -10554 -132651
rect -10510 -132695 -10454 -132651
rect -10410 -132695 -10354 -132651
rect -10310 -132695 -10254 -132651
rect -10210 -132695 -10154 -132651
rect -10110 -132695 -10054 -132651
rect -10010 -132695 -9954 -132651
rect -9910 -132695 -9854 -132651
rect -9810 -132695 -9354 -132651
rect -9310 -132695 -9254 -132651
rect -9210 -132695 -9154 -132651
rect -9110 -132695 -9054 -132651
rect -9010 -132695 -8954 -132651
rect -8910 -132695 -8854 -132651
rect -8810 -132695 -8754 -132651
rect -8710 -132695 -8654 -132651
rect -8610 -132695 -8554 -132651
rect -8510 -132695 -8454 -132651
rect -8410 -132695 -8354 -132651
rect -8310 -132695 -8254 -132651
rect -8210 -132695 -8154 -132651
rect -8110 -132695 -8054 -132651
rect -8010 -132695 -7954 -132651
rect -7910 -132695 -7854 -132651
rect -7810 -132695 -7354 -132651
rect -7310 -132695 -7254 -132651
rect -7210 -132695 -7154 -132651
rect -7110 -132695 -7054 -132651
rect -7010 -132695 -6954 -132651
rect -6910 -132695 -6854 -132651
rect -6810 -132695 -6754 -132651
rect -6710 -132695 -6654 -132651
rect -6610 -132695 -6554 -132651
rect -6510 -132695 -6454 -132651
rect -6410 -132695 -6354 -132651
rect -6310 -132695 -6254 -132651
rect -6210 -132695 -6154 -132651
rect -6110 -132695 -6054 -132651
rect -6010 -132695 -5954 -132651
rect -5910 -132695 -5854 -132651
rect -5810 -132685 177664 -132651
rect -5810 -132695 37387 -132685
rect -108812 -132729 37387 -132695
rect 37431 -132729 37487 -132685
rect 37531 -132729 37587 -132685
rect 37631 -132729 37687 -132685
rect 37731 -132729 37787 -132685
rect 37831 -132729 37887 -132685
rect 37931 -132729 37987 -132685
rect 38031 -132729 38087 -132685
rect 38131 -132729 38187 -132685
rect 38231 -132729 38287 -132685
rect 38331 -132729 38387 -132685
rect 38431 -132729 38487 -132685
rect 38531 -132729 38587 -132685
rect 38631 -132729 38687 -132685
rect 38731 -132729 38787 -132685
rect 38831 -132729 38887 -132685
rect 38931 -132729 39387 -132685
rect 39431 -132729 39487 -132685
rect 39531 -132729 39587 -132685
rect 39631 -132729 39687 -132685
rect 39731 -132729 39787 -132685
rect 39831 -132729 39887 -132685
rect 39931 -132729 39987 -132685
rect 40031 -132729 40087 -132685
rect 40131 -132729 40187 -132685
rect 40231 -132729 40287 -132685
rect 40331 -132729 40387 -132685
rect 40431 -132729 40487 -132685
rect 40531 -132729 40587 -132685
rect 40631 -132729 40687 -132685
rect 40731 -132729 40787 -132685
rect 40831 -132729 40887 -132685
rect 40931 -132729 41387 -132685
rect 41431 -132729 41487 -132685
rect 41531 -132729 41587 -132685
rect 41631 -132729 41687 -132685
rect 41731 -132729 41787 -132685
rect 41831 -132729 41887 -132685
rect 41931 -132729 41987 -132685
rect 42031 -132729 42087 -132685
rect 42131 -132729 42187 -132685
rect 42231 -132729 42287 -132685
rect 42331 -132729 42387 -132685
rect 42431 -132729 42487 -132685
rect 42531 -132729 42587 -132685
rect 42631 -132729 42687 -132685
rect 42731 -132729 42787 -132685
rect 42831 -132729 42887 -132685
rect 42931 -132729 43387 -132685
rect 43431 -132729 43487 -132685
rect 43531 -132729 43587 -132685
rect 43631 -132729 43687 -132685
rect 43731 -132729 43787 -132685
rect 43831 -132729 43887 -132685
rect 43931 -132729 43987 -132685
rect 44031 -132729 44087 -132685
rect 44131 -132729 44187 -132685
rect 44231 -132729 44287 -132685
rect 44331 -132729 44387 -132685
rect 44431 -132729 44487 -132685
rect 44531 -132729 44587 -132685
rect 44631 -132729 44687 -132685
rect 44731 -132729 44787 -132685
rect 44831 -132729 44887 -132685
rect 44931 -132729 177664 -132685
rect -108812 -132751 177664 -132729
rect -108812 -132795 -13354 -132751
rect -13310 -132795 -13254 -132751
rect -13210 -132795 -13154 -132751
rect -13110 -132795 -13054 -132751
rect -13010 -132795 -12954 -132751
rect -12910 -132795 -12854 -132751
rect -12810 -132795 -12754 -132751
rect -12710 -132795 -12654 -132751
rect -12610 -132795 -12554 -132751
rect -12510 -132795 -12454 -132751
rect -12410 -132795 -12354 -132751
rect -12310 -132795 -12254 -132751
rect -12210 -132795 -12154 -132751
rect -12110 -132795 -12054 -132751
rect -12010 -132795 -11954 -132751
rect -11910 -132795 -11854 -132751
rect -11810 -132795 -11354 -132751
rect -11310 -132795 -11254 -132751
rect -11210 -132795 -11154 -132751
rect -11110 -132795 -11054 -132751
rect -11010 -132795 -10954 -132751
rect -10910 -132795 -10854 -132751
rect -10810 -132795 -10754 -132751
rect -10710 -132795 -10654 -132751
rect -10610 -132795 -10554 -132751
rect -10510 -132795 -10454 -132751
rect -10410 -132795 -10354 -132751
rect -10310 -132795 -10254 -132751
rect -10210 -132795 -10154 -132751
rect -10110 -132795 -10054 -132751
rect -10010 -132795 -9954 -132751
rect -9910 -132795 -9854 -132751
rect -9810 -132795 -9354 -132751
rect -9310 -132795 -9254 -132751
rect -9210 -132795 -9154 -132751
rect -9110 -132795 -9054 -132751
rect -9010 -132795 -8954 -132751
rect -8910 -132795 -8854 -132751
rect -8810 -132795 -8754 -132751
rect -8710 -132795 -8654 -132751
rect -8610 -132795 -8554 -132751
rect -8510 -132795 -8454 -132751
rect -8410 -132795 -8354 -132751
rect -8310 -132795 -8254 -132751
rect -8210 -132795 -8154 -132751
rect -8110 -132795 -8054 -132751
rect -8010 -132795 -7954 -132751
rect -7910 -132795 -7854 -132751
rect -7810 -132795 -7354 -132751
rect -7310 -132795 -7254 -132751
rect -7210 -132795 -7154 -132751
rect -7110 -132795 -7054 -132751
rect -7010 -132795 -6954 -132751
rect -6910 -132795 -6854 -132751
rect -6810 -132795 -6754 -132751
rect -6710 -132795 -6654 -132751
rect -6610 -132795 -6554 -132751
rect -6510 -132795 -6454 -132751
rect -6410 -132795 -6354 -132751
rect -6310 -132795 -6254 -132751
rect -6210 -132795 -6154 -132751
rect -6110 -132795 -6054 -132751
rect -6010 -132795 -5954 -132751
rect -5910 -132795 -5854 -132751
rect -5810 -132785 177664 -132751
rect -5810 -132795 37387 -132785
rect -108812 -132829 37387 -132795
rect 37431 -132829 37487 -132785
rect 37531 -132829 37587 -132785
rect 37631 -132829 37687 -132785
rect 37731 -132829 37787 -132785
rect 37831 -132829 37887 -132785
rect 37931 -132829 37987 -132785
rect 38031 -132829 38087 -132785
rect 38131 -132829 38187 -132785
rect 38231 -132829 38287 -132785
rect 38331 -132829 38387 -132785
rect 38431 -132829 38487 -132785
rect 38531 -132829 38587 -132785
rect 38631 -132829 38687 -132785
rect 38731 -132829 38787 -132785
rect 38831 -132829 38887 -132785
rect 38931 -132829 39387 -132785
rect 39431 -132829 39487 -132785
rect 39531 -132829 39587 -132785
rect 39631 -132829 39687 -132785
rect 39731 -132829 39787 -132785
rect 39831 -132829 39887 -132785
rect 39931 -132829 39987 -132785
rect 40031 -132829 40087 -132785
rect 40131 -132829 40187 -132785
rect 40231 -132829 40287 -132785
rect 40331 -132829 40387 -132785
rect 40431 -132829 40487 -132785
rect 40531 -132829 40587 -132785
rect 40631 -132829 40687 -132785
rect 40731 -132829 40787 -132785
rect 40831 -132829 40887 -132785
rect 40931 -132829 41387 -132785
rect 41431 -132829 41487 -132785
rect 41531 -132829 41587 -132785
rect 41631 -132829 41687 -132785
rect 41731 -132829 41787 -132785
rect 41831 -132829 41887 -132785
rect 41931 -132829 41987 -132785
rect 42031 -132829 42087 -132785
rect 42131 -132829 42187 -132785
rect 42231 -132829 42287 -132785
rect 42331 -132829 42387 -132785
rect 42431 -132829 42487 -132785
rect 42531 -132829 42587 -132785
rect 42631 -132829 42687 -132785
rect 42731 -132829 42787 -132785
rect 42831 -132829 42887 -132785
rect 42931 -132829 43387 -132785
rect 43431 -132829 43487 -132785
rect 43531 -132829 43587 -132785
rect 43631 -132829 43687 -132785
rect 43731 -132829 43787 -132785
rect 43831 -132829 43887 -132785
rect 43931 -132829 43987 -132785
rect 44031 -132829 44087 -132785
rect 44131 -132829 44187 -132785
rect 44231 -132829 44287 -132785
rect 44331 -132829 44387 -132785
rect 44431 -132829 44487 -132785
rect 44531 -132829 44587 -132785
rect 44631 -132829 44687 -132785
rect 44731 -132829 44787 -132785
rect 44831 -132829 44887 -132785
rect 44931 -132829 177664 -132785
rect -108812 -132885 177664 -132829
rect -108812 -132929 37387 -132885
rect 37431 -132929 37487 -132885
rect 37531 -132929 37587 -132885
rect 37631 -132929 37687 -132885
rect 37731 -132929 37787 -132885
rect 37831 -132929 37887 -132885
rect 37931 -132929 37987 -132885
rect 38031 -132929 38087 -132885
rect 38131 -132929 38187 -132885
rect 38231 -132929 38287 -132885
rect 38331 -132929 38387 -132885
rect 38431 -132929 38487 -132885
rect 38531 -132929 38587 -132885
rect 38631 -132929 38687 -132885
rect 38731 -132929 38787 -132885
rect 38831 -132929 38887 -132885
rect 38931 -132929 39387 -132885
rect 39431 -132929 39487 -132885
rect 39531 -132929 39587 -132885
rect 39631 -132929 39687 -132885
rect 39731 -132929 39787 -132885
rect 39831 -132929 39887 -132885
rect 39931 -132929 39987 -132885
rect 40031 -132929 40087 -132885
rect 40131 -132929 40187 -132885
rect 40231 -132929 40287 -132885
rect 40331 -132929 40387 -132885
rect 40431 -132929 40487 -132885
rect 40531 -132929 40587 -132885
rect 40631 -132929 40687 -132885
rect 40731 -132929 40787 -132885
rect 40831 -132929 40887 -132885
rect 40931 -132929 41387 -132885
rect 41431 -132929 41487 -132885
rect 41531 -132929 41587 -132885
rect 41631 -132929 41687 -132885
rect 41731 -132929 41787 -132885
rect 41831 -132929 41887 -132885
rect 41931 -132929 41987 -132885
rect 42031 -132929 42087 -132885
rect 42131 -132929 42187 -132885
rect 42231 -132929 42287 -132885
rect 42331 -132929 42387 -132885
rect 42431 -132929 42487 -132885
rect 42531 -132929 42587 -132885
rect 42631 -132929 42687 -132885
rect 42731 -132929 42787 -132885
rect 42831 -132929 42887 -132885
rect 42931 -132929 43387 -132885
rect 43431 -132929 43487 -132885
rect 43531 -132929 43587 -132885
rect 43631 -132929 43687 -132885
rect 43731 -132929 43787 -132885
rect 43831 -132929 43887 -132885
rect 43931 -132929 43987 -132885
rect 44031 -132929 44087 -132885
rect 44131 -132929 44187 -132885
rect 44231 -132929 44287 -132885
rect 44331 -132929 44387 -132885
rect 44431 -132929 44487 -132885
rect 44531 -132929 44587 -132885
rect 44631 -132929 44687 -132885
rect 44731 -132929 44787 -132885
rect 44831 -132929 44887 -132885
rect 44931 -132929 177664 -132885
rect -108812 -133867 177664 -132929
rect -105360 -135314 -95895 -134569
rect -105360 -135358 -104783 -135314
rect -104739 -135358 -104683 -135314
rect -104639 -135358 -104583 -135314
rect -104539 -135358 -104483 -135314
rect -104439 -135358 -104383 -135314
rect -104339 -135358 -104283 -135314
rect -104239 -135358 -104183 -135314
rect -104139 -135358 -104083 -135314
rect -104039 -135358 -103983 -135314
rect -103939 -135358 -103883 -135314
rect -103839 -135358 -103783 -135314
rect -103739 -135358 -103683 -135314
rect -103639 -135358 -103583 -135314
rect -103539 -135358 -103483 -135314
rect -103439 -135358 -103383 -135314
rect -103339 -135358 -103283 -135314
rect -103239 -135358 -102783 -135314
rect -102739 -135358 -102683 -135314
rect -102639 -135358 -102583 -135314
rect -102539 -135358 -102483 -135314
rect -102439 -135358 -102383 -135314
rect -102339 -135358 -102283 -135314
rect -102239 -135358 -102183 -135314
rect -102139 -135358 -102083 -135314
rect -102039 -135358 -101983 -135314
rect -101939 -135358 -101883 -135314
rect -101839 -135358 -101783 -135314
rect -101739 -135358 -101683 -135314
rect -101639 -135358 -101583 -135314
rect -101539 -135358 -101483 -135314
rect -101439 -135358 -101383 -135314
rect -101339 -135358 -101283 -135314
rect -101239 -135358 -100783 -135314
rect -100739 -135358 -100683 -135314
rect -100639 -135358 -100583 -135314
rect -100539 -135358 -100483 -135314
rect -100439 -135358 -100383 -135314
rect -100339 -135358 -100283 -135314
rect -100239 -135358 -100183 -135314
rect -100139 -135358 -100083 -135314
rect -100039 -135358 -99983 -135314
rect -99939 -135358 -99883 -135314
rect -99839 -135358 -99783 -135314
rect -99739 -135358 -99683 -135314
rect -99639 -135358 -99583 -135314
rect -99539 -135358 -99483 -135314
rect -99439 -135358 -99383 -135314
rect -99339 -135358 -99283 -135314
rect -99239 -135358 -98783 -135314
rect -98739 -135358 -98683 -135314
rect -98639 -135358 -98583 -135314
rect -98539 -135358 -98483 -135314
rect -98439 -135358 -98383 -135314
rect -98339 -135358 -98283 -135314
rect -98239 -135358 -98183 -135314
rect -98139 -135358 -98083 -135314
rect -98039 -135358 -97983 -135314
rect -97939 -135358 -97883 -135314
rect -97839 -135358 -97783 -135314
rect -97739 -135358 -97683 -135314
rect -97639 -135358 -97583 -135314
rect -97539 -135358 -97483 -135314
rect -97439 -135358 -97383 -135314
rect -97339 -135358 -97283 -135314
rect -97239 -135358 -95895 -135314
rect -105360 -135414 -95895 -135358
rect -105360 -135458 -104783 -135414
rect -104739 -135458 -104683 -135414
rect -104639 -135458 -104583 -135414
rect -104539 -135458 -104483 -135414
rect -104439 -135458 -104383 -135414
rect -104339 -135458 -104283 -135414
rect -104239 -135458 -104183 -135414
rect -104139 -135458 -104083 -135414
rect -104039 -135458 -103983 -135414
rect -103939 -135458 -103883 -135414
rect -103839 -135458 -103783 -135414
rect -103739 -135458 -103683 -135414
rect -103639 -135458 -103583 -135414
rect -103539 -135458 -103483 -135414
rect -103439 -135458 -103383 -135414
rect -103339 -135458 -103283 -135414
rect -103239 -135458 -102783 -135414
rect -102739 -135458 -102683 -135414
rect -102639 -135458 -102583 -135414
rect -102539 -135458 -102483 -135414
rect -102439 -135458 -102383 -135414
rect -102339 -135458 -102283 -135414
rect -102239 -135458 -102183 -135414
rect -102139 -135458 -102083 -135414
rect -102039 -135458 -101983 -135414
rect -101939 -135458 -101883 -135414
rect -101839 -135458 -101783 -135414
rect -101739 -135458 -101683 -135414
rect -101639 -135458 -101583 -135414
rect -101539 -135458 -101483 -135414
rect -101439 -135458 -101383 -135414
rect -101339 -135458 -101283 -135414
rect -101239 -135458 -100783 -135414
rect -100739 -135458 -100683 -135414
rect -100639 -135458 -100583 -135414
rect -100539 -135458 -100483 -135414
rect -100439 -135458 -100383 -135414
rect -100339 -135458 -100283 -135414
rect -100239 -135458 -100183 -135414
rect -100139 -135458 -100083 -135414
rect -100039 -135458 -99983 -135414
rect -99939 -135458 -99883 -135414
rect -99839 -135458 -99783 -135414
rect -99739 -135458 -99683 -135414
rect -99639 -135458 -99583 -135414
rect -99539 -135458 -99483 -135414
rect -99439 -135458 -99383 -135414
rect -99339 -135458 -99283 -135414
rect -99239 -135458 -98783 -135414
rect -98739 -135458 -98683 -135414
rect -98639 -135458 -98583 -135414
rect -98539 -135458 -98483 -135414
rect -98439 -135458 -98383 -135414
rect -98339 -135458 -98283 -135414
rect -98239 -135458 -98183 -135414
rect -98139 -135458 -98083 -135414
rect -98039 -135458 -97983 -135414
rect -97939 -135458 -97883 -135414
rect -97839 -135458 -97783 -135414
rect -97739 -135458 -97683 -135414
rect -97639 -135458 -97583 -135414
rect -97539 -135458 -97483 -135414
rect -97439 -135458 -97383 -135414
rect -97339 -135458 -97283 -135414
rect -97239 -135458 -95895 -135414
rect -105360 -135514 -95895 -135458
rect -105360 -135558 -104783 -135514
rect -104739 -135558 -104683 -135514
rect -104639 -135558 -104583 -135514
rect -104539 -135558 -104483 -135514
rect -104439 -135558 -104383 -135514
rect -104339 -135558 -104283 -135514
rect -104239 -135558 -104183 -135514
rect -104139 -135558 -104083 -135514
rect -104039 -135558 -103983 -135514
rect -103939 -135558 -103883 -135514
rect -103839 -135558 -103783 -135514
rect -103739 -135558 -103683 -135514
rect -103639 -135558 -103583 -135514
rect -103539 -135558 -103483 -135514
rect -103439 -135558 -103383 -135514
rect -103339 -135558 -103283 -135514
rect -103239 -135558 -102783 -135514
rect -102739 -135558 -102683 -135514
rect -102639 -135558 -102583 -135514
rect -102539 -135558 -102483 -135514
rect -102439 -135558 -102383 -135514
rect -102339 -135558 -102283 -135514
rect -102239 -135558 -102183 -135514
rect -102139 -135558 -102083 -135514
rect -102039 -135558 -101983 -135514
rect -101939 -135558 -101883 -135514
rect -101839 -135558 -101783 -135514
rect -101739 -135558 -101683 -135514
rect -101639 -135558 -101583 -135514
rect -101539 -135558 -101483 -135514
rect -101439 -135558 -101383 -135514
rect -101339 -135558 -101283 -135514
rect -101239 -135558 -100783 -135514
rect -100739 -135558 -100683 -135514
rect -100639 -135558 -100583 -135514
rect -100539 -135558 -100483 -135514
rect -100439 -135558 -100383 -135514
rect -100339 -135558 -100283 -135514
rect -100239 -135558 -100183 -135514
rect -100139 -135558 -100083 -135514
rect -100039 -135558 -99983 -135514
rect -99939 -135558 -99883 -135514
rect -99839 -135558 -99783 -135514
rect -99739 -135558 -99683 -135514
rect -99639 -135558 -99583 -135514
rect -99539 -135558 -99483 -135514
rect -99439 -135558 -99383 -135514
rect -99339 -135558 -99283 -135514
rect -99239 -135558 -98783 -135514
rect -98739 -135558 -98683 -135514
rect -98639 -135558 -98583 -135514
rect -98539 -135558 -98483 -135514
rect -98439 -135558 -98383 -135514
rect -98339 -135558 -98283 -135514
rect -98239 -135558 -98183 -135514
rect -98139 -135558 -98083 -135514
rect -98039 -135558 -97983 -135514
rect -97939 -135558 -97883 -135514
rect -97839 -135558 -97783 -135514
rect -97739 -135558 -97683 -135514
rect -97639 -135558 -97583 -135514
rect -97539 -135558 -97483 -135514
rect -97439 -135558 -97383 -135514
rect -97339 -135558 -97283 -135514
rect -97239 -135558 -95895 -135514
rect -105360 -135614 -95895 -135558
rect -105360 -135658 -104783 -135614
rect -104739 -135658 -104683 -135614
rect -104639 -135658 -104583 -135614
rect -104539 -135658 -104483 -135614
rect -104439 -135658 -104383 -135614
rect -104339 -135658 -104283 -135614
rect -104239 -135658 -104183 -135614
rect -104139 -135658 -104083 -135614
rect -104039 -135658 -103983 -135614
rect -103939 -135658 -103883 -135614
rect -103839 -135658 -103783 -135614
rect -103739 -135658 -103683 -135614
rect -103639 -135658 -103583 -135614
rect -103539 -135658 -103483 -135614
rect -103439 -135658 -103383 -135614
rect -103339 -135658 -103283 -135614
rect -103239 -135658 -102783 -135614
rect -102739 -135658 -102683 -135614
rect -102639 -135658 -102583 -135614
rect -102539 -135658 -102483 -135614
rect -102439 -135658 -102383 -135614
rect -102339 -135658 -102283 -135614
rect -102239 -135658 -102183 -135614
rect -102139 -135658 -102083 -135614
rect -102039 -135658 -101983 -135614
rect -101939 -135658 -101883 -135614
rect -101839 -135658 -101783 -135614
rect -101739 -135658 -101683 -135614
rect -101639 -135658 -101583 -135614
rect -101539 -135658 -101483 -135614
rect -101439 -135658 -101383 -135614
rect -101339 -135658 -101283 -135614
rect -101239 -135658 -100783 -135614
rect -100739 -135658 -100683 -135614
rect -100639 -135658 -100583 -135614
rect -100539 -135658 -100483 -135614
rect -100439 -135658 -100383 -135614
rect -100339 -135658 -100283 -135614
rect -100239 -135658 -100183 -135614
rect -100139 -135658 -100083 -135614
rect -100039 -135658 -99983 -135614
rect -99939 -135658 -99883 -135614
rect -99839 -135658 -99783 -135614
rect -99739 -135658 -99683 -135614
rect -99639 -135658 -99583 -135614
rect -99539 -135658 -99483 -135614
rect -99439 -135658 -99383 -135614
rect -99339 -135658 -99283 -135614
rect -99239 -135658 -98783 -135614
rect -98739 -135658 -98683 -135614
rect -98639 -135658 -98583 -135614
rect -98539 -135658 -98483 -135614
rect -98439 -135658 -98383 -135614
rect -98339 -135658 -98283 -135614
rect -98239 -135658 -98183 -135614
rect -98139 -135658 -98083 -135614
rect -98039 -135658 -97983 -135614
rect -97939 -135658 -97883 -135614
rect -97839 -135658 -97783 -135614
rect -97739 -135658 -97683 -135614
rect -97639 -135658 -97583 -135614
rect -97539 -135658 -97483 -135614
rect -97439 -135658 -97383 -135614
rect -97339 -135658 -97283 -135614
rect -97239 -135658 -95895 -135614
rect -105360 -135714 -95895 -135658
rect -105360 -135758 -104783 -135714
rect -104739 -135758 -104683 -135714
rect -104639 -135758 -104583 -135714
rect -104539 -135758 -104483 -135714
rect -104439 -135758 -104383 -135714
rect -104339 -135758 -104283 -135714
rect -104239 -135758 -104183 -135714
rect -104139 -135758 -104083 -135714
rect -104039 -135758 -103983 -135714
rect -103939 -135758 -103883 -135714
rect -103839 -135758 -103783 -135714
rect -103739 -135758 -103683 -135714
rect -103639 -135758 -103583 -135714
rect -103539 -135758 -103483 -135714
rect -103439 -135758 -103383 -135714
rect -103339 -135758 -103283 -135714
rect -103239 -135758 -102783 -135714
rect -102739 -135758 -102683 -135714
rect -102639 -135758 -102583 -135714
rect -102539 -135758 -102483 -135714
rect -102439 -135758 -102383 -135714
rect -102339 -135758 -102283 -135714
rect -102239 -135758 -102183 -135714
rect -102139 -135758 -102083 -135714
rect -102039 -135758 -101983 -135714
rect -101939 -135758 -101883 -135714
rect -101839 -135758 -101783 -135714
rect -101739 -135758 -101683 -135714
rect -101639 -135758 -101583 -135714
rect -101539 -135758 -101483 -135714
rect -101439 -135758 -101383 -135714
rect -101339 -135758 -101283 -135714
rect -101239 -135758 -100783 -135714
rect -100739 -135758 -100683 -135714
rect -100639 -135758 -100583 -135714
rect -100539 -135758 -100483 -135714
rect -100439 -135758 -100383 -135714
rect -100339 -135758 -100283 -135714
rect -100239 -135758 -100183 -135714
rect -100139 -135758 -100083 -135714
rect -100039 -135758 -99983 -135714
rect -99939 -135758 -99883 -135714
rect -99839 -135758 -99783 -135714
rect -99739 -135758 -99683 -135714
rect -99639 -135758 -99583 -135714
rect -99539 -135758 -99483 -135714
rect -99439 -135758 -99383 -135714
rect -99339 -135758 -99283 -135714
rect -99239 -135758 -98783 -135714
rect -98739 -135758 -98683 -135714
rect -98639 -135758 -98583 -135714
rect -98539 -135758 -98483 -135714
rect -98439 -135758 -98383 -135714
rect -98339 -135758 -98283 -135714
rect -98239 -135758 -98183 -135714
rect -98139 -135758 -98083 -135714
rect -98039 -135758 -97983 -135714
rect -97939 -135758 -97883 -135714
rect -97839 -135758 -97783 -135714
rect -97739 -135758 -97683 -135714
rect -97639 -135758 -97583 -135714
rect -97539 -135758 -97483 -135714
rect -97439 -135758 -97383 -135714
rect -97339 -135758 -97283 -135714
rect -97239 -135758 -95895 -135714
rect -105360 -135814 -95895 -135758
rect -105360 -135858 -104783 -135814
rect -104739 -135858 -104683 -135814
rect -104639 -135858 -104583 -135814
rect -104539 -135858 -104483 -135814
rect -104439 -135858 -104383 -135814
rect -104339 -135858 -104283 -135814
rect -104239 -135858 -104183 -135814
rect -104139 -135858 -104083 -135814
rect -104039 -135858 -103983 -135814
rect -103939 -135858 -103883 -135814
rect -103839 -135858 -103783 -135814
rect -103739 -135858 -103683 -135814
rect -103639 -135858 -103583 -135814
rect -103539 -135858 -103483 -135814
rect -103439 -135858 -103383 -135814
rect -103339 -135858 -103283 -135814
rect -103239 -135858 -102783 -135814
rect -102739 -135858 -102683 -135814
rect -102639 -135858 -102583 -135814
rect -102539 -135858 -102483 -135814
rect -102439 -135858 -102383 -135814
rect -102339 -135858 -102283 -135814
rect -102239 -135858 -102183 -135814
rect -102139 -135858 -102083 -135814
rect -102039 -135858 -101983 -135814
rect -101939 -135858 -101883 -135814
rect -101839 -135858 -101783 -135814
rect -101739 -135858 -101683 -135814
rect -101639 -135858 -101583 -135814
rect -101539 -135858 -101483 -135814
rect -101439 -135858 -101383 -135814
rect -101339 -135858 -101283 -135814
rect -101239 -135858 -100783 -135814
rect -100739 -135858 -100683 -135814
rect -100639 -135858 -100583 -135814
rect -100539 -135858 -100483 -135814
rect -100439 -135858 -100383 -135814
rect -100339 -135858 -100283 -135814
rect -100239 -135858 -100183 -135814
rect -100139 -135858 -100083 -135814
rect -100039 -135858 -99983 -135814
rect -99939 -135858 -99883 -135814
rect -99839 -135858 -99783 -135814
rect -99739 -135858 -99683 -135814
rect -99639 -135858 -99583 -135814
rect -99539 -135858 -99483 -135814
rect -99439 -135858 -99383 -135814
rect -99339 -135858 -99283 -135814
rect -99239 -135858 -98783 -135814
rect -98739 -135858 -98683 -135814
rect -98639 -135858 -98583 -135814
rect -98539 -135858 -98483 -135814
rect -98439 -135858 -98383 -135814
rect -98339 -135858 -98283 -135814
rect -98239 -135858 -98183 -135814
rect -98139 -135858 -98083 -135814
rect -98039 -135858 -97983 -135814
rect -97939 -135858 -97883 -135814
rect -97839 -135858 -97783 -135814
rect -97739 -135858 -97683 -135814
rect -97639 -135858 -97583 -135814
rect -97539 -135858 -97483 -135814
rect -97439 -135858 -97383 -135814
rect -97339 -135858 -97283 -135814
rect -97239 -135858 -95895 -135814
rect -105360 -135914 -95895 -135858
rect -105360 -135958 -104783 -135914
rect -104739 -135958 -104683 -135914
rect -104639 -135958 -104583 -135914
rect -104539 -135958 -104483 -135914
rect -104439 -135958 -104383 -135914
rect -104339 -135958 -104283 -135914
rect -104239 -135958 -104183 -135914
rect -104139 -135958 -104083 -135914
rect -104039 -135958 -103983 -135914
rect -103939 -135958 -103883 -135914
rect -103839 -135958 -103783 -135914
rect -103739 -135958 -103683 -135914
rect -103639 -135958 -103583 -135914
rect -103539 -135958 -103483 -135914
rect -103439 -135958 -103383 -135914
rect -103339 -135958 -103283 -135914
rect -103239 -135958 -102783 -135914
rect -102739 -135958 -102683 -135914
rect -102639 -135958 -102583 -135914
rect -102539 -135958 -102483 -135914
rect -102439 -135958 -102383 -135914
rect -102339 -135958 -102283 -135914
rect -102239 -135958 -102183 -135914
rect -102139 -135958 -102083 -135914
rect -102039 -135958 -101983 -135914
rect -101939 -135958 -101883 -135914
rect -101839 -135958 -101783 -135914
rect -101739 -135958 -101683 -135914
rect -101639 -135958 -101583 -135914
rect -101539 -135958 -101483 -135914
rect -101439 -135958 -101383 -135914
rect -101339 -135958 -101283 -135914
rect -101239 -135958 -100783 -135914
rect -100739 -135958 -100683 -135914
rect -100639 -135958 -100583 -135914
rect -100539 -135958 -100483 -135914
rect -100439 -135958 -100383 -135914
rect -100339 -135958 -100283 -135914
rect -100239 -135958 -100183 -135914
rect -100139 -135958 -100083 -135914
rect -100039 -135958 -99983 -135914
rect -99939 -135958 -99883 -135914
rect -99839 -135958 -99783 -135914
rect -99739 -135958 -99683 -135914
rect -99639 -135958 -99583 -135914
rect -99539 -135958 -99483 -135914
rect -99439 -135958 -99383 -135914
rect -99339 -135958 -99283 -135914
rect -99239 -135958 -98783 -135914
rect -98739 -135958 -98683 -135914
rect -98639 -135958 -98583 -135914
rect -98539 -135958 -98483 -135914
rect -98439 -135958 -98383 -135914
rect -98339 -135958 -98283 -135914
rect -98239 -135958 -98183 -135914
rect -98139 -135958 -98083 -135914
rect -98039 -135958 -97983 -135914
rect -97939 -135958 -97883 -135914
rect -97839 -135958 -97783 -135914
rect -97739 -135958 -97683 -135914
rect -97639 -135958 -97583 -135914
rect -97539 -135958 -97483 -135914
rect -97439 -135958 -97383 -135914
rect -97339 -135958 -97283 -135914
rect -97239 -135958 -95895 -135914
rect -105360 -136014 -95895 -135958
rect -105360 -136058 -104783 -136014
rect -104739 -136058 -104683 -136014
rect -104639 -136058 -104583 -136014
rect -104539 -136058 -104483 -136014
rect -104439 -136058 -104383 -136014
rect -104339 -136058 -104283 -136014
rect -104239 -136058 -104183 -136014
rect -104139 -136058 -104083 -136014
rect -104039 -136058 -103983 -136014
rect -103939 -136058 -103883 -136014
rect -103839 -136058 -103783 -136014
rect -103739 -136058 -103683 -136014
rect -103639 -136058 -103583 -136014
rect -103539 -136058 -103483 -136014
rect -103439 -136058 -103383 -136014
rect -103339 -136058 -103283 -136014
rect -103239 -136058 -102783 -136014
rect -102739 -136058 -102683 -136014
rect -102639 -136058 -102583 -136014
rect -102539 -136058 -102483 -136014
rect -102439 -136058 -102383 -136014
rect -102339 -136058 -102283 -136014
rect -102239 -136058 -102183 -136014
rect -102139 -136058 -102083 -136014
rect -102039 -136058 -101983 -136014
rect -101939 -136058 -101883 -136014
rect -101839 -136058 -101783 -136014
rect -101739 -136058 -101683 -136014
rect -101639 -136058 -101583 -136014
rect -101539 -136058 -101483 -136014
rect -101439 -136058 -101383 -136014
rect -101339 -136058 -101283 -136014
rect -101239 -136058 -100783 -136014
rect -100739 -136058 -100683 -136014
rect -100639 -136058 -100583 -136014
rect -100539 -136058 -100483 -136014
rect -100439 -136058 -100383 -136014
rect -100339 -136058 -100283 -136014
rect -100239 -136058 -100183 -136014
rect -100139 -136058 -100083 -136014
rect -100039 -136058 -99983 -136014
rect -99939 -136058 -99883 -136014
rect -99839 -136058 -99783 -136014
rect -99739 -136058 -99683 -136014
rect -99639 -136058 -99583 -136014
rect -99539 -136058 -99483 -136014
rect -99439 -136058 -99383 -136014
rect -99339 -136058 -99283 -136014
rect -99239 -136058 -98783 -136014
rect -98739 -136058 -98683 -136014
rect -98639 -136058 -98583 -136014
rect -98539 -136058 -98483 -136014
rect -98439 -136058 -98383 -136014
rect -98339 -136058 -98283 -136014
rect -98239 -136058 -98183 -136014
rect -98139 -136058 -98083 -136014
rect -98039 -136058 -97983 -136014
rect -97939 -136058 -97883 -136014
rect -97839 -136058 -97783 -136014
rect -97739 -136058 -97683 -136014
rect -97639 -136058 -97583 -136014
rect -97539 -136058 -97483 -136014
rect -97439 -136058 -97383 -136014
rect -97339 -136058 -97283 -136014
rect -97239 -136058 -95895 -136014
rect -105360 -136114 -95895 -136058
rect -105360 -136158 -104783 -136114
rect -104739 -136158 -104683 -136114
rect -104639 -136158 -104583 -136114
rect -104539 -136158 -104483 -136114
rect -104439 -136158 -104383 -136114
rect -104339 -136158 -104283 -136114
rect -104239 -136158 -104183 -136114
rect -104139 -136158 -104083 -136114
rect -104039 -136158 -103983 -136114
rect -103939 -136158 -103883 -136114
rect -103839 -136158 -103783 -136114
rect -103739 -136158 -103683 -136114
rect -103639 -136158 -103583 -136114
rect -103539 -136158 -103483 -136114
rect -103439 -136158 -103383 -136114
rect -103339 -136158 -103283 -136114
rect -103239 -136158 -102783 -136114
rect -102739 -136158 -102683 -136114
rect -102639 -136158 -102583 -136114
rect -102539 -136158 -102483 -136114
rect -102439 -136158 -102383 -136114
rect -102339 -136158 -102283 -136114
rect -102239 -136158 -102183 -136114
rect -102139 -136158 -102083 -136114
rect -102039 -136158 -101983 -136114
rect -101939 -136158 -101883 -136114
rect -101839 -136158 -101783 -136114
rect -101739 -136158 -101683 -136114
rect -101639 -136158 -101583 -136114
rect -101539 -136158 -101483 -136114
rect -101439 -136158 -101383 -136114
rect -101339 -136158 -101283 -136114
rect -101239 -136158 -100783 -136114
rect -100739 -136158 -100683 -136114
rect -100639 -136158 -100583 -136114
rect -100539 -136158 -100483 -136114
rect -100439 -136158 -100383 -136114
rect -100339 -136158 -100283 -136114
rect -100239 -136158 -100183 -136114
rect -100139 -136158 -100083 -136114
rect -100039 -136158 -99983 -136114
rect -99939 -136158 -99883 -136114
rect -99839 -136158 -99783 -136114
rect -99739 -136158 -99683 -136114
rect -99639 -136158 -99583 -136114
rect -99539 -136158 -99483 -136114
rect -99439 -136158 -99383 -136114
rect -99339 -136158 -99283 -136114
rect -99239 -136158 -98783 -136114
rect -98739 -136158 -98683 -136114
rect -98639 -136158 -98583 -136114
rect -98539 -136158 -98483 -136114
rect -98439 -136158 -98383 -136114
rect -98339 -136158 -98283 -136114
rect -98239 -136158 -98183 -136114
rect -98139 -136158 -98083 -136114
rect -98039 -136158 -97983 -136114
rect -97939 -136158 -97883 -136114
rect -97839 -136158 -97783 -136114
rect -97739 -136158 -97683 -136114
rect -97639 -136158 -97583 -136114
rect -97539 -136158 -97483 -136114
rect -97439 -136158 -97383 -136114
rect -97339 -136158 -97283 -136114
rect -97239 -136158 -95895 -136114
rect -105360 -136214 -95895 -136158
rect -105360 -136258 -104783 -136214
rect -104739 -136258 -104683 -136214
rect -104639 -136258 -104583 -136214
rect -104539 -136258 -104483 -136214
rect -104439 -136258 -104383 -136214
rect -104339 -136258 -104283 -136214
rect -104239 -136258 -104183 -136214
rect -104139 -136258 -104083 -136214
rect -104039 -136258 -103983 -136214
rect -103939 -136258 -103883 -136214
rect -103839 -136258 -103783 -136214
rect -103739 -136258 -103683 -136214
rect -103639 -136258 -103583 -136214
rect -103539 -136258 -103483 -136214
rect -103439 -136258 -103383 -136214
rect -103339 -136258 -103283 -136214
rect -103239 -136258 -102783 -136214
rect -102739 -136258 -102683 -136214
rect -102639 -136258 -102583 -136214
rect -102539 -136258 -102483 -136214
rect -102439 -136258 -102383 -136214
rect -102339 -136258 -102283 -136214
rect -102239 -136258 -102183 -136214
rect -102139 -136258 -102083 -136214
rect -102039 -136258 -101983 -136214
rect -101939 -136258 -101883 -136214
rect -101839 -136258 -101783 -136214
rect -101739 -136258 -101683 -136214
rect -101639 -136258 -101583 -136214
rect -101539 -136258 -101483 -136214
rect -101439 -136258 -101383 -136214
rect -101339 -136258 -101283 -136214
rect -101239 -136258 -100783 -136214
rect -100739 -136258 -100683 -136214
rect -100639 -136258 -100583 -136214
rect -100539 -136258 -100483 -136214
rect -100439 -136258 -100383 -136214
rect -100339 -136258 -100283 -136214
rect -100239 -136258 -100183 -136214
rect -100139 -136258 -100083 -136214
rect -100039 -136258 -99983 -136214
rect -99939 -136258 -99883 -136214
rect -99839 -136258 -99783 -136214
rect -99739 -136258 -99683 -136214
rect -99639 -136258 -99583 -136214
rect -99539 -136258 -99483 -136214
rect -99439 -136258 -99383 -136214
rect -99339 -136258 -99283 -136214
rect -99239 -136258 -98783 -136214
rect -98739 -136258 -98683 -136214
rect -98639 -136258 -98583 -136214
rect -98539 -136258 -98483 -136214
rect -98439 -136258 -98383 -136214
rect -98339 -136258 -98283 -136214
rect -98239 -136258 -98183 -136214
rect -98139 -136258 -98083 -136214
rect -98039 -136258 -97983 -136214
rect -97939 -136258 -97883 -136214
rect -97839 -136258 -97783 -136214
rect -97739 -136258 -97683 -136214
rect -97639 -136258 -97583 -136214
rect -97539 -136258 -97483 -136214
rect -97439 -136258 -97383 -136214
rect -97339 -136258 -97283 -136214
rect -97239 -136258 -95895 -136214
rect -105360 -136314 -95895 -136258
rect -105360 -136358 -104783 -136314
rect -104739 -136358 -104683 -136314
rect -104639 -136358 -104583 -136314
rect -104539 -136358 -104483 -136314
rect -104439 -136358 -104383 -136314
rect -104339 -136358 -104283 -136314
rect -104239 -136358 -104183 -136314
rect -104139 -136358 -104083 -136314
rect -104039 -136358 -103983 -136314
rect -103939 -136358 -103883 -136314
rect -103839 -136358 -103783 -136314
rect -103739 -136358 -103683 -136314
rect -103639 -136358 -103583 -136314
rect -103539 -136358 -103483 -136314
rect -103439 -136358 -103383 -136314
rect -103339 -136358 -103283 -136314
rect -103239 -136358 -102783 -136314
rect -102739 -136358 -102683 -136314
rect -102639 -136358 -102583 -136314
rect -102539 -136358 -102483 -136314
rect -102439 -136358 -102383 -136314
rect -102339 -136358 -102283 -136314
rect -102239 -136358 -102183 -136314
rect -102139 -136358 -102083 -136314
rect -102039 -136358 -101983 -136314
rect -101939 -136358 -101883 -136314
rect -101839 -136358 -101783 -136314
rect -101739 -136358 -101683 -136314
rect -101639 -136358 -101583 -136314
rect -101539 -136358 -101483 -136314
rect -101439 -136358 -101383 -136314
rect -101339 -136358 -101283 -136314
rect -101239 -136358 -100783 -136314
rect -100739 -136358 -100683 -136314
rect -100639 -136358 -100583 -136314
rect -100539 -136358 -100483 -136314
rect -100439 -136358 -100383 -136314
rect -100339 -136358 -100283 -136314
rect -100239 -136358 -100183 -136314
rect -100139 -136358 -100083 -136314
rect -100039 -136358 -99983 -136314
rect -99939 -136358 -99883 -136314
rect -99839 -136358 -99783 -136314
rect -99739 -136358 -99683 -136314
rect -99639 -136358 -99583 -136314
rect -99539 -136358 -99483 -136314
rect -99439 -136358 -99383 -136314
rect -99339 -136358 -99283 -136314
rect -99239 -136358 -98783 -136314
rect -98739 -136358 -98683 -136314
rect -98639 -136358 -98583 -136314
rect -98539 -136358 -98483 -136314
rect -98439 -136358 -98383 -136314
rect -98339 -136358 -98283 -136314
rect -98239 -136358 -98183 -136314
rect -98139 -136358 -98083 -136314
rect -98039 -136358 -97983 -136314
rect -97939 -136358 -97883 -136314
rect -97839 -136358 -97783 -136314
rect -97739 -136358 -97683 -136314
rect -97639 -136358 -97583 -136314
rect -97539 -136358 -97483 -136314
rect -97439 -136358 -97383 -136314
rect -97339 -136358 -97283 -136314
rect -97239 -136358 -95895 -136314
rect -105360 -136414 -95895 -136358
rect -105360 -136458 -104783 -136414
rect -104739 -136458 -104683 -136414
rect -104639 -136458 -104583 -136414
rect -104539 -136458 -104483 -136414
rect -104439 -136458 -104383 -136414
rect -104339 -136458 -104283 -136414
rect -104239 -136458 -104183 -136414
rect -104139 -136458 -104083 -136414
rect -104039 -136458 -103983 -136414
rect -103939 -136458 -103883 -136414
rect -103839 -136458 -103783 -136414
rect -103739 -136458 -103683 -136414
rect -103639 -136458 -103583 -136414
rect -103539 -136458 -103483 -136414
rect -103439 -136458 -103383 -136414
rect -103339 -136458 -103283 -136414
rect -103239 -136458 -102783 -136414
rect -102739 -136458 -102683 -136414
rect -102639 -136458 -102583 -136414
rect -102539 -136458 -102483 -136414
rect -102439 -136458 -102383 -136414
rect -102339 -136458 -102283 -136414
rect -102239 -136458 -102183 -136414
rect -102139 -136458 -102083 -136414
rect -102039 -136458 -101983 -136414
rect -101939 -136458 -101883 -136414
rect -101839 -136458 -101783 -136414
rect -101739 -136458 -101683 -136414
rect -101639 -136458 -101583 -136414
rect -101539 -136458 -101483 -136414
rect -101439 -136458 -101383 -136414
rect -101339 -136458 -101283 -136414
rect -101239 -136458 -100783 -136414
rect -100739 -136458 -100683 -136414
rect -100639 -136458 -100583 -136414
rect -100539 -136458 -100483 -136414
rect -100439 -136458 -100383 -136414
rect -100339 -136458 -100283 -136414
rect -100239 -136458 -100183 -136414
rect -100139 -136458 -100083 -136414
rect -100039 -136458 -99983 -136414
rect -99939 -136458 -99883 -136414
rect -99839 -136458 -99783 -136414
rect -99739 -136458 -99683 -136414
rect -99639 -136458 -99583 -136414
rect -99539 -136458 -99483 -136414
rect -99439 -136458 -99383 -136414
rect -99339 -136458 -99283 -136414
rect -99239 -136458 -98783 -136414
rect -98739 -136458 -98683 -136414
rect -98639 -136458 -98583 -136414
rect -98539 -136458 -98483 -136414
rect -98439 -136458 -98383 -136414
rect -98339 -136458 -98283 -136414
rect -98239 -136458 -98183 -136414
rect -98139 -136458 -98083 -136414
rect -98039 -136458 -97983 -136414
rect -97939 -136458 -97883 -136414
rect -97839 -136458 -97783 -136414
rect -97739 -136458 -97683 -136414
rect -97639 -136458 -97583 -136414
rect -97539 -136458 -97483 -136414
rect -97439 -136458 -97383 -136414
rect -97339 -136458 -97283 -136414
rect -97239 -136458 -95895 -136414
rect -105360 -136514 -95895 -136458
rect -105360 -136558 -104783 -136514
rect -104739 -136558 -104683 -136514
rect -104639 -136558 -104583 -136514
rect -104539 -136558 -104483 -136514
rect -104439 -136558 -104383 -136514
rect -104339 -136558 -104283 -136514
rect -104239 -136558 -104183 -136514
rect -104139 -136558 -104083 -136514
rect -104039 -136558 -103983 -136514
rect -103939 -136558 -103883 -136514
rect -103839 -136558 -103783 -136514
rect -103739 -136558 -103683 -136514
rect -103639 -136558 -103583 -136514
rect -103539 -136558 -103483 -136514
rect -103439 -136558 -103383 -136514
rect -103339 -136558 -103283 -136514
rect -103239 -136558 -102783 -136514
rect -102739 -136558 -102683 -136514
rect -102639 -136558 -102583 -136514
rect -102539 -136558 -102483 -136514
rect -102439 -136558 -102383 -136514
rect -102339 -136558 -102283 -136514
rect -102239 -136558 -102183 -136514
rect -102139 -136558 -102083 -136514
rect -102039 -136558 -101983 -136514
rect -101939 -136558 -101883 -136514
rect -101839 -136558 -101783 -136514
rect -101739 -136558 -101683 -136514
rect -101639 -136558 -101583 -136514
rect -101539 -136558 -101483 -136514
rect -101439 -136558 -101383 -136514
rect -101339 -136558 -101283 -136514
rect -101239 -136558 -100783 -136514
rect -100739 -136558 -100683 -136514
rect -100639 -136558 -100583 -136514
rect -100539 -136558 -100483 -136514
rect -100439 -136558 -100383 -136514
rect -100339 -136558 -100283 -136514
rect -100239 -136558 -100183 -136514
rect -100139 -136558 -100083 -136514
rect -100039 -136558 -99983 -136514
rect -99939 -136558 -99883 -136514
rect -99839 -136558 -99783 -136514
rect -99739 -136558 -99683 -136514
rect -99639 -136558 -99583 -136514
rect -99539 -136558 -99483 -136514
rect -99439 -136558 -99383 -136514
rect -99339 -136558 -99283 -136514
rect -99239 -136558 -98783 -136514
rect -98739 -136558 -98683 -136514
rect -98639 -136558 -98583 -136514
rect -98539 -136558 -98483 -136514
rect -98439 -136558 -98383 -136514
rect -98339 -136558 -98283 -136514
rect -98239 -136558 -98183 -136514
rect -98139 -136558 -98083 -136514
rect -98039 -136558 -97983 -136514
rect -97939 -136558 -97883 -136514
rect -97839 -136558 -97783 -136514
rect -97739 -136558 -97683 -136514
rect -97639 -136558 -97583 -136514
rect -97539 -136558 -97483 -136514
rect -97439 -136558 -97383 -136514
rect -97339 -136558 -97283 -136514
rect -97239 -136558 -95895 -136514
rect -105360 -136614 -95895 -136558
rect -105360 -136658 -104783 -136614
rect -104739 -136658 -104683 -136614
rect -104639 -136658 -104583 -136614
rect -104539 -136658 -104483 -136614
rect -104439 -136658 -104383 -136614
rect -104339 -136658 -104283 -136614
rect -104239 -136658 -104183 -136614
rect -104139 -136658 -104083 -136614
rect -104039 -136658 -103983 -136614
rect -103939 -136658 -103883 -136614
rect -103839 -136658 -103783 -136614
rect -103739 -136658 -103683 -136614
rect -103639 -136658 -103583 -136614
rect -103539 -136658 -103483 -136614
rect -103439 -136658 -103383 -136614
rect -103339 -136658 -103283 -136614
rect -103239 -136658 -102783 -136614
rect -102739 -136658 -102683 -136614
rect -102639 -136658 -102583 -136614
rect -102539 -136658 -102483 -136614
rect -102439 -136658 -102383 -136614
rect -102339 -136658 -102283 -136614
rect -102239 -136658 -102183 -136614
rect -102139 -136658 -102083 -136614
rect -102039 -136658 -101983 -136614
rect -101939 -136658 -101883 -136614
rect -101839 -136658 -101783 -136614
rect -101739 -136658 -101683 -136614
rect -101639 -136658 -101583 -136614
rect -101539 -136658 -101483 -136614
rect -101439 -136658 -101383 -136614
rect -101339 -136658 -101283 -136614
rect -101239 -136658 -100783 -136614
rect -100739 -136658 -100683 -136614
rect -100639 -136658 -100583 -136614
rect -100539 -136658 -100483 -136614
rect -100439 -136658 -100383 -136614
rect -100339 -136658 -100283 -136614
rect -100239 -136658 -100183 -136614
rect -100139 -136658 -100083 -136614
rect -100039 -136658 -99983 -136614
rect -99939 -136658 -99883 -136614
rect -99839 -136658 -99783 -136614
rect -99739 -136658 -99683 -136614
rect -99639 -136658 -99583 -136614
rect -99539 -136658 -99483 -136614
rect -99439 -136658 -99383 -136614
rect -99339 -136658 -99283 -136614
rect -99239 -136658 -98783 -136614
rect -98739 -136658 -98683 -136614
rect -98639 -136658 -98583 -136614
rect -98539 -136658 -98483 -136614
rect -98439 -136658 -98383 -136614
rect -98339 -136658 -98283 -136614
rect -98239 -136658 -98183 -136614
rect -98139 -136658 -98083 -136614
rect -98039 -136658 -97983 -136614
rect -97939 -136658 -97883 -136614
rect -97839 -136658 -97783 -136614
rect -97739 -136658 -97683 -136614
rect -97639 -136658 -97583 -136614
rect -97539 -136658 -97483 -136614
rect -97439 -136658 -97383 -136614
rect -97339 -136658 -97283 -136614
rect -97239 -136658 -95895 -136614
rect -105360 -136714 -95895 -136658
rect -105360 -136758 -104783 -136714
rect -104739 -136758 -104683 -136714
rect -104639 -136758 -104583 -136714
rect -104539 -136758 -104483 -136714
rect -104439 -136758 -104383 -136714
rect -104339 -136758 -104283 -136714
rect -104239 -136758 -104183 -136714
rect -104139 -136758 -104083 -136714
rect -104039 -136758 -103983 -136714
rect -103939 -136758 -103883 -136714
rect -103839 -136758 -103783 -136714
rect -103739 -136758 -103683 -136714
rect -103639 -136758 -103583 -136714
rect -103539 -136758 -103483 -136714
rect -103439 -136758 -103383 -136714
rect -103339 -136758 -103283 -136714
rect -103239 -136758 -102783 -136714
rect -102739 -136758 -102683 -136714
rect -102639 -136758 -102583 -136714
rect -102539 -136758 -102483 -136714
rect -102439 -136758 -102383 -136714
rect -102339 -136758 -102283 -136714
rect -102239 -136758 -102183 -136714
rect -102139 -136758 -102083 -136714
rect -102039 -136758 -101983 -136714
rect -101939 -136758 -101883 -136714
rect -101839 -136758 -101783 -136714
rect -101739 -136758 -101683 -136714
rect -101639 -136758 -101583 -136714
rect -101539 -136758 -101483 -136714
rect -101439 -136758 -101383 -136714
rect -101339 -136758 -101283 -136714
rect -101239 -136758 -100783 -136714
rect -100739 -136758 -100683 -136714
rect -100639 -136758 -100583 -136714
rect -100539 -136758 -100483 -136714
rect -100439 -136758 -100383 -136714
rect -100339 -136758 -100283 -136714
rect -100239 -136758 -100183 -136714
rect -100139 -136758 -100083 -136714
rect -100039 -136758 -99983 -136714
rect -99939 -136758 -99883 -136714
rect -99839 -136758 -99783 -136714
rect -99739 -136758 -99683 -136714
rect -99639 -136758 -99583 -136714
rect -99539 -136758 -99483 -136714
rect -99439 -136758 -99383 -136714
rect -99339 -136758 -99283 -136714
rect -99239 -136758 -98783 -136714
rect -98739 -136758 -98683 -136714
rect -98639 -136758 -98583 -136714
rect -98539 -136758 -98483 -136714
rect -98439 -136758 -98383 -136714
rect -98339 -136758 -98283 -136714
rect -98239 -136758 -98183 -136714
rect -98139 -136758 -98083 -136714
rect -98039 -136758 -97983 -136714
rect -97939 -136758 -97883 -136714
rect -97839 -136758 -97783 -136714
rect -97739 -136758 -97683 -136714
rect -97639 -136758 -97583 -136714
rect -97539 -136758 -97483 -136714
rect -97439 -136758 -97383 -136714
rect -97339 -136758 -97283 -136714
rect -97239 -136758 -95895 -136714
rect -105360 -136814 -95895 -136758
rect -105360 -136858 -104783 -136814
rect -104739 -136858 -104683 -136814
rect -104639 -136858 -104583 -136814
rect -104539 -136858 -104483 -136814
rect -104439 -136858 -104383 -136814
rect -104339 -136858 -104283 -136814
rect -104239 -136858 -104183 -136814
rect -104139 -136858 -104083 -136814
rect -104039 -136858 -103983 -136814
rect -103939 -136858 -103883 -136814
rect -103839 -136858 -103783 -136814
rect -103739 -136858 -103683 -136814
rect -103639 -136858 -103583 -136814
rect -103539 -136858 -103483 -136814
rect -103439 -136858 -103383 -136814
rect -103339 -136858 -103283 -136814
rect -103239 -136858 -102783 -136814
rect -102739 -136858 -102683 -136814
rect -102639 -136858 -102583 -136814
rect -102539 -136858 -102483 -136814
rect -102439 -136858 -102383 -136814
rect -102339 -136858 -102283 -136814
rect -102239 -136858 -102183 -136814
rect -102139 -136858 -102083 -136814
rect -102039 -136858 -101983 -136814
rect -101939 -136858 -101883 -136814
rect -101839 -136858 -101783 -136814
rect -101739 -136858 -101683 -136814
rect -101639 -136858 -101583 -136814
rect -101539 -136858 -101483 -136814
rect -101439 -136858 -101383 -136814
rect -101339 -136858 -101283 -136814
rect -101239 -136858 -100783 -136814
rect -100739 -136858 -100683 -136814
rect -100639 -136858 -100583 -136814
rect -100539 -136858 -100483 -136814
rect -100439 -136858 -100383 -136814
rect -100339 -136858 -100283 -136814
rect -100239 -136858 -100183 -136814
rect -100139 -136858 -100083 -136814
rect -100039 -136858 -99983 -136814
rect -99939 -136858 -99883 -136814
rect -99839 -136858 -99783 -136814
rect -99739 -136858 -99683 -136814
rect -99639 -136858 -99583 -136814
rect -99539 -136858 -99483 -136814
rect -99439 -136858 -99383 -136814
rect -99339 -136858 -99283 -136814
rect -99239 -136858 -98783 -136814
rect -98739 -136858 -98683 -136814
rect -98639 -136858 -98583 -136814
rect -98539 -136858 -98483 -136814
rect -98439 -136858 -98383 -136814
rect -98339 -136858 -98283 -136814
rect -98239 -136858 -98183 -136814
rect -98139 -136858 -98083 -136814
rect -98039 -136858 -97983 -136814
rect -97939 -136858 -97883 -136814
rect -97839 -136858 -97783 -136814
rect -97739 -136858 -97683 -136814
rect -97639 -136858 -97583 -136814
rect -97539 -136858 -97483 -136814
rect -97439 -136858 -97383 -136814
rect -97339 -136858 -97283 -136814
rect -97239 -136858 -95895 -136814
rect -107141 -171279 -105588 -138781
rect -105360 -142610 -95895 -136858
rect -60256 -137966 174378 -136015
rect -60256 -138010 81632 -137966
rect 81676 -138010 81732 -137966
rect 81776 -138010 81832 -137966
rect 81876 -138010 81932 -137966
rect 81976 -138010 82032 -137966
rect 82076 -138010 82132 -137966
rect 82176 -138010 82232 -137966
rect 82276 -138010 82332 -137966
rect 82376 -138010 82432 -137966
rect 82476 -138010 82532 -137966
rect 82576 -138010 82632 -137966
rect 82676 -138010 82732 -137966
rect 82776 -138010 82832 -137966
rect 82876 -138010 82932 -137966
rect 82976 -138010 83032 -137966
rect 83076 -138010 83132 -137966
rect 83176 -138010 83632 -137966
rect 83676 -138010 83732 -137966
rect 83776 -138010 83832 -137966
rect 83876 -138010 83932 -137966
rect 83976 -138010 84032 -137966
rect 84076 -138010 84132 -137966
rect 84176 -138010 84232 -137966
rect 84276 -138010 84332 -137966
rect 84376 -138010 84432 -137966
rect 84476 -138010 84532 -137966
rect 84576 -138010 84632 -137966
rect 84676 -138010 84732 -137966
rect 84776 -138010 84832 -137966
rect 84876 -138010 84932 -137966
rect 84976 -138010 85032 -137966
rect 85076 -138010 85132 -137966
rect 85176 -138010 85632 -137966
rect 85676 -138010 85732 -137966
rect 85776 -138010 85832 -137966
rect 85876 -138010 85932 -137966
rect 85976 -138010 86032 -137966
rect 86076 -138010 86132 -137966
rect 86176 -138010 86232 -137966
rect 86276 -138010 86332 -137966
rect 86376 -138010 86432 -137966
rect 86476 -138010 86532 -137966
rect 86576 -138010 86632 -137966
rect 86676 -138010 86732 -137966
rect 86776 -138010 86832 -137966
rect 86876 -138010 86932 -137966
rect 86976 -138010 87032 -137966
rect 87076 -138010 87132 -137966
rect 87176 -138010 87632 -137966
rect 87676 -138010 87732 -137966
rect 87776 -138010 87832 -137966
rect 87876 -138010 87932 -137966
rect 87976 -138010 88032 -137966
rect 88076 -138010 88132 -137966
rect 88176 -138010 88232 -137966
rect 88276 -138010 88332 -137966
rect 88376 -138010 88432 -137966
rect 88476 -138010 88532 -137966
rect 88576 -138010 88632 -137966
rect 88676 -138010 88732 -137966
rect 88776 -138010 88832 -137966
rect 88876 -138010 88932 -137966
rect 88976 -138010 89032 -137966
rect 89076 -138010 89132 -137966
rect 89176 -138010 174378 -137966
rect -60256 -138066 174378 -138010
rect -60256 -138110 81632 -138066
rect 81676 -138110 81732 -138066
rect 81776 -138110 81832 -138066
rect 81876 -138110 81932 -138066
rect 81976 -138110 82032 -138066
rect 82076 -138110 82132 -138066
rect 82176 -138110 82232 -138066
rect 82276 -138110 82332 -138066
rect 82376 -138110 82432 -138066
rect 82476 -138110 82532 -138066
rect 82576 -138110 82632 -138066
rect 82676 -138110 82732 -138066
rect 82776 -138110 82832 -138066
rect 82876 -138110 82932 -138066
rect 82976 -138110 83032 -138066
rect 83076 -138110 83132 -138066
rect 83176 -138110 83632 -138066
rect 83676 -138110 83732 -138066
rect 83776 -138110 83832 -138066
rect 83876 -138110 83932 -138066
rect 83976 -138110 84032 -138066
rect 84076 -138110 84132 -138066
rect 84176 -138110 84232 -138066
rect 84276 -138110 84332 -138066
rect 84376 -138110 84432 -138066
rect 84476 -138110 84532 -138066
rect 84576 -138110 84632 -138066
rect 84676 -138110 84732 -138066
rect 84776 -138110 84832 -138066
rect 84876 -138110 84932 -138066
rect 84976 -138110 85032 -138066
rect 85076 -138110 85132 -138066
rect 85176 -138110 85632 -138066
rect 85676 -138110 85732 -138066
rect 85776 -138110 85832 -138066
rect 85876 -138110 85932 -138066
rect 85976 -138110 86032 -138066
rect 86076 -138110 86132 -138066
rect 86176 -138110 86232 -138066
rect 86276 -138110 86332 -138066
rect 86376 -138110 86432 -138066
rect 86476 -138110 86532 -138066
rect 86576 -138110 86632 -138066
rect 86676 -138110 86732 -138066
rect 86776 -138110 86832 -138066
rect 86876 -138110 86932 -138066
rect 86976 -138110 87032 -138066
rect 87076 -138110 87132 -138066
rect 87176 -138110 87632 -138066
rect 87676 -138110 87732 -138066
rect 87776 -138110 87832 -138066
rect 87876 -138110 87932 -138066
rect 87976 -138110 88032 -138066
rect 88076 -138110 88132 -138066
rect 88176 -138110 88232 -138066
rect 88276 -138110 88332 -138066
rect 88376 -138110 88432 -138066
rect 88476 -138110 88532 -138066
rect 88576 -138110 88632 -138066
rect 88676 -138110 88732 -138066
rect 88776 -138110 88832 -138066
rect 88876 -138110 88932 -138066
rect 88976 -138110 89032 -138066
rect 89076 -138110 89132 -138066
rect 89176 -138110 174378 -138066
rect -60256 -138166 174378 -138110
rect -60256 -138210 81632 -138166
rect 81676 -138210 81732 -138166
rect 81776 -138210 81832 -138166
rect 81876 -138210 81932 -138166
rect 81976 -138210 82032 -138166
rect 82076 -138210 82132 -138166
rect 82176 -138210 82232 -138166
rect 82276 -138210 82332 -138166
rect 82376 -138210 82432 -138166
rect 82476 -138210 82532 -138166
rect 82576 -138210 82632 -138166
rect 82676 -138210 82732 -138166
rect 82776 -138210 82832 -138166
rect 82876 -138210 82932 -138166
rect 82976 -138210 83032 -138166
rect 83076 -138210 83132 -138166
rect 83176 -138210 83632 -138166
rect 83676 -138210 83732 -138166
rect 83776 -138210 83832 -138166
rect 83876 -138210 83932 -138166
rect 83976 -138210 84032 -138166
rect 84076 -138210 84132 -138166
rect 84176 -138210 84232 -138166
rect 84276 -138210 84332 -138166
rect 84376 -138210 84432 -138166
rect 84476 -138210 84532 -138166
rect 84576 -138210 84632 -138166
rect 84676 -138210 84732 -138166
rect 84776 -138210 84832 -138166
rect 84876 -138210 84932 -138166
rect 84976 -138210 85032 -138166
rect 85076 -138210 85132 -138166
rect 85176 -138210 85632 -138166
rect 85676 -138210 85732 -138166
rect 85776 -138210 85832 -138166
rect 85876 -138210 85932 -138166
rect 85976 -138210 86032 -138166
rect 86076 -138210 86132 -138166
rect 86176 -138210 86232 -138166
rect 86276 -138210 86332 -138166
rect 86376 -138210 86432 -138166
rect 86476 -138210 86532 -138166
rect 86576 -138210 86632 -138166
rect 86676 -138210 86732 -138166
rect 86776 -138210 86832 -138166
rect 86876 -138210 86932 -138166
rect 86976 -138210 87032 -138166
rect 87076 -138210 87132 -138166
rect 87176 -138210 87632 -138166
rect 87676 -138210 87732 -138166
rect 87776 -138210 87832 -138166
rect 87876 -138210 87932 -138166
rect 87976 -138210 88032 -138166
rect 88076 -138210 88132 -138166
rect 88176 -138210 88232 -138166
rect 88276 -138210 88332 -138166
rect 88376 -138210 88432 -138166
rect 88476 -138210 88532 -138166
rect 88576 -138210 88632 -138166
rect 88676 -138210 88732 -138166
rect 88776 -138210 88832 -138166
rect 88876 -138210 88932 -138166
rect 88976 -138210 89032 -138166
rect 89076 -138210 89132 -138166
rect 89176 -138210 174378 -138166
rect -60256 -138266 174378 -138210
rect -105360 -143556 -103394 -142610
rect -102448 -143556 -95895 -142610
rect -105360 -144550 -95895 -143556
rect -85973 -140231 -72506 -138270
rect -85973 -140275 -83265 -140231
rect -83221 -140275 -83165 -140231
rect -83121 -140275 -83065 -140231
rect -83021 -140275 -82965 -140231
rect -82921 -140275 -82865 -140231
rect -82821 -140275 -82765 -140231
rect -82721 -140275 -82665 -140231
rect -82621 -140275 -82565 -140231
rect -82521 -140275 -82465 -140231
rect -82421 -140275 -82365 -140231
rect -82321 -140275 -82265 -140231
rect -82221 -140275 -82165 -140231
rect -82121 -140275 -82065 -140231
rect -82021 -140275 -81965 -140231
rect -81921 -140275 -81865 -140231
rect -81821 -140275 -81765 -140231
rect -81721 -140275 -81265 -140231
rect -81221 -140275 -81165 -140231
rect -81121 -140275 -81065 -140231
rect -81021 -140275 -80965 -140231
rect -80921 -140275 -80865 -140231
rect -80821 -140275 -80765 -140231
rect -80721 -140275 -80665 -140231
rect -80621 -140275 -80565 -140231
rect -80521 -140275 -80465 -140231
rect -80421 -140275 -80365 -140231
rect -80321 -140275 -80265 -140231
rect -80221 -140275 -80165 -140231
rect -80121 -140275 -80065 -140231
rect -80021 -140275 -79965 -140231
rect -79921 -140275 -79865 -140231
rect -79821 -140275 -79765 -140231
rect -79721 -140275 -79265 -140231
rect -79221 -140275 -79165 -140231
rect -79121 -140275 -79065 -140231
rect -79021 -140275 -78965 -140231
rect -78921 -140275 -78865 -140231
rect -78821 -140275 -78765 -140231
rect -78721 -140275 -78665 -140231
rect -78621 -140275 -78565 -140231
rect -78521 -140275 -78465 -140231
rect -78421 -140275 -78365 -140231
rect -78321 -140275 -78265 -140231
rect -78221 -140275 -78165 -140231
rect -78121 -140275 -78065 -140231
rect -78021 -140275 -77965 -140231
rect -77921 -140275 -77865 -140231
rect -77821 -140275 -77765 -140231
rect -77721 -140275 -77265 -140231
rect -77221 -140275 -77165 -140231
rect -77121 -140275 -77065 -140231
rect -77021 -140275 -76965 -140231
rect -76921 -140275 -76865 -140231
rect -76821 -140275 -76765 -140231
rect -76721 -140275 -76665 -140231
rect -76621 -140275 -76565 -140231
rect -76521 -140275 -76465 -140231
rect -76421 -140275 -76365 -140231
rect -76321 -140275 -76265 -140231
rect -76221 -140275 -76165 -140231
rect -76121 -140275 -76065 -140231
rect -76021 -140275 -75965 -140231
rect -75921 -140275 -75865 -140231
rect -75821 -140275 -75765 -140231
rect -75721 -140275 -72506 -140231
rect -85973 -140331 -72506 -140275
rect -85973 -140375 -83265 -140331
rect -83221 -140375 -83165 -140331
rect -83121 -140375 -83065 -140331
rect -83021 -140375 -82965 -140331
rect -82921 -140375 -82865 -140331
rect -82821 -140375 -82765 -140331
rect -82721 -140375 -82665 -140331
rect -82621 -140375 -82565 -140331
rect -82521 -140375 -82465 -140331
rect -82421 -140375 -82365 -140331
rect -82321 -140375 -82265 -140331
rect -82221 -140375 -82165 -140331
rect -82121 -140375 -82065 -140331
rect -82021 -140375 -81965 -140331
rect -81921 -140375 -81865 -140331
rect -81821 -140375 -81765 -140331
rect -81721 -140375 -81265 -140331
rect -81221 -140375 -81165 -140331
rect -81121 -140375 -81065 -140331
rect -81021 -140375 -80965 -140331
rect -80921 -140375 -80865 -140331
rect -80821 -140375 -80765 -140331
rect -80721 -140375 -80665 -140331
rect -80621 -140375 -80565 -140331
rect -80521 -140375 -80465 -140331
rect -80421 -140375 -80365 -140331
rect -80321 -140375 -80265 -140331
rect -80221 -140375 -80165 -140331
rect -80121 -140375 -80065 -140331
rect -80021 -140375 -79965 -140331
rect -79921 -140375 -79865 -140331
rect -79821 -140375 -79765 -140331
rect -79721 -140375 -79265 -140331
rect -79221 -140375 -79165 -140331
rect -79121 -140375 -79065 -140331
rect -79021 -140375 -78965 -140331
rect -78921 -140375 -78865 -140331
rect -78821 -140375 -78765 -140331
rect -78721 -140375 -78665 -140331
rect -78621 -140375 -78565 -140331
rect -78521 -140375 -78465 -140331
rect -78421 -140375 -78365 -140331
rect -78321 -140375 -78265 -140331
rect -78221 -140375 -78165 -140331
rect -78121 -140375 -78065 -140331
rect -78021 -140375 -77965 -140331
rect -77921 -140375 -77865 -140331
rect -77821 -140375 -77765 -140331
rect -77721 -140375 -77265 -140331
rect -77221 -140375 -77165 -140331
rect -77121 -140375 -77065 -140331
rect -77021 -140375 -76965 -140331
rect -76921 -140375 -76865 -140331
rect -76821 -140375 -76765 -140331
rect -76721 -140375 -76665 -140331
rect -76621 -140375 -76565 -140331
rect -76521 -140375 -76465 -140331
rect -76421 -140375 -76365 -140331
rect -76321 -140375 -76265 -140331
rect -76221 -140375 -76165 -140331
rect -76121 -140375 -76065 -140331
rect -76021 -140375 -75965 -140331
rect -75921 -140375 -75865 -140331
rect -75821 -140375 -75765 -140331
rect -75721 -140375 -72506 -140331
rect -85973 -140431 -72506 -140375
rect -85973 -140475 -83265 -140431
rect -83221 -140475 -83165 -140431
rect -83121 -140475 -83065 -140431
rect -83021 -140475 -82965 -140431
rect -82921 -140475 -82865 -140431
rect -82821 -140475 -82765 -140431
rect -82721 -140475 -82665 -140431
rect -82621 -140475 -82565 -140431
rect -82521 -140475 -82465 -140431
rect -82421 -140475 -82365 -140431
rect -82321 -140475 -82265 -140431
rect -82221 -140475 -82165 -140431
rect -82121 -140475 -82065 -140431
rect -82021 -140475 -81965 -140431
rect -81921 -140475 -81865 -140431
rect -81821 -140475 -81765 -140431
rect -81721 -140475 -81265 -140431
rect -81221 -140475 -81165 -140431
rect -81121 -140475 -81065 -140431
rect -81021 -140475 -80965 -140431
rect -80921 -140475 -80865 -140431
rect -80821 -140475 -80765 -140431
rect -80721 -140475 -80665 -140431
rect -80621 -140475 -80565 -140431
rect -80521 -140475 -80465 -140431
rect -80421 -140475 -80365 -140431
rect -80321 -140475 -80265 -140431
rect -80221 -140475 -80165 -140431
rect -80121 -140475 -80065 -140431
rect -80021 -140475 -79965 -140431
rect -79921 -140475 -79865 -140431
rect -79821 -140475 -79765 -140431
rect -79721 -140475 -79265 -140431
rect -79221 -140475 -79165 -140431
rect -79121 -140475 -79065 -140431
rect -79021 -140475 -78965 -140431
rect -78921 -140475 -78865 -140431
rect -78821 -140475 -78765 -140431
rect -78721 -140475 -78665 -140431
rect -78621 -140475 -78565 -140431
rect -78521 -140475 -78465 -140431
rect -78421 -140475 -78365 -140431
rect -78321 -140475 -78265 -140431
rect -78221 -140475 -78165 -140431
rect -78121 -140475 -78065 -140431
rect -78021 -140475 -77965 -140431
rect -77921 -140475 -77865 -140431
rect -77821 -140475 -77765 -140431
rect -77721 -140475 -77265 -140431
rect -77221 -140475 -77165 -140431
rect -77121 -140475 -77065 -140431
rect -77021 -140475 -76965 -140431
rect -76921 -140475 -76865 -140431
rect -76821 -140475 -76765 -140431
rect -76721 -140475 -76665 -140431
rect -76621 -140475 -76565 -140431
rect -76521 -140475 -76465 -140431
rect -76421 -140475 -76365 -140431
rect -76321 -140475 -76265 -140431
rect -76221 -140475 -76165 -140431
rect -76121 -140475 -76065 -140431
rect -76021 -140475 -75965 -140431
rect -75921 -140475 -75865 -140431
rect -75821 -140475 -75765 -140431
rect -75721 -140475 -72506 -140431
rect -85973 -140531 -72506 -140475
rect -85973 -140575 -83265 -140531
rect -83221 -140575 -83165 -140531
rect -83121 -140575 -83065 -140531
rect -83021 -140575 -82965 -140531
rect -82921 -140575 -82865 -140531
rect -82821 -140575 -82765 -140531
rect -82721 -140575 -82665 -140531
rect -82621 -140575 -82565 -140531
rect -82521 -140575 -82465 -140531
rect -82421 -140575 -82365 -140531
rect -82321 -140575 -82265 -140531
rect -82221 -140575 -82165 -140531
rect -82121 -140575 -82065 -140531
rect -82021 -140575 -81965 -140531
rect -81921 -140575 -81865 -140531
rect -81821 -140575 -81765 -140531
rect -81721 -140575 -81265 -140531
rect -81221 -140575 -81165 -140531
rect -81121 -140575 -81065 -140531
rect -81021 -140575 -80965 -140531
rect -80921 -140575 -80865 -140531
rect -80821 -140575 -80765 -140531
rect -80721 -140575 -80665 -140531
rect -80621 -140575 -80565 -140531
rect -80521 -140575 -80465 -140531
rect -80421 -140575 -80365 -140531
rect -80321 -140575 -80265 -140531
rect -80221 -140575 -80165 -140531
rect -80121 -140575 -80065 -140531
rect -80021 -140575 -79965 -140531
rect -79921 -140575 -79865 -140531
rect -79821 -140575 -79765 -140531
rect -79721 -140575 -79265 -140531
rect -79221 -140575 -79165 -140531
rect -79121 -140575 -79065 -140531
rect -79021 -140575 -78965 -140531
rect -78921 -140575 -78865 -140531
rect -78821 -140575 -78765 -140531
rect -78721 -140575 -78665 -140531
rect -78621 -140575 -78565 -140531
rect -78521 -140575 -78465 -140531
rect -78421 -140575 -78365 -140531
rect -78321 -140575 -78265 -140531
rect -78221 -140575 -78165 -140531
rect -78121 -140575 -78065 -140531
rect -78021 -140575 -77965 -140531
rect -77921 -140575 -77865 -140531
rect -77821 -140575 -77765 -140531
rect -77721 -140575 -77265 -140531
rect -77221 -140575 -77165 -140531
rect -77121 -140575 -77065 -140531
rect -77021 -140575 -76965 -140531
rect -76921 -140575 -76865 -140531
rect -76821 -140575 -76765 -140531
rect -76721 -140575 -76665 -140531
rect -76621 -140575 -76565 -140531
rect -76521 -140575 -76465 -140531
rect -76421 -140575 -76365 -140531
rect -76321 -140575 -76265 -140531
rect -76221 -140575 -76165 -140531
rect -76121 -140575 -76065 -140531
rect -76021 -140575 -75965 -140531
rect -75921 -140575 -75865 -140531
rect -75821 -140575 -75765 -140531
rect -75721 -140575 -72506 -140531
rect -85973 -140631 -72506 -140575
rect -85973 -140675 -83265 -140631
rect -83221 -140675 -83165 -140631
rect -83121 -140675 -83065 -140631
rect -83021 -140675 -82965 -140631
rect -82921 -140675 -82865 -140631
rect -82821 -140675 -82765 -140631
rect -82721 -140675 -82665 -140631
rect -82621 -140675 -82565 -140631
rect -82521 -140675 -82465 -140631
rect -82421 -140675 -82365 -140631
rect -82321 -140675 -82265 -140631
rect -82221 -140675 -82165 -140631
rect -82121 -140675 -82065 -140631
rect -82021 -140675 -81965 -140631
rect -81921 -140675 -81865 -140631
rect -81821 -140675 -81765 -140631
rect -81721 -140675 -81265 -140631
rect -81221 -140675 -81165 -140631
rect -81121 -140675 -81065 -140631
rect -81021 -140675 -80965 -140631
rect -80921 -140675 -80865 -140631
rect -80821 -140675 -80765 -140631
rect -80721 -140675 -80665 -140631
rect -80621 -140675 -80565 -140631
rect -80521 -140675 -80465 -140631
rect -80421 -140675 -80365 -140631
rect -80321 -140675 -80265 -140631
rect -80221 -140675 -80165 -140631
rect -80121 -140675 -80065 -140631
rect -80021 -140675 -79965 -140631
rect -79921 -140675 -79865 -140631
rect -79821 -140675 -79765 -140631
rect -79721 -140675 -79265 -140631
rect -79221 -140675 -79165 -140631
rect -79121 -140675 -79065 -140631
rect -79021 -140675 -78965 -140631
rect -78921 -140675 -78865 -140631
rect -78821 -140675 -78765 -140631
rect -78721 -140675 -78665 -140631
rect -78621 -140675 -78565 -140631
rect -78521 -140675 -78465 -140631
rect -78421 -140675 -78365 -140631
rect -78321 -140675 -78265 -140631
rect -78221 -140675 -78165 -140631
rect -78121 -140675 -78065 -140631
rect -78021 -140675 -77965 -140631
rect -77921 -140675 -77865 -140631
rect -77821 -140675 -77765 -140631
rect -77721 -140675 -77265 -140631
rect -77221 -140675 -77165 -140631
rect -77121 -140675 -77065 -140631
rect -77021 -140675 -76965 -140631
rect -76921 -140675 -76865 -140631
rect -76821 -140675 -76765 -140631
rect -76721 -140675 -76665 -140631
rect -76621 -140675 -76565 -140631
rect -76521 -140675 -76465 -140631
rect -76421 -140675 -76365 -140631
rect -76321 -140675 -76265 -140631
rect -76221 -140675 -76165 -140631
rect -76121 -140675 -76065 -140631
rect -76021 -140675 -75965 -140631
rect -75921 -140675 -75865 -140631
rect -75821 -140675 -75765 -140631
rect -75721 -140675 -72506 -140631
rect -85973 -140731 -72506 -140675
rect -85973 -140775 -83265 -140731
rect -83221 -140775 -83165 -140731
rect -83121 -140775 -83065 -140731
rect -83021 -140775 -82965 -140731
rect -82921 -140775 -82865 -140731
rect -82821 -140775 -82765 -140731
rect -82721 -140775 -82665 -140731
rect -82621 -140775 -82565 -140731
rect -82521 -140775 -82465 -140731
rect -82421 -140775 -82365 -140731
rect -82321 -140775 -82265 -140731
rect -82221 -140775 -82165 -140731
rect -82121 -140775 -82065 -140731
rect -82021 -140775 -81965 -140731
rect -81921 -140775 -81865 -140731
rect -81821 -140775 -81765 -140731
rect -81721 -140775 -81265 -140731
rect -81221 -140775 -81165 -140731
rect -81121 -140775 -81065 -140731
rect -81021 -140775 -80965 -140731
rect -80921 -140775 -80865 -140731
rect -80821 -140775 -80765 -140731
rect -80721 -140775 -80665 -140731
rect -80621 -140775 -80565 -140731
rect -80521 -140775 -80465 -140731
rect -80421 -140775 -80365 -140731
rect -80321 -140775 -80265 -140731
rect -80221 -140775 -80165 -140731
rect -80121 -140775 -80065 -140731
rect -80021 -140775 -79965 -140731
rect -79921 -140775 -79865 -140731
rect -79821 -140775 -79765 -140731
rect -79721 -140775 -79265 -140731
rect -79221 -140775 -79165 -140731
rect -79121 -140775 -79065 -140731
rect -79021 -140775 -78965 -140731
rect -78921 -140775 -78865 -140731
rect -78821 -140775 -78765 -140731
rect -78721 -140775 -78665 -140731
rect -78621 -140775 -78565 -140731
rect -78521 -140775 -78465 -140731
rect -78421 -140775 -78365 -140731
rect -78321 -140775 -78265 -140731
rect -78221 -140775 -78165 -140731
rect -78121 -140775 -78065 -140731
rect -78021 -140775 -77965 -140731
rect -77921 -140775 -77865 -140731
rect -77821 -140775 -77765 -140731
rect -77721 -140775 -77265 -140731
rect -77221 -140775 -77165 -140731
rect -77121 -140775 -77065 -140731
rect -77021 -140775 -76965 -140731
rect -76921 -140775 -76865 -140731
rect -76821 -140775 -76765 -140731
rect -76721 -140775 -76665 -140731
rect -76621 -140775 -76565 -140731
rect -76521 -140775 -76465 -140731
rect -76421 -140775 -76365 -140731
rect -76321 -140775 -76265 -140731
rect -76221 -140775 -76165 -140731
rect -76121 -140775 -76065 -140731
rect -76021 -140775 -75965 -140731
rect -75921 -140775 -75865 -140731
rect -75821 -140775 -75765 -140731
rect -75721 -140775 -72506 -140731
rect -85973 -140831 -72506 -140775
rect -85973 -140875 -83265 -140831
rect -83221 -140875 -83165 -140831
rect -83121 -140875 -83065 -140831
rect -83021 -140875 -82965 -140831
rect -82921 -140875 -82865 -140831
rect -82821 -140875 -82765 -140831
rect -82721 -140875 -82665 -140831
rect -82621 -140875 -82565 -140831
rect -82521 -140875 -82465 -140831
rect -82421 -140875 -82365 -140831
rect -82321 -140875 -82265 -140831
rect -82221 -140875 -82165 -140831
rect -82121 -140875 -82065 -140831
rect -82021 -140875 -81965 -140831
rect -81921 -140875 -81865 -140831
rect -81821 -140875 -81765 -140831
rect -81721 -140875 -81265 -140831
rect -81221 -140875 -81165 -140831
rect -81121 -140875 -81065 -140831
rect -81021 -140875 -80965 -140831
rect -80921 -140875 -80865 -140831
rect -80821 -140875 -80765 -140831
rect -80721 -140875 -80665 -140831
rect -80621 -140875 -80565 -140831
rect -80521 -140875 -80465 -140831
rect -80421 -140875 -80365 -140831
rect -80321 -140875 -80265 -140831
rect -80221 -140875 -80165 -140831
rect -80121 -140875 -80065 -140831
rect -80021 -140875 -79965 -140831
rect -79921 -140875 -79865 -140831
rect -79821 -140875 -79765 -140831
rect -79721 -140875 -79265 -140831
rect -79221 -140875 -79165 -140831
rect -79121 -140875 -79065 -140831
rect -79021 -140875 -78965 -140831
rect -78921 -140875 -78865 -140831
rect -78821 -140875 -78765 -140831
rect -78721 -140875 -78665 -140831
rect -78621 -140875 -78565 -140831
rect -78521 -140875 -78465 -140831
rect -78421 -140875 -78365 -140831
rect -78321 -140875 -78265 -140831
rect -78221 -140875 -78165 -140831
rect -78121 -140875 -78065 -140831
rect -78021 -140875 -77965 -140831
rect -77921 -140875 -77865 -140831
rect -77821 -140875 -77765 -140831
rect -77721 -140875 -77265 -140831
rect -77221 -140875 -77165 -140831
rect -77121 -140875 -77065 -140831
rect -77021 -140875 -76965 -140831
rect -76921 -140875 -76865 -140831
rect -76821 -140875 -76765 -140831
rect -76721 -140875 -76665 -140831
rect -76621 -140875 -76565 -140831
rect -76521 -140875 -76465 -140831
rect -76421 -140875 -76365 -140831
rect -76321 -140875 -76265 -140831
rect -76221 -140875 -76165 -140831
rect -76121 -140875 -76065 -140831
rect -76021 -140875 -75965 -140831
rect -75921 -140875 -75865 -140831
rect -75821 -140875 -75765 -140831
rect -75721 -140875 -72506 -140831
rect -85973 -140931 -72506 -140875
rect -85973 -140975 -83265 -140931
rect -83221 -140975 -83165 -140931
rect -83121 -140975 -83065 -140931
rect -83021 -140975 -82965 -140931
rect -82921 -140975 -82865 -140931
rect -82821 -140975 -82765 -140931
rect -82721 -140975 -82665 -140931
rect -82621 -140975 -82565 -140931
rect -82521 -140975 -82465 -140931
rect -82421 -140975 -82365 -140931
rect -82321 -140975 -82265 -140931
rect -82221 -140975 -82165 -140931
rect -82121 -140975 -82065 -140931
rect -82021 -140975 -81965 -140931
rect -81921 -140975 -81865 -140931
rect -81821 -140975 -81765 -140931
rect -81721 -140975 -81265 -140931
rect -81221 -140975 -81165 -140931
rect -81121 -140975 -81065 -140931
rect -81021 -140975 -80965 -140931
rect -80921 -140975 -80865 -140931
rect -80821 -140975 -80765 -140931
rect -80721 -140975 -80665 -140931
rect -80621 -140975 -80565 -140931
rect -80521 -140975 -80465 -140931
rect -80421 -140975 -80365 -140931
rect -80321 -140975 -80265 -140931
rect -80221 -140975 -80165 -140931
rect -80121 -140975 -80065 -140931
rect -80021 -140975 -79965 -140931
rect -79921 -140975 -79865 -140931
rect -79821 -140975 -79765 -140931
rect -79721 -140975 -79265 -140931
rect -79221 -140975 -79165 -140931
rect -79121 -140975 -79065 -140931
rect -79021 -140975 -78965 -140931
rect -78921 -140975 -78865 -140931
rect -78821 -140975 -78765 -140931
rect -78721 -140975 -78665 -140931
rect -78621 -140975 -78565 -140931
rect -78521 -140975 -78465 -140931
rect -78421 -140975 -78365 -140931
rect -78321 -140975 -78265 -140931
rect -78221 -140975 -78165 -140931
rect -78121 -140975 -78065 -140931
rect -78021 -140975 -77965 -140931
rect -77921 -140975 -77865 -140931
rect -77821 -140975 -77765 -140931
rect -77721 -140975 -77265 -140931
rect -77221 -140975 -77165 -140931
rect -77121 -140975 -77065 -140931
rect -77021 -140975 -76965 -140931
rect -76921 -140975 -76865 -140931
rect -76821 -140975 -76765 -140931
rect -76721 -140975 -76665 -140931
rect -76621 -140975 -76565 -140931
rect -76521 -140975 -76465 -140931
rect -76421 -140975 -76365 -140931
rect -76321 -140975 -76265 -140931
rect -76221 -140975 -76165 -140931
rect -76121 -140975 -76065 -140931
rect -76021 -140975 -75965 -140931
rect -75921 -140975 -75865 -140931
rect -75821 -140975 -75765 -140931
rect -75721 -140975 -72506 -140931
rect -85973 -141031 -72506 -140975
rect -85973 -141075 -83265 -141031
rect -83221 -141075 -83165 -141031
rect -83121 -141075 -83065 -141031
rect -83021 -141075 -82965 -141031
rect -82921 -141075 -82865 -141031
rect -82821 -141075 -82765 -141031
rect -82721 -141075 -82665 -141031
rect -82621 -141075 -82565 -141031
rect -82521 -141075 -82465 -141031
rect -82421 -141075 -82365 -141031
rect -82321 -141075 -82265 -141031
rect -82221 -141075 -82165 -141031
rect -82121 -141075 -82065 -141031
rect -82021 -141075 -81965 -141031
rect -81921 -141075 -81865 -141031
rect -81821 -141075 -81765 -141031
rect -81721 -141075 -81265 -141031
rect -81221 -141075 -81165 -141031
rect -81121 -141075 -81065 -141031
rect -81021 -141075 -80965 -141031
rect -80921 -141075 -80865 -141031
rect -80821 -141075 -80765 -141031
rect -80721 -141075 -80665 -141031
rect -80621 -141075 -80565 -141031
rect -80521 -141075 -80465 -141031
rect -80421 -141075 -80365 -141031
rect -80321 -141075 -80265 -141031
rect -80221 -141075 -80165 -141031
rect -80121 -141075 -80065 -141031
rect -80021 -141075 -79965 -141031
rect -79921 -141075 -79865 -141031
rect -79821 -141075 -79765 -141031
rect -79721 -141075 -79265 -141031
rect -79221 -141075 -79165 -141031
rect -79121 -141075 -79065 -141031
rect -79021 -141075 -78965 -141031
rect -78921 -141075 -78865 -141031
rect -78821 -141075 -78765 -141031
rect -78721 -141075 -78665 -141031
rect -78621 -141075 -78565 -141031
rect -78521 -141075 -78465 -141031
rect -78421 -141075 -78365 -141031
rect -78321 -141075 -78265 -141031
rect -78221 -141075 -78165 -141031
rect -78121 -141075 -78065 -141031
rect -78021 -141075 -77965 -141031
rect -77921 -141075 -77865 -141031
rect -77821 -141075 -77765 -141031
rect -77721 -141075 -77265 -141031
rect -77221 -141075 -77165 -141031
rect -77121 -141075 -77065 -141031
rect -77021 -141075 -76965 -141031
rect -76921 -141075 -76865 -141031
rect -76821 -141075 -76765 -141031
rect -76721 -141075 -76665 -141031
rect -76621 -141075 -76565 -141031
rect -76521 -141075 -76465 -141031
rect -76421 -141075 -76365 -141031
rect -76321 -141075 -76265 -141031
rect -76221 -141075 -76165 -141031
rect -76121 -141075 -76065 -141031
rect -76021 -141075 -75965 -141031
rect -75921 -141075 -75865 -141031
rect -75821 -141075 -75765 -141031
rect -75721 -141075 -72506 -141031
rect -85973 -141131 -72506 -141075
rect -85973 -141175 -83265 -141131
rect -83221 -141175 -83165 -141131
rect -83121 -141175 -83065 -141131
rect -83021 -141175 -82965 -141131
rect -82921 -141175 -82865 -141131
rect -82821 -141175 -82765 -141131
rect -82721 -141175 -82665 -141131
rect -82621 -141175 -82565 -141131
rect -82521 -141175 -82465 -141131
rect -82421 -141175 -82365 -141131
rect -82321 -141175 -82265 -141131
rect -82221 -141175 -82165 -141131
rect -82121 -141175 -82065 -141131
rect -82021 -141175 -81965 -141131
rect -81921 -141175 -81865 -141131
rect -81821 -141175 -81765 -141131
rect -81721 -141175 -81265 -141131
rect -81221 -141175 -81165 -141131
rect -81121 -141175 -81065 -141131
rect -81021 -141175 -80965 -141131
rect -80921 -141175 -80865 -141131
rect -80821 -141175 -80765 -141131
rect -80721 -141175 -80665 -141131
rect -80621 -141175 -80565 -141131
rect -80521 -141175 -80465 -141131
rect -80421 -141175 -80365 -141131
rect -80321 -141175 -80265 -141131
rect -80221 -141175 -80165 -141131
rect -80121 -141175 -80065 -141131
rect -80021 -141175 -79965 -141131
rect -79921 -141175 -79865 -141131
rect -79821 -141175 -79765 -141131
rect -79721 -141175 -79265 -141131
rect -79221 -141175 -79165 -141131
rect -79121 -141175 -79065 -141131
rect -79021 -141175 -78965 -141131
rect -78921 -141175 -78865 -141131
rect -78821 -141175 -78765 -141131
rect -78721 -141175 -78665 -141131
rect -78621 -141175 -78565 -141131
rect -78521 -141175 -78465 -141131
rect -78421 -141175 -78365 -141131
rect -78321 -141175 -78265 -141131
rect -78221 -141175 -78165 -141131
rect -78121 -141175 -78065 -141131
rect -78021 -141175 -77965 -141131
rect -77921 -141175 -77865 -141131
rect -77821 -141175 -77765 -141131
rect -77721 -141175 -77265 -141131
rect -77221 -141175 -77165 -141131
rect -77121 -141175 -77065 -141131
rect -77021 -141175 -76965 -141131
rect -76921 -141175 -76865 -141131
rect -76821 -141175 -76765 -141131
rect -76721 -141175 -76665 -141131
rect -76621 -141175 -76565 -141131
rect -76521 -141175 -76465 -141131
rect -76421 -141175 -76365 -141131
rect -76321 -141175 -76265 -141131
rect -76221 -141175 -76165 -141131
rect -76121 -141175 -76065 -141131
rect -76021 -141175 -75965 -141131
rect -75921 -141175 -75865 -141131
rect -75821 -141175 -75765 -141131
rect -75721 -141175 -72506 -141131
rect -85973 -141231 -72506 -141175
rect -85973 -141275 -83265 -141231
rect -83221 -141275 -83165 -141231
rect -83121 -141275 -83065 -141231
rect -83021 -141275 -82965 -141231
rect -82921 -141275 -82865 -141231
rect -82821 -141275 -82765 -141231
rect -82721 -141275 -82665 -141231
rect -82621 -141275 -82565 -141231
rect -82521 -141275 -82465 -141231
rect -82421 -141275 -82365 -141231
rect -82321 -141275 -82265 -141231
rect -82221 -141275 -82165 -141231
rect -82121 -141275 -82065 -141231
rect -82021 -141275 -81965 -141231
rect -81921 -141275 -81865 -141231
rect -81821 -141275 -81765 -141231
rect -81721 -141275 -81265 -141231
rect -81221 -141275 -81165 -141231
rect -81121 -141275 -81065 -141231
rect -81021 -141275 -80965 -141231
rect -80921 -141275 -80865 -141231
rect -80821 -141275 -80765 -141231
rect -80721 -141275 -80665 -141231
rect -80621 -141275 -80565 -141231
rect -80521 -141275 -80465 -141231
rect -80421 -141275 -80365 -141231
rect -80321 -141275 -80265 -141231
rect -80221 -141275 -80165 -141231
rect -80121 -141275 -80065 -141231
rect -80021 -141275 -79965 -141231
rect -79921 -141275 -79865 -141231
rect -79821 -141275 -79765 -141231
rect -79721 -141275 -79265 -141231
rect -79221 -141275 -79165 -141231
rect -79121 -141275 -79065 -141231
rect -79021 -141275 -78965 -141231
rect -78921 -141275 -78865 -141231
rect -78821 -141275 -78765 -141231
rect -78721 -141275 -78665 -141231
rect -78621 -141275 -78565 -141231
rect -78521 -141275 -78465 -141231
rect -78421 -141275 -78365 -141231
rect -78321 -141275 -78265 -141231
rect -78221 -141275 -78165 -141231
rect -78121 -141275 -78065 -141231
rect -78021 -141275 -77965 -141231
rect -77921 -141275 -77865 -141231
rect -77821 -141275 -77765 -141231
rect -77721 -141275 -77265 -141231
rect -77221 -141275 -77165 -141231
rect -77121 -141275 -77065 -141231
rect -77021 -141275 -76965 -141231
rect -76921 -141275 -76865 -141231
rect -76821 -141275 -76765 -141231
rect -76721 -141275 -76665 -141231
rect -76621 -141275 -76565 -141231
rect -76521 -141275 -76465 -141231
rect -76421 -141275 -76365 -141231
rect -76321 -141275 -76265 -141231
rect -76221 -141275 -76165 -141231
rect -76121 -141275 -76065 -141231
rect -76021 -141275 -75965 -141231
rect -75921 -141275 -75865 -141231
rect -75821 -141275 -75765 -141231
rect -75721 -141275 -72506 -141231
rect -85973 -141331 -72506 -141275
rect -85973 -141375 -83265 -141331
rect -83221 -141375 -83165 -141331
rect -83121 -141375 -83065 -141331
rect -83021 -141375 -82965 -141331
rect -82921 -141375 -82865 -141331
rect -82821 -141375 -82765 -141331
rect -82721 -141375 -82665 -141331
rect -82621 -141375 -82565 -141331
rect -82521 -141375 -82465 -141331
rect -82421 -141375 -82365 -141331
rect -82321 -141375 -82265 -141331
rect -82221 -141375 -82165 -141331
rect -82121 -141375 -82065 -141331
rect -82021 -141375 -81965 -141331
rect -81921 -141375 -81865 -141331
rect -81821 -141375 -81765 -141331
rect -81721 -141375 -81265 -141331
rect -81221 -141375 -81165 -141331
rect -81121 -141375 -81065 -141331
rect -81021 -141375 -80965 -141331
rect -80921 -141375 -80865 -141331
rect -80821 -141375 -80765 -141331
rect -80721 -141375 -80665 -141331
rect -80621 -141375 -80565 -141331
rect -80521 -141375 -80465 -141331
rect -80421 -141375 -80365 -141331
rect -80321 -141375 -80265 -141331
rect -80221 -141375 -80165 -141331
rect -80121 -141375 -80065 -141331
rect -80021 -141375 -79965 -141331
rect -79921 -141375 -79865 -141331
rect -79821 -141375 -79765 -141331
rect -79721 -141375 -79265 -141331
rect -79221 -141375 -79165 -141331
rect -79121 -141375 -79065 -141331
rect -79021 -141375 -78965 -141331
rect -78921 -141375 -78865 -141331
rect -78821 -141375 -78765 -141331
rect -78721 -141375 -78665 -141331
rect -78621 -141375 -78565 -141331
rect -78521 -141375 -78465 -141331
rect -78421 -141375 -78365 -141331
rect -78321 -141375 -78265 -141331
rect -78221 -141375 -78165 -141331
rect -78121 -141375 -78065 -141331
rect -78021 -141375 -77965 -141331
rect -77921 -141375 -77865 -141331
rect -77821 -141375 -77765 -141331
rect -77721 -141375 -77265 -141331
rect -77221 -141375 -77165 -141331
rect -77121 -141375 -77065 -141331
rect -77021 -141375 -76965 -141331
rect -76921 -141375 -76865 -141331
rect -76821 -141375 -76765 -141331
rect -76721 -141375 -76665 -141331
rect -76621 -141375 -76565 -141331
rect -76521 -141375 -76465 -141331
rect -76421 -141375 -76365 -141331
rect -76321 -141375 -76265 -141331
rect -76221 -141375 -76165 -141331
rect -76121 -141375 -76065 -141331
rect -76021 -141375 -75965 -141331
rect -75921 -141375 -75865 -141331
rect -75821 -141375 -75765 -141331
rect -75721 -141375 -72506 -141331
rect -85973 -141431 -72506 -141375
rect -85973 -141475 -83265 -141431
rect -83221 -141475 -83165 -141431
rect -83121 -141475 -83065 -141431
rect -83021 -141475 -82965 -141431
rect -82921 -141475 -82865 -141431
rect -82821 -141475 -82765 -141431
rect -82721 -141475 -82665 -141431
rect -82621 -141475 -82565 -141431
rect -82521 -141475 -82465 -141431
rect -82421 -141475 -82365 -141431
rect -82321 -141475 -82265 -141431
rect -82221 -141475 -82165 -141431
rect -82121 -141475 -82065 -141431
rect -82021 -141475 -81965 -141431
rect -81921 -141475 -81865 -141431
rect -81821 -141475 -81765 -141431
rect -81721 -141475 -81265 -141431
rect -81221 -141475 -81165 -141431
rect -81121 -141475 -81065 -141431
rect -81021 -141475 -80965 -141431
rect -80921 -141475 -80865 -141431
rect -80821 -141475 -80765 -141431
rect -80721 -141475 -80665 -141431
rect -80621 -141475 -80565 -141431
rect -80521 -141475 -80465 -141431
rect -80421 -141475 -80365 -141431
rect -80321 -141475 -80265 -141431
rect -80221 -141475 -80165 -141431
rect -80121 -141475 -80065 -141431
rect -80021 -141475 -79965 -141431
rect -79921 -141475 -79865 -141431
rect -79821 -141475 -79765 -141431
rect -79721 -141475 -79265 -141431
rect -79221 -141475 -79165 -141431
rect -79121 -141475 -79065 -141431
rect -79021 -141475 -78965 -141431
rect -78921 -141475 -78865 -141431
rect -78821 -141475 -78765 -141431
rect -78721 -141475 -78665 -141431
rect -78621 -141475 -78565 -141431
rect -78521 -141475 -78465 -141431
rect -78421 -141475 -78365 -141431
rect -78321 -141475 -78265 -141431
rect -78221 -141475 -78165 -141431
rect -78121 -141475 -78065 -141431
rect -78021 -141475 -77965 -141431
rect -77921 -141475 -77865 -141431
rect -77821 -141475 -77765 -141431
rect -77721 -141475 -77265 -141431
rect -77221 -141475 -77165 -141431
rect -77121 -141475 -77065 -141431
rect -77021 -141475 -76965 -141431
rect -76921 -141475 -76865 -141431
rect -76821 -141475 -76765 -141431
rect -76721 -141475 -76665 -141431
rect -76621 -141475 -76565 -141431
rect -76521 -141475 -76465 -141431
rect -76421 -141475 -76365 -141431
rect -76321 -141475 -76265 -141431
rect -76221 -141475 -76165 -141431
rect -76121 -141475 -76065 -141431
rect -76021 -141475 -75965 -141431
rect -75921 -141475 -75865 -141431
rect -75821 -141475 -75765 -141431
rect -75721 -141475 -72506 -141431
rect -85973 -141531 -72506 -141475
rect -85973 -141575 -83265 -141531
rect -83221 -141575 -83165 -141531
rect -83121 -141575 -83065 -141531
rect -83021 -141575 -82965 -141531
rect -82921 -141575 -82865 -141531
rect -82821 -141575 -82765 -141531
rect -82721 -141575 -82665 -141531
rect -82621 -141575 -82565 -141531
rect -82521 -141575 -82465 -141531
rect -82421 -141575 -82365 -141531
rect -82321 -141575 -82265 -141531
rect -82221 -141575 -82165 -141531
rect -82121 -141575 -82065 -141531
rect -82021 -141575 -81965 -141531
rect -81921 -141575 -81865 -141531
rect -81821 -141575 -81765 -141531
rect -81721 -141575 -81265 -141531
rect -81221 -141575 -81165 -141531
rect -81121 -141575 -81065 -141531
rect -81021 -141575 -80965 -141531
rect -80921 -141575 -80865 -141531
rect -80821 -141575 -80765 -141531
rect -80721 -141575 -80665 -141531
rect -80621 -141575 -80565 -141531
rect -80521 -141575 -80465 -141531
rect -80421 -141575 -80365 -141531
rect -80321 -141575 -80265 -141531
rect -80221 -141575 -80165 -141531
rect -80121 -141575 -80065 -141531
rect -80021 -141575 -79965 -141531
rect -79921 -141575 -79865 -141531
rect -79821 -141575 -79765 -141531
rect -79721 -141575 -79265 -141531
rect -79221 -141575 -79165 -141531
rect -79121 -141575 -79065 -141531
rect -79021 -141575 -78965 -141531
rect -78921 -141575 -78865 -141531
rect -78821 -141575 -78765 -141531
rect -78721 -141575 -78665 -141531
rect -78621 -141575 -78565 -141531
rect -78521 -141575 -78465 -141531
rect -78421 -141575 -78365 -141531
rect -78321 -141575 -78265 -141531
rect -78221 -141575 -78165 -141531
rect -78121 -141575 -78065 -141531
rect -78021 -141575 -77965 -141531
rect -77921 -141575 -77865 -141531
rect -77821 -141575 -77765 -141531
rect -77721 -141575 -77265 -141531
rect -77221 -141575 -77165 -141531
rect -77121 -141575 -77065 -141531
rect -77021 -141575 -76965 -141531
rect -76921 -141575 -76865 -141531
rect -76821 -141575 -76765 -141531
rect -76721 -141575 -76665 -141531
rect -76621 -141575 -76565 -141531
rect -76521 -141575 -76465 -141531
rect -76421 -141575 -76365 -141531
rect -76321 -141575 -76265 -141531
rect -76221 -141575 -76165 -141531
rect -76121 -141575 -76065 -141531
rect -76021 -141575 -75965 -141531
rect -75921 -141575 -75865 -141531
rect -75821 -141575 -75765 -141531
rect -75721 -141575 -72506 -141531
rect -85973 -141631 -72506 -141575
rect -85973 -141675 -83265 -141631
rect -83221 -141675 -83165 -141631
rect -83121 -141675 -83065 -141631
rect -83021 -141675 -82965 -141631
rect -82921 -141675 -82865 -141631
rect -82821 -141675 -82765 -141631
rect -82721 -141675 -82665 -141631
rect -82621 -141675 -82565 -141631
rect -82521 -141675 -82465 -141631
rect -82421 -141675 -82365 -141631
rect -82321 -141675 -82265 -141631
rect -82221 -141675 -82165 -141631
rect -82121 -141675 -82065 -141631
rect -82021 -141675 -81965 -141631
rect -81921 -141675 -81865 -141631
rect -81821 -141675 -81765 -141631
rect -81721 -141675 -81265 -141631
rect -81221 -141675 -81165 -141631
rect -81121 -141675 -81065 -141631
rect -81021 -141675 -80965 -141631
rect -80921 -141675 -80865 -141631
rect -80821 -141675 -80765 -141631
rect -80721 -141675 -80665 -141631
rect -80621 -141675 -80565 -141631
rect -80521 -141675 -80465 -141631
rect -80421 -141675 -80365 -141631
rect -80321 -141675 -80265 -141631
rect -80221 -141675 -80165 -141631
rect -80121 -141675 -80065 -141631
rect -80021 -141675 -79965 -141631
rect -79921 -141675 -79865 -141631
rect -79821 -141675 -79765 -141631
rect -79721 -141675 -79265 -141631
rect -79221 -141675 -79165 -141631
rect -79121 -141675 -79065 -141631
rect -79021 -141675 -78965 -141631
rect -78921 -141675 -78865 -141631
rect -78821 -141675 -78765 -141631
rect -78721 -141675 -78665 -141631
rect -78621 -141675 -78565 -141631
rect -78521 -141675 -78465 -141631
rect -78421 -141675 -78365 -141631
rect -78321 -141675 -78265 -141631
rect -78221 -141675 -78165 -141631
rect -78121 -141675 -78065 -141631
rect -78021 -141675 -77965 -141631
rect -77921 -141675 -77865 -141631
rect -77821 -141675 -77765 -141631
rect -77721 -141675 -77265 -141631
rect -77221 -141675 -77165 -141631
rect -77121 -141675 -77065 -141631
rect -77021 -141675 -76965 -141631
rect -76921 -141675 -76865 -141631
rect -76821 -141675 -76765 -141631
rect -76721 -141675 -76665 -141631
rect -76621 -141675 -76565 -141631
rect -76521 -141675 -76465 -141631
rect -76421 -141675 -76365 -141631
rect -76321 -141675 -76265 -141631
rect -76221 -141675 -76165 -141631
rect -76121 -141675 -76065 -141631
rect -76021 -141675 -75965 -141631
rect -75921 -141675 -75865 -141631
rect -75821 -141675 -75765 -141631
rect -75721 -141675 -72506 -141631
rect -85973 -141731 -72506 -141675
rect -85973 -141775 -83265 -141731
rect -83221 -141775 -83165 -141731
rect -83121 -141775 -83065 -141731
rect -83021 -141775 -82965 -141731
rect -82921 -141775 -82865 -141731
rect -82821 -141775 -82765 -141731
rect -82721 -141775 -82665 -141731
rect -82621 -141775 -82565 -141731
rect -82521 -141775 -82465 -141731
rect -82421 -141775 -82365 -141731
rect -82321 -141775 -82265 -141731
rect -82221 -141775 -82165 -141731
rect -82121 -141775 -82065 -141731
rect -82021 -141775 -81965 -141731
rect -81921 -141775 -81865 -141731
rect -81821 -141775 -81765 -141731
rect -81721 -141775 -81265 -141731
rect -81221 -141775 -81165 -141731
rect -81121 -141775 -81065 -141731
rect -81021 -141775 -80965 -141731
rect -80921 -141775 -80865 -141731
rect -80821 -141775 -80765 -141731
rect -80721 -141775 -80665 -141731
rect -80621 -141775 -80565 -141731
rect -80521 -141775 -80465 -141731
rect -80421 -141775 -80365 -141731
rect -80321 -141775 -80265 -141731
rect -80221 -141775 -80165 -141731
rect -80121 -141775 -80065 -141731
rect -80021 -141775 -79965 -141731
rect -79921 -141775 -79865 -141731
rect -79821 -141775 -79765 -141731
rect -79721 -141775 -79265 -141731
rect -79221 -141775 -79165 -141731
rect -79121 -141775 -79065 -141731
rect -79021 -141775 -78965 -141731
rect -78921 -141775 -78865 -141731
rect -78821 -141775 -78765 -141731
rect -78721 -141775 -78665 -141731
rect -78621 -141775 -78565 -141731
rect -78521 -141775 -78465 -141731
rect -78421 -141775 -78365 -141731
rect -78321 -141775 -78265 -141731
rect -78221 -141775 -78165 -141731
rect -78121 -141775 -78065 -141731
rect -78021 -141775 -77965 -141731
rect -77921 -141775 -77865 -141731
rect -77821 -141775 -77765 -141731
rect -77721 -141775 -77265 -141731
rect -77221 -141775 -77165 -141731
rect -77121 -141775 -77065 -141731
rect -77021 -141775 -76965 -141731
rect -76921 -141775 -76865 -141731
rect -76821 -141775 -76765 -141731
rect -76721 -141775 -76665 -141731
rect -76621 -141775 -76565 -141731
rect -76521 -141775 -76465 -141731
rect -76421 -141775 -76365 -141731
rect -76321 -141775 -76265 -141731
rect -76221 -141775 -76165 -141731
rect -76121 -141775 -76065 -141731
rect -76021 -141775 -75965 -141731
rect -75921 -141775 -75865 -141731
rect -75821 -141775 -75765 -141731
rect -75721 -141775 -72506 -141731
rect -85973 -143750 -72506 -141775
rect -103327 -149974 -79660 -148766
rect -103327 -162685 -97900 -149974
rect -97368 -150681 -97292 -149974
rect -96760 -150681 -96684 -149974
rect -96152 -150681 -96076 -149974
rect -95544 -150681 -95468 -149974
rect -94936 -150681 -94860 -149974
rect -94328 -150681 -94252 -149974
rect -93720 -150681 -93644 -149974
rect -93112 -150681 -93036 -149974
rect -92504 -150681 -92428 -149974
rect -91896 -150681 -91820 -149974
rect -91288 -150681 -91212 -149974
rect -90680 -150681 -90604 -149974
rect -90072 -150681 -89996 -149974
rect -89464 -150681 -89388 -149974
rect -88856 -150681 -88780 -149974
rect -88248 -150681 -88172 -149974
rect -87640 -150681 -87564 -149974
rect -87032 -150681 -86956 -149974
rect -86424 -150681 -86348 -149974
rect -85816 -150681 -85740 -149974
rect -85208 -150681 -85132 -149974
rect -84600 -150681 -84524 -149974
rect -83992 -150681 -83916 -149974
rect -83384 -150681 -83308 -149974
rect -82776 -150681 -82700 -149974
rect -82168 -150681 -82092 -149974
rect -81560 -150681 -81484 -149974
rect -80952 -150681 -80876 -149974
rect -80344 -150681 -80268 -149974
rect -79736 -150681 -79660 -149974
rect -103327 -171279 -98134 -162685
rect -97672 -163392 -97596 -162685
rect -97064 -163392 -96988 -162685
rect -96456 -163392 -96380 -162685
rect -95848 -163392 -95772 -162685
rect -95240 -163392 -95164 -162685
rect -94632 -163392 -94556 -162685
rect -94024 -163392 -93948 -162685
rect -93416 -163392 -93340 -162685
rect -92808 -163392 -92732 -162685
rect -92200 -163392 -92124 -162685
rect -91592 -163392 -91516 -162685
rect -90984 -163392 -90908 -162685
rect -90376 -163392 -90300 -162685
rect -89768 -163392 -89692 -162685
rect -89160 -163392 -89084 -162685
rect -88552 -163392 -88476 -162685
rect -87944 -163392 -87868 -162685
rect -87336 -163392 -87260 -162685
rect -86728 -163392 -86652 -162685
rect -86120 -163392 -86044 -162685
rect -85512 -163392 -85436 -162685
rect -84904 -163392 -84828 -162685
rect -84296 -163392 -84220 -162685
rect -83688 -163392 -83612 -162685
rect -83080 -163392 -83004 -162685
rect -82472 -163392 -82396 -162685
rect -81864 -163392 -81788 -162685
rect -81256 -163392 -81180 -162685
rect -80648 -163392 -80572 -162685
rect -80040 -163392 -79964 -162685
rect -77671 -163392 -72506 -143750
rect -60256 -138310 81632 -138266
rect 81676 -138310 81732 -138266
rect 81776 -138310 81832 -138266
rect 81876 -138310 81932 -138266
rect 81976 -138310 82032 -138266
rect 82076 -138310 82132 -138266
rect 82176 -138310 82232 -138266
rect 82276 -138310 82332 -138266
rect 82376 -138310 82432 -138266
rect 82476 -138310 82532 -138266
rect 82576 -138310 82632 -138266
rect 82676 -138310 82732 -138266
rect 82776 -138310 82832 -138266
rect 82876 -138310 82932 -138266
rect 82976 -138310 83032 -138266
rect 83076 -138310 83132 -138266
rect 83176 -138310 83632 -138266
rect 83676 -138310 83732 -138266
rect 83776 -138310 83832 -138266
rect 83876 -138310 83932 -138266
rect 83976 -138310 84032 -138266
rect 84076 -138310 84132 -138266
rect 84176 -138310 84232 -138266
rect 84276 -138310 84332 -138266
rect 84376 -138310 84432 -138266
rect 84476 -138310 84532 -138266
rect 84576 -138310 84632 -138266
rect 84676 -138310 84732 -138266
rect 84776 -138310 84832 -138266
rect 84876 -138310 84932 -138266
rect 84976 -138310 85032 -138266
rect 85076 -138310 85132 -138266
rect 85176 -138310 85632 -138266
rect 85676 -138310 85732 -138266
rect 85776 -138310 85832 -138266
rect 85876 -138310 85932 -138266
rect 85976 -138310 86032 -138266
rect 86076 -138310 86132 -138266
rect 86176 -138310 86232 -138266
rect 86276 -138310 86332 -138266
rect 86376 -138310 86432 -138266
rect 86476 -138310 86532 -138266
rect 86576 -138310 86632 -138266
rect 86676 -138310 86732 -138266
rect 86776 -138310 86832 -138266
rect 86876 -138310 86932 -138266
rect 86976 -138310 87032 -138266
rect 87076 -138310 87132 -138266
rect 87176 -138310 87632 -138266
rect 87676 -138310 87732 -138266
rect 87776 -138310 87832 -138266
rect 87876 -138310 87932 -138266
rect 87976 -138310 88032 -138266
rect 88076 -138310 88132 -138266
rect 88176 -138310 88232 -138266
rect 88276 -138310 88332 -138266
rect 88376 -138310 88432 -138266
rect 88476 -138310 88532 -138266
rect 88576 -138310 88632 -138266
rect 88676 -138310 88732 -138266
rect 88776 -138310 88832 -138266
rect 88876 -138310 88932 -138266
rect 88976 -138310 89032 -138266
rect 89076 -138310 89132 -138266
rect 89176 -138310 174378 -138266
rect -60256 -138366 174378 -138310
rect -60256 -138410 81632 -138366
rect 81676 -138410 81732 -138366
rect 81776 -138410 81832 -138366
rect 81876 -138410 81932 -138366
rect 81976 -138410 82032 -138366
rect 82076 -138410 82132 -138366
rect 82176 -138410 82232 -138366
rect 82276 -138410 82332 -138366
rect 82376 -138410 82432 -138366
rect 82476 -138410 82532 -138366
rect 82576 -138410 82632 -138366
rect 82676 -138410 82732 -138366
rect 82776 -138410 82832 -138366
rect 82876 -138410 82932 -138366
rect 82976 -138410 83032 -138366
rect 83076 -138410 83132 -138366
rect 83176 -138410 83632 -138366
rect 83676 -138410 83732 -138366
rect 83776 -138410 83832 -138366
rect 83876 -138410 83932 -138366
rect 83976 -138410 84032 -138366
rect 84076 -138410 84132 -138366
rect 84176 -138410 84232 -138366
rect 84276 -138410 84332 -138366
rect 84376 -138410 84432 -138366
rect 84476 -138410 84532 -138366
rect 84576 -138410 84632 -138366
rect 84676 -138410 84732 -138366
rect 84776 -138410 84832 -138366
rect 84876 -138410 84932 -138366
rect 84976 -138410 85032 -138366
rect 85076 -138410 85132 -138366
rect 85176 -138410 85632 -138366
rect 85676 -138410 85732 -138366
rect 85776 -138410 85832 -138366
rect 85876 -138410 85932 -138366
rect 85976 -138410 86032 -138366
rect 86076 -138410 86132 -138366
rect 86176 -138410 86232 -138366
rect 86276 -138410 86332 -138366
rect 86376 -138410 86432 -138366
rect 86476 -138410 86532 -138366
rect 86576 -138410 86632 -138366
rect 86676 -138410 86732 -138366
rect 86776 -138410 86832 -138366
rect 86876 -138410 86932 -138366
rect 86976 -138410 87032 -138366
rect 87076 -138410 87132 -138366
rect 87176 -138410 87632 -138366
rect 87676 -138410 87732 -138366
rect 87776 -138410 87832 -138366
rect 87876 -138410 87932 -138366
rect 87976 -138410 88032 -138366
rect 88076 -138410 88132 -138366
rect 88176 -138410 88232 -138366
rect 88276 -138410 88332 -138366
rect 88376 -138410 88432 -138366
rect 88476 -138410 88532 -138366
rect 88576 -138410 88632 -138366
rect 88676 -138410 88732 -138366
rect 88776 -138410 88832 -138366
rect 88876 -138410 88932 -138366
rect 88976 -138410 89032 -138366
rect 89076 -138410 89132 -138366
rect 89176 -138410 174378 -138366
rect -60256 -138466 174378 -138410
rect -60256 -138510 81632 -138466
rect 81676 -138510 81732 -138466
rect 81776 -138510 81832 -138466
rect 81876 -138510 81932 -138466
rect 81976 -138510 82032 -138466
rect 82076 -138510 82132 -138466
rect 82176 -138510 82232 -138466
rect 82276 -138510 82332 -138466
rect 82376 -138510 82432 -138466
rect 82476 -138510 82532 -138466
rect 82576 -138510 82632 -138466
rect 82676 -138510 82732 -138466
rect 82776 -138510 82832 -138466
rect 82876 -138510 82932 -138466
rect 82976 -138510 83032 -138466
rect 83076 -138510 83132 -138466
rect 83176 -138510 83632 -138466
rect 83676 -138510 83732 -138466
rect 83776 -138510 83832 -138466
rect 83876 -138510 83932 -138466
rect 83976 -138510 84032 -138466
rect 84076 -138510 84132 -138466
rect 84176 -138510 84232 -138466
rect 84276 -138510 84332 -138466
rect 84376 -138510 84432 -138466
rect 84476 -138510 84532 -138466
rect 84576 -138510 84632 -138466
rect 84676 -138510 84732 -138466
rect 84776 -138510 84832 -138466
rect 84876 -138510 84932 -138466
rect 84976 -138510 85032 -138466
rect 85076 -138510 85132 -138466
rect 85176 -138510 85632 -138466
rect 85676 -138510 85732 -138466
rect 85776 -138510 85832 -138466
rect 85876 -138510 85932 -138466
rect 85976 -138510 86032 -138466
rect 86076 -138510 86132 -138466
rect 86176 -138510 86232 -138466
rect 86276 -138510 86332 -138466
rect 86376 -138510 86432 -138466
rect 86476 -138510 86532 -138466
rect 86576 -138510 86632 -138466
rect 86676 -138510 86732 -138466
rect 86776 -138510 86832 -138466
rect 86876 -138510 86932 -138466
rect 86976 -138510 87032 -138466
rect 87076 -138510 87132 -138466
rect 87176 -138510 87632 -138466
rect 87676 -138510 87732 -138466
rect 87776 -138510 87832 -138466
rect 87876 -138510 87932 -138466
rect 87976 -138510 88032 -138466
rect 88076 -138510 88132 -138466
rect 88176 -138510 88232 -138466
rect 88276 -138510 88332 -138466
rect 88376 -138510 88432 -138466
rect 88476 -138510 88532 -138466
rect 88576 -138510 88632 -138466
rect 88676 -138510 88732 -138466
rect 88776 -138510 88832 -138466
rect 88876 -138510 88932 -138466
rect 88976 -138510 89032 -138466
rect 89076 -138510 89132 -138466
rect 89176 -138510 174378 -138466
rect -60256 -138566 174378 -138510
rect -60256 -138610 81632 -138566
rect 81676 -138610 81732 -138566
rect 81776 -138610 81832 -138566
rect 81876 -138610 81932 -138566
rect 81976 -138610 82032 -138566
rect 82076 -138610 82132 -138566
rect 82176 -138610 82232 -138566
rect 82276 -138610 82332 -138566
rect 82376 -138610 82432 -138566
rect 82476 -138610 82532 -138566
rect 82576 -138610 82632 -138566
rect 82676 -138610 82732 -138566
rect 82776 -138610 82832 -138566
rect 82876 -138610 82932 -138566
rect 82976 -138610 83032 -138566
rect 83076 -138610 83132 -138566
rect 83176 -138610 83632 -138566
rect 83676 -138610 83732 -138566
rect 83776 -138610 83832 -138566
rect 83876 -138610 83932 -138566
rect 83976 -138610 84032 -138566
rect 84076 -138610 84132 -138566
rect 84176 -138610 84232 -138566
rect 84276 -138610 84332 -138566
rect 84376 -138610 84432 -138566
rect 84476 -138610 84532 -138566
rect 84576 -138610 84632 -138566
rect 84676 -138610 84732 -138566
rect 84776 -138610 84832 -138566
rect 84876 -138610 84932 -138566
rect 84976 -138610 85032 -138566
rect 85076 -138610 85132 -138566
rect 85176 -138610 85632 -138566
rect 85676 -138610 85732 -138566
rect 85776 -138610 85832 -138566
rect 85876 -138610 85932 -138566
rect 85976 -138610 86032 -138566
rect 86076 -138610 86132 -138566
rect 86176 -138610 86232 -138566
rect 86276 -138610 86332 -138566
rect 86376 -138610 86432 -138566
rect 86476 -138610 86532 -138566
rect 86576 -138610 86632 -138566
rect 86676 -138610 86732 -138566
rect 86776 -138610 86832 -138566
rect 86876 -138610 86932 -138566
rect 86976 -138610 87032 -138566
rect 87076 -138610 87132 -138566
rect 87176 -138610 87632 -138566
rect 87676 -138610 87732 -138566
rect 87776 -138610 87832 -138566
rect 87876 -138610 87932 -138566
rect 87976 -138610 88032 -138566
rect 88076 -138610 88132 -138566
rect 88176 -138610 88232 -138566
rect 88276 -138610 88332 -138566
rect 88376 -138610 88432 -138566
rect 88476 -138610 88532 -138566
rect 88576 -138610 88632 -138566
rect 88676 -138610 88732 -138566
rect 88776 -138610 88832 -138566
rect 88876 -138610 88932 -138566
rect 88976 -138610 89032 -138566
rect 89076 -138610 89132 -138566
rect 89176 -138610 174378 -138566
rect -60256 -138666 174378 -138610
rect -60256 -138710 81632 -138666
rect 81676 -138710 81732 -138666
rect 81776 -138710 81832 -138666
rect 81876 -138710 81932 -138666
rect 81976 -138710 82032 -138666
rect 82076 -138710 82132 -138666
rect 82176 -138710 82232 -138666
rect 82276 -138710 82332 -138666
rect 82376 -138710 82432 -138666
rect 82476 -138710 82532 -138666
rect 82576 -138710 82632 -138666
rect 82676 -138710 82732 -138666
rect 82776 -138710 82832 -138666
rect 82876 -138710 82932 -138666
rect 82976 -138710 83032 -138666
rect 83076 -138710 83132 -138666
rect 83176 -138710 83632 -138666
rect 83676 -138710 83732 -138666
rect 83776 -138710 83832 -138666
rect 83876 -138710 83932 -138666
rect 83976 -138710 84032 -138666
rect 84076 -138710 84132 -138666
rect 84176 -138710 84232 -138666
rect 84276 -138710 84332 -138666
rect 84376 -138710 84432 -138666
rect 84476 -138710 84532 -138666
rect 84576 -138710 84632 -138666
rect 84676 -138710 84732 -138666
rect 84776 -138710 84832 -138666
rect 84876 -138710 84932 -138666
rect 84976 -138710 85032 -138666
rect 85076 -138710 85132 -138666
rect 85176 -138710 85632 -138666
rect 85676 -138710 85732 -138666
rect 85776 -138710 85832 -138666
rect 85876 -138710 85932 -138666
rect 85976 -138710 86032 -138666
rect 86076 -138710 86132 -138666
rect 86176 -138710 86232 -138666
rect 86276 -138710 86332 -138666
rect 86376 -138710 86432 -138666
rect 86476 -138710 86532 -138666
rect 86576 -138710 86632 -138666
rect 86676 -138710 86732 -138666
rect 86776 -138710 86832 -138666
rect 86876 -138710 86932 -138666
rect 86976 -138710 87032 -138666
rect 87076 -138710 87132 -138666
rect 87176 -138710 87632 -138666
rect 87676 -138710 87732 -138666
rect 87776 -138710 87832 -138666
rect 87876 -138710 87932 -138666
rect 87976 -138710 88032 -138666
rect 88076 -138710 88132 -138666
rect 88176 -138710 88232 -138666
rect 88276 -138710 88332 -138666
rect 88376 -138710 88432 -138666
rect 88476 -138710 88532 -138666
rect 88576 -138710 88632 -138666
rect 88676 -138710 88732 -138666
rect 88776 -138710 88832 -138666
rect 88876 -138710 88932 -138666
rect 88976 -138710 89032 -138666
rect 89076 -138710 89132 -138666
rect 89176 -138710 174378 -138666
rect -60256 -138766 174378 -138710
rect -60256 -138810 81632 -138766
rect 81676 -138810 81732 -138766
rect 81776 -138810 81832 -138766
rect 81876 -138810 81932 -138766
rect 81976 -138810 82032 -138766
rect 82076 -138810 82132 -138766
rect 82176 -138810 82232 -138766
rect 82276 -138810 82332 -138766
rect 82376 -138810 82432 -138766
rect 82476 -138810 82532 -138766
rect 82576 -138810 82632 -138766
rect 82676 -138810 82732 -138766
rect 82776 -138810 82832 -138766
rect 82876 -138810 82932 -138766
rect 82976 -138810 83032 -138766
rect 83076 -138810 83132 -138766
rect 83176 -138810 83632 -138766
rect 83676 -138810 83732 -138766
rect 83776 -138810 83832 -138766
rect 83876 -138810 83932 -138766
rect 83976 -138810 84032 -138766
rect 84076 -138810 84132 -138766
rect 84176 -138810 84232 -138766
rect 84276 -138810 84332 -138766
rect 84376 -138810 84432 -138766
rect 84476 -138810 84532 -138766
rect 84576 -138810 84632 -138766
rect 84676 -138810 84732 -138766
rect 84776 -138810 84832 -138766
rect 84876 -138810 84932 -138766
rect 84976 -138810 85032 -138766
rect 85076 -138810 85132 -138766
rect 85176 -138810 85632 -138766
rect 85676 -138810 85732 -138766
rect 85776 -138810 85832 -138766
rect 85876 -138810 85932 -138766
rect 85976 -138810 86032 -138766
rect 86076 -138810 86132 -138766
rect 86176 -138810 86232 -138766
rect 86276 -138810 86332 -138766
rect 86376 -138810 86432 -138766
rect 86476 -138810 86532 -138766
rect 86576 -138810 86632 -138766
rect 86676 -138810 86732 -138766
rect 86776 -138810 86832 -138766
rect 86876 -138810 86932 -138766
rect 86976 -138810 87032 -138766
rect 87076 -138810 87132 -138766
rect 87176 -138810 87632 -138766
rect 87676 -138810 87732 -138766
rect 87776 -138810 87832 -138766
rect 87876 -138810 87932 -138766
rect 87976 -138810 88032 -138766
rect 88076 -138810 88132 -138766
rect 88176 -138810 88232 -138766
rect 88276 -138810 88332 -138766
rect 88376 -138810 88432 -138766
rect 88476 -138810 88532 -138766
rect 88576 -138810 88632 -138766
rect 88676 -138810 88732 -138766
rect 88776 -138810 88832 -138766
rect 88876 -138810 88932 -138766
rect 88976 -138810 89032 -138766
rect 89076 -138810 89132 -138766
rect 89176 -138810 174378 -138766
rect -60256 -138866 174378 -138810
rect -60256 -138910 81632 -138866
rect 81676 -138910 81732 -138866
rect 81776 -138910 81832 -138866
rect 81876 -138910 81932 -138866
rect 81976 -138910 82032 -138866
rect 82076 -138910 82132 -138866
rect 82176 -138910 82232 -138866
rect 82276 -138910 82332 -138866
rect 82376 -138910 82432 -138866
rect 82476 -138910 82532 -138866
rect 82576 -138910 82632 -138866
rect 82676 -138910 82732 -138866
rect 82776 -138910 82832 -138866
rect 82876 -138910 82932 -138866
rect 82976 -138910 83032 -138866
rect 83076 -138910 83132 -138866
rect 83176 -138910 83632 -138866
rect 83676 -138910 83732 -138866
rect 83776 -138910 83832 -138866
rect 83876 -138910 83932 -138866
rect 83976 -138910 84032 -138866
rect 84076 -138910 84132 -138866
rect 84176 -138910 84232 -138866
rect 84276 -138910 84332 -138866
rect 84376 -138910 84432 -138866
rect 84476 -138910 84532 -138866
rect 84576 -138910 84632 -138866
rect 84676 -138910 84732 -138866
rect 84776 -138910 84832 -138866
rect 84876 -138910 84932 -138866
rect 84976 -138910 85032 -138866
rect 85076 -138910 85132 -138866
rect 85176 -138910 85632 -138866
rect 85676 -138910 85732 -138866
rect 85776 -138910 85832 -138866
rect 85876 -138910 85932 -138866
rect 85976 -138910 86032 -138866
rect 86076 -138910 86132 -138866
rect 86176 -138910 86232 -138866
rect 86276 -138910 86332 -138866
rect 86376 -138910 86432 -138866
rect 86476 -138910 86532 -138866
rect 86576 -138910 86632 -138866
rect 86676 -138910 86732 -138866
rect 86776 -138910 86832 -138866
rect 86876 -138910 86932 -138866
rect 86976 -138910 87032 -138866
rect 87076 -138910 87132 -138866
rect 87176 -138910 87632 -138866
rect 87676 -138910 87732 -138866
rect 87776 -138910 87832 -138866
rect 87876 -138910 87932 -138866
rect 87976 -138910 88032 -138866
rect 88076 -138910 88132 -138866
rect 88176 -138910 88232 -138866
rect 88276 -138910 88332 -138866
rect 88376 -138910 88432 -138866
rect 88476 -138910 88532 -138866
rect 88576 -138910 88632 -138866
rect 88676 -138910 88732 -138866
rect 88776 -138910 88832 -138866
rect 88876 -138910 88932 -138866
rect 88976 -138910 89032 -138866
rect 89076 -138910 89132 -138866
rect 89176 -138910 174378 -138866
rect -60256 -138966 174378 -138910
rect -60256 -139010 81632 -138966
rect 81676 -139010 81732 -138966
rect 81776 -139010 81832 -138966
rect 81876 -139010 81932 -138966
rect 81976 -139010 82032 -138966
rect 82076 -139010 82132 -138966
rect 82176 -139010 82232 -138966
rect 82276 -139010 82332 -138966
rect 82376 -139010 82432 -138966
rect 82476 -139010 82532 -138966
rect 82576 -139010 82632 -138966
rect 82676 -139010 82732 -138966
rect 82776 -139010 82832 -138966
rect 82876 -139010 82932 -138966
rect 82976 -139010 83032 -138966
rect 83076 -139010 83132 -138966
rect 83176 -139010 83632 -138966
rect 83676 -139010 83732 -138966
rect 83776 -139010 83832 -138966
rect 83876 -139010 83932 -138966
rect 83976 -139010 84032 -138966
rect 84076 -139010 84132 -138966
rect 84176 -139010 84232 -138966
rect 84276 -139010 84332 -138966
rect 84376 -139010 84432 -138966
rect 84476 -139010 84532 -138966
rect 84576 -139010 84632 -138966
rect 84676 -139010 84732 -138966
rect 84776 -139010 84832 -138966
rect 84876 -139010 84932 -138966
rect 84976 -139010 85032 -138966
rect 85076 -139010 85132 -138966
rect 85176 -139010 85632 -138966
rect 85676 -139010 85732 -138966
rect 85776 -139010 85832 -138966
rect 85876 -139010 85932 -138966
rect 85976 -139010 86032 -138966
rect 86076 -139010 86132 -138966
rect 86176 -139010 86232 -138966
rect 86276 -139010 86332 -138966
rect 86376 -139010 86432 -138966
rect 86476 -139010 86532 -138966
rect 86576 -139010 86632 -138966
rect 86676 -139010 86732 -138966
rect 86776 -139010 86832 -138966
rect 86876 -139010 86932 -138966
rect 86976 -139010 87032 -138966
rect 87076 -139010 87132 -138966
rect 87176 -139010 87632 -138966
rect 87676 -139010 87732 -138966
rect 87776 -139010 87832 -138966
rect 87876 -139010 87932 -138966
rect 87976 -139010 88032 -138966
rect 88076 -139010 88132 -138966
rect 88176 -139010 88232 -138966
rect 88276 -139010 88332 -138966
rect 88376 -139010 88432 -138966
rect 88476 -139010 88532 -138966
rect 88576 -139010 88632 -138966
rect 88676 -139010 88732 -138966
rect 88776 -139010 88832 -138966
rect 88876 -139010 88932 -138966
rect 88976 -139010 89032 -138966
rect 89076 -139010 89132 -138966
rect 89176 -139010 174378 -138966
rect -60256 -139066 174378 -139010
rect -60256 -139110 81632 -139066
rect 81676 -139110 81732 -139066
rect 81776 -139110 81832 -139066
rect 81876 -139110 81932 -139066
rect 81976 -139110 82032 -139066
rect 82076 -139110 82132 -139066
rect 82176 -139110 82232 -139066
rect 82276 -139110 82332 -139066
rect 82376 -139110 82432 -139066
rect 82476 -139110 82532 -139066
rect 82576 -139110 82632 -139066
rect 82676 -139110 82732 -139066
rect 82776 -139110 82832 -139066
rect 82876 -139110 82932 -139066
rect 82976 -139110 83032 -139066
rect 83076 -139110 83132 -139066
rect 83176 -139110 83632 -139066
rect 83676 -139110 83732 -139066
rect 83776 -139110 83832 -139066
rect 83876 -139110 83932 -139066
rect 83976 -139110 84032 -139066
rect 84076 -139110 84132 -139066
rect 84176 -139110 84232 -139066
rect 84276 -139110 84332 -139066
rect 84376 -139110 84432 -139066
rect 84476 -139110 84532 -139066
rect 84576 -139110 84632 -139066
rect 84676 -139110 84732 -139066
rect 84776 -139110 84832 -139066
rect 84876 -139110 84932 -139066
rect 84976 -139110 85032 -139066
rect 85076 -139110 85132 -139066
rect 85176 -139110 85632 -139066
rect 85676 -139110 85732 -139066
rect 85776 -139110 85832 -139066
rect 85876 -139110 85932 -139066
rect 85976 -139110 86032 -139066
rect 86076 -139110 86132 -139066
rect 86176 -139110 86232 -139066
rect 86276 -139110 86332 -139066
rect 86376 -139110 86432 -139066
rect 86476 -139110 86532 -139066
rect 86576 -139110 86632 -139066
rect 86676 -139110 86732 -139066
rect 86776 -139110 86832 -139066
rect 86876 -139110 86932 -139066
rect 86976 -139110 87032 -139066
rect 87076 -139110 87132 -139066
rect 87176 -139110 87632 -139066
rect 87676 -139110 87732 -139066
rect 87776 -139110 87832 -139066
rect 87876 -139110 87932 -139066
rect 87976 -139110 88032 -139066
rect 88076 -139110 88132 -139066
rect 88176 -139110 88232 -139066
rect 88276 -139110 88332 -139066
rect 88376 -139110 88432 -139066
rect 88476 -139110 88532 -139066
rect 88576 -139110 88632 -139066
rect 88676 -139110 88732 -139066
rect 88776 -139110 88832 -139066
rect 88876 -139110 88932 -139066
rect 88976 -139110 89032 -139066
rect 89076 -139110 89132 -139066
rect 89176 -139110 174378 -139066
rect -60256 -139166 174378 -139110
rect -60256 -139210 81632 -139166
rect 81676 -139210 81732 -139166
rect 81776 -139210 81832 -139166
rect 81876 -139210 81932 -139166
rect 81976 -139210 82032 -139166
rect 82076 -139210 82132 -139166
rect 82176 -139210 82232 -139166
rect 82276 -139210 82332 -139166
rect 82376 -139210 82432 -139166
rect 82476 -139210 82532 -139166
rect 82576 -139210 82632 -139166
rect 82676 -139210 82732 -139166
rect 82776 -139210 82832 -139166
rect 82876 -139210 82932 -139166
rect 82976 -139210 83032 -139166
rect 83076 -139210 83132 -139166
rect 83176 -139210 83632 -139166
rect 83676 -139210 83732 -139166
rect 83776 -139210 83832 -139166
rect 83876 -139210 83932 -139166
rect 83976 -139210 84032 -139166
rect 84076 -139210 84132 -139166
rect 84176 -139210 84232 -139166
rect 84276 -139210 84332 -139166
rect 84376 -139210 84432 -139166
rect 84476 -139210 84532 -139166
rect 84576 -139210 84632 -139166
rect 84676 -139210 84732 -139166
rect 84776 -139210 84832 -139166
rect 84876 -139210 84932 -139166
rect 84976 -139210 85032 -139166
rect 85076 -139210 85132 -139166
rect 85176 -139210 85632 -139166
rect 85676 -139210 85732 -139166
rect 85776 -139210 85832 -139166
rect 85876 -139210 85932 -139166
rect 85976 -139210 86032 -139166
rect 86076 -139210 86132 -139166
rect 86176 -139210 86232 -139166
rect 86276 -139210 86332 -139166
rect 86376 -139210 86432 -139166
rect 86476 -139210 86532 -139166
rect 86576 -139210 86632 -139166
rect 86676 -139210 86732 -139166
rect 86776 -139210 86832 -139166
rect 86876 -139210 86932 -139166
rect 86976 -139210 87032 -139166
rect 87076 -139210 87132 -139166
rect 87176 -139210 87632 -139166
rect 87676 -139210 87732 -139166
rect 87776 -139210 87832 -139166
rect 87876 -139210 87932 -139166
rect 87976 -139210 88032 -139166
rect 88076 -139210 88132 -139166
rect 88176 -139210 88232 -139166
rect 88276 -139210 88332 -139166
rect 88376 -139210 88432 -139166
rect 88476 -139210 88532 -139166
rect 88576 -139210 88632 -139166
rect 88676 -139210 88732 -139166
rect 88776 -139210 88832 -139166
rect 88876 -139210 88932 -139166
rect 88976 -139210 89032 -139166
rect 89076 -139210 89132 -139166
rect 89176 -139210 174378 -139166
rect -60256 -139266 174378 -139210
rect -60256 -139310 81632 -139266
rect 81676 -139310 81732 -139266
rect 81776 -139310 81832 -139266
rect 81876 -139310 81932 -139266
rect 81976 -139310 82032 -139266
rect 82076 -139310 82132 -139266
rect 82176 -139310 82232 -139266
rect 82276 -139310 82332 -139266
rect 82376 -139310 82432 -139266
rect 82476 -139310 82532 -139266
rect 82576 -139310 82632 -139266
rect 82676 -139310 82732 -139266
rect 82776 -139310 82832 -139266
rect 82876 -139310 82932 -139266
rect 82976 -139310 83032 -139266
rect 83076 -139310 83132 -139266
rect 83176 -139310 83632 -139266
rect 83676 -139310 83732 -139266
rect 83776 -139310 83832 -139266
rect 83876 -139310 83932 -139266
rect 83976 -139310 84032 -139266
rect 84076 -139310 84132 -139266
rect 84176 -139310 84232 -139266
rect 84276 -139310 84332 -139266
rect 84376 -139310 84432 -139266
rect 84476 -139310 84532 -139266
rect 84576 -139310 84632 -139266
rect 84676 -139310 84732 -139266
rect 84776 -139310 84832 -139266
rect 84876 -139310 84932 -139266
rect 84976 -139310 85032 -139266
rect 85076 -139310 85132 -139266
rect 85176 -139310 85632 -139266
rect 85676 -139310 85732 -139266
rect 85776 -139310 85832 -139266
rect 85876 -139310 85932 -139266
rect 85976 -139310 86032 -139266
rect 86076 -139310 86132 -139266
rect 86176 -139310 86232 -139266
rect 86276 -139310 86332 -139266
rect 86376 -139310 86432 -139266
rect 86476 -139310 86532 -139266
rect 86576 -139310 86632 -139266
rect 86676 -139310 86732 -139266
rect 86776 -139310 86832 -139266
rect 86876 -139310 86932 -139266
rect 86976 -139310 87032 -139266
rect 87076 -139310 87132 -139266
rect 87176 -139310 87632 -139266
rect 87676 -139310 87732 -139266
rect 87776 -139310 87832 -139266
rect 87876 -139310 87932 -139266
rect 87976 -139310 88032 -139266
rect 88076 -139310 88132 -139266
rect 88176 -139310 88232 -139266
rect 88276 -139310 88332 -139266
rect 88376 -139310 88432 -139266
rect 88476 -139310 88532 -139266
rect 88576 -139310 88632 -139266
rect 88676 -139310 88732 -139266
rect 88776 -139310 88832 -139266
rect 88876 -139310 88932 -139266
rect 88976 -139310 89032 -139266
rect 89076 -139310 89132 -139266
rect 89176 -139310 174378 -139266
rect -60256 -139366 174378 -139310
rect -60256 -139410 81632 -139366
rect 81676 -139410 81732 -139366
rect 81776 -139410 81832 -139366
rect 81876 -139410 81932 -139366
rect 81976 -139410 82032 -139366
rect 82076 -139410 82132 -139366
rect 82176 -139410 82232 -139366
rect 82276 -139410 82332 -139366
rect 82376 -139410 82432 -139366
rect 82476 -139410 82532 -139366
rect 82576 -139410 82632 -139366
rect 82676 -139410 82732 -139366
rect 82776 -139410 82832 -139366
rect 82876 -139410 82932 -139366
rect 82976 -139410 83032 -139366
rect 83076 -139410 83132 -139366
rect 83176 -139410 83632 -139366
rect 83676 -139410 83732 -139366
rect 83776 -139410 83832 -139366
rect 83876 -139410 83932 -139366
rect 83976 -139410 84032 -139366
rect 84076 -139410 84132 -139366
rect 84176 -139410 84232 -139366
rect 84276 -139410 84332 -139366
rect 84376 -139410 84432 -139366
rect 84476 -139410 84532 -139366
rect 84576 -139410 84632 -139366
rect 84676 -139410 84732 -139366
rect 84776 -139410 84832 -139366
rect 84876 -139410 84932 -139366
rect 84976 -139410 85032 -139366
rect 85076 -139410 85132 -139366
rect 85176 -139410 85632 -139366
rect 85676 -139410 85732 -139366
rect 85776 -139410 85832 -139366
rect 85876 -139410 85932 -139366
rect 85976 -139410 86032 -139366
rect 86076 -139410 86132 -139366
rect 86176 -139410 86232 -139366
rect 86276 -139410 86332 -139366
rect 86376 -139410 86432 -139366
rect 86476 -139410 86532 -139366
rect 86576 -139410 86632 -139366
rect 86676 -139410 86732 -139366
rect 86776 -139410 86832 -139366
rect 86876 -139410 86932 -139366
rect 86976 -139410 87032 -139366
rect 87076 -139410 87132 -139366
rect 87176 -139410 87632 -139366
rect 87676 -139410 87732 -139366
rect 87776 -139410 87832 -139366
rect 87876 -139410 87932 -139366
rect 87976 -139410 88032 -139366
rect 88076 -139410 88132 -139366
rect 88176 -139410 88232 -139366
rect 88276 -139410 88332 -139366
rect 88376 -139410 88432 -139366
rect 88476 -139410 88532 -139366
rect 88576 -139410 88632 -139366
rect 88676 -139410 88732 -139366
rect 88776 -139410 88832 -139366
rect 88876 -139410 88932 -139366
rect 88976 -139410 89032 -139366
rect 89076 -139410 89132 -139366
rect 89176 -139410 174378 -139366
rect -60256 -139466 174378 -139410
rect -60256 -139510 81632 -139466
rect 81676 -139510 81732 -139466
rect 81776 -139510 81832 -139466
rect 81876 -139510 81932 -139466
rect 81976 -139510 82032 -139466
rect 82076 -139510 82132 -139466
rect 82176 -139510 82232 -139466
rect 82276 -139510 82332 -139466
rect 82376 -139510 82432 -139466
rect 82476 -139510 82532 -139466
rect 82576 -139510 82632 -139466
rect 82676 -139510 82732 -139466
rect 82776 -139510 82832 -139466
rect 82876 -139510 82932 -139466
rect 82976 -139510 83032 -139466
rect 83076 -139510 83132 -139466
rect 83176 -139510 83632 -139466
rect 83676 -139510 83732 -139466
rect 83776 -139510 83832 -139466
rect 83876 -139510 83932 -139466
rect 83976 -139510 84032 -139466
rect 84076 -139510 84132 -139466
rect 84176 -139510 84232 -139466
rect 84276 -139510 84332 -139466
rect 84376 -139510 84432 -139466
rect 84476 -139510 84532 -139466
rect 84576 -139510 84632 -139466
rect 84676 -139510 84732 -139466
rect 84776 -139510 84832 -139466
rect 84876 -139510 84932 -139466
rect 84976 -139510 85032 -139466
rect 85076 -139510 85132 -139466
rect 85176 -139510 85632 -139466
rect 85676 -139510 85732 -139466
rect 85776 -139510 85832 -139466
rect 85876 -139510 85932 -139466
rect 85976 -139510 86032 -139466
rect 86076 -139510 86132 -139466
rect 86176 -139510 86232 -139466
rect 86276 -139510 86332 -139466
rect 86376 -139510 86432 -139466
rect 86476 -139510 86532 -139466
rect 86576 -139510 86632 -139466
rect 86676 -139510 86732 -139466
rect 86776 -139510 86832 -139466
rect 86876 -139510 86932 -139466
rect 86976 -139510 87032 -139466
rect 87076 -139510 87132 -139466
rect 87176 -139510 87632 -139466
rect 87676 -139510 87732 -139466
rect 87776 -139510 87832 -139466
rect 87876 -139510 87932 -139466
rect 87976 -139510 88032 -139466
rect 88076 -139510 88132 -139466
rect 88176 -139510 88232 -139466
rect 88276 -139510 88332 -139466
rect 88376 -139510 88432 -139466
rect 88476 -139510 88532 -139466
rect 88576 -139510 88632 -139466
rect 88676 -139510 88732 -139466
rect 88776 -139510 88832 -139466
rect 88876 -139510 88932 -139466
rect 88976 -139510 89032 -139466
rect 89076 -139510 89132 -139466
rect 89176 -139510 174378 -139466
rect -60256 -141107 174378 -139510
rect -60256 -162352 -60022 -141107
rect -59490 -142350 -59414 -141107
rect -58882 -142350 -58806 -141107
rect -58274 -142350 -58198 -141107
rect -57666 -142350 -57590 -141107
rect -57058 -142350 -56982 -141107
rect -56450 -142350 -56374 -141107
rect -55842 -142350 -55766 -141107
rect -55234 -142350 -55158 -141107
rect -54626 -142350 -54550 -141107
rect -54018 -142350 -53942 -141107
rect -53410 -142350 -53334 -141107
rect -52802 -142350 -52726 -141107
rect -52194 -142350 -52118 -141107
rect -51586 -142350 -51510 -141107
rect -50978 -142350 -50902 -141107
rect -50370 -142350 -50294 -141107
rect -49762 -142350 -49686 -141107
rect -49154 -142350 -49078 -141107
rect -48546 -142350 -48470 -141107
rect -47938 -142350 -47862 -141107
rect -47330 -142350 -47254 -141107
rect -46722 -142350 -46646 -141107
rect -46114 -142350 -46038 -141107
rect -45506 -142350 -45430 -141107
rect -44898 -142350 -44822 -141107
rect -44290 -142350 -44214 -141107
rect -43682 -142350 -43606 -141107
rect -43074 -142350 -42998 -141107
rect -42466 -142350 -42390 -141107
rect -41858 -142350 -41782 -141107
rect -41250 -142350 -41174 -141107
rect -40642 -142350 -40566 -141107
rect -40034 -142350 -39958 -141107
rect -39426 -142350 -39350 -141107
rect -38818 -142350 -38742 -141107
rect -38210 -142350 -38134 -141107
rect -37602 -142350 -37526 -141107
rect -36994 -142350 -36918 -141107
rect -36386 -142350 -36310 -141107
rect -35778 -142350 -35702 -141107
rect -35170 -142350 -35094 -141107
rect -34562 -142350 -34486 -141107
rect -33954 -142350 -33878 -141107
rect -33346 -142350 -33270 -141107
rect -32738 -142350 -32662 -141107
rect -32130 -142350 -32054 -141107
rect -31522 -142350 -31446 -141107
rect -30914 -142350 -30838 -141107
rect -30306 -142350 -30230 -141107
rect -29698 -142350 -29622 -141107
rect -26256 -162352 -26022 -141107
rect -25490 -142350 -25414 -141107
rect -24882 -142350 -24806 -141107
rect -24274 -142350 -24198 -141107
rect -23666 -142350 -23590 -141107
rect -23058 -142350 -22982 -141107
rect -22450 -142350 -22374 -141107
rect -21842 -142350 -21766 -141107
rect -21234 -142350 -21158 -141107
rect -20626 -142350 -20550 -141107
rect -20018 -142350 -19942 -141107
rect -19410 -142350 -19334 -141107
rect -18802 -142350 -18726 -141107
rect -18194 -142350 -18118 -141107
rect -17586 -142350 -17510 -141107
rect -16978 -142350 -16902 -141107
rect -16370 -142350 -16294 -141107
rect -15762 -142350 -15686 -141107
rect -15154 -142350 -15078 -141107
rect -14546 -142350 -14470 -141107
rect -13938 -142350 -13862 -141107
rect -13330 -142350 -13254 -141107
rect -12722 -142350 -12646 -141107
rect -12114 -142350 -12038 -141107
rect -11506 -142350 -11430 -141107
rect -10898 -142350 -10822 -141107
rect -10290 -142350 -10214 -141107
rect -9682 -142350 -9606 -141107
rect -9074 -142350 -8998 -141107
rect -8466 -142350 -8390 -141107
rect -7858 -142350 -7782 -141107
rect -7250 -142350 -7174 -141107
rect -6642 -142350 -6566 -141107
rect -6034 -142350 -5958 -141107
rect -5426 -142350 -5350 -141107
rect -4818 -142350 -4742 -141107
rect -4210 -142350 -4134 -141107
rect -3602 -142350 -3526 -141107
rect -2994 -142350 -2918 -141107
rect -2386 -142350 -2310 -141107
rect -1778 -142350 -1702 -141107
rect -1170 -142350 -1094 -141107
rect -562 -142350 -486 -141107
rect 46 -142350 122 -141107
rect 654 -142350 730 -141107
rect 1262 -142350 1338 -141107
rect 1870 -142350 1946 -141107
rect 2478 -142350 2554 -141107
rect 3086 -142350 3162 -141107
rect 3694 -142350 3770 -141107
rect 4302 -142350 4378 -141107
rect 7744 -162352 7978 -141107
rect 8510 -142350 8586 -141107
rect 9118 -142350 9194 -141107
rect 9726 -142350 9802 -141107
rect 10334 -142350 10410 -141107
rect 10942 -142350 11018 -141107
rect 11550 -142350 11626 -141107
rect 12158 -142350 12234 -141107
rect 12766 -142350 12842 -141107
rect 13374 -142350 13450 -141107
rect 13982 -142350 14058 -141107
rect 14590 -142350 14666 -141107
rect 15198 -142350 15274 -141107
rect 15806 -142350 15882 -141107
rect 16414 -142350 16490 -141107
rect 17022 -142350 17098 -141107
rect 17630 -142350 17706 -141107
rect 18238 -142350 18314 -141107
rect 18846 -142350 18922 -141107
rect 19454 -142350 19530 -141107
rect 20062 -142350 20138 -141107
rect 20670 -142350 20746 -141107
rect 21278 -142350 21354 -141107
rect 21886 -142350 21962 -141107
rect 22494 -142350 22570 -141107
rect 23102 -142350 23178 -141107
rect 23710 -142350 23786 -141107
rect 24318 -142350 24394 -141107
rect 24926 -142350 25002 -141107
rect 25534 -142350 25610 -141107
rect 26142 -142350 26218 -141107
rect 26750 -142350 26826 -141107
rect 27358 -142350 27434 -141107
rect 27966 -142350 28042 -141107
rect 28574 -142350 28650 -141107
rect 29182 -142350 29258 -141107
rect 29790 -142350 29866 -141107
rect 30398 -142350 30474 -141107
rect 31006 -142350 31082 -141107
rect 31614 -142350 31690 -141107
rect 32222 -142350 32298 -141107
rect 32830 -142350 32906 -141107
rect 33438 -142350 33514 -141107
rect 34046 -142350 34122 -141107
rect 34654 -142350 34730 -141107
rect 35262 -142350 35338 -141107
rect 35870 -142350 35946 -141107
rect 36478 -142350 36554 -141107
rect 37086 -142350 37162 -141107
rect 37694 -142350 37770 -141107
rect 38302 -142350 38378 -141107
rect 41744 -162352 41978 -141107
rect 42510 -142350 42586 -141107
rect 43118 -142350 43194 -141107
rect 43726 -142350 43802 -141107
rect 44334 -142350 44410 -141107
rect 44942 -142350 45018 -141107
rect 45550 -142350 45626 -141107
rect 46158 -142350 46234 -141107
rect 46766 -142350 46842 -141107
rect 47374 -142350 47450 -141107
rect 47982 -142350 48058 -141107
rect 48590 -142350 48666 -141107
rect 49198 -142350 49274 -141107
rect 49806 -142350 49882 -141107
rect 50414 -142350 50490 -141107
rect 51022 -142350 51098 -141107
rect 51630 -142350 51706 -141107
rect 52238 -142350 52314 -141107
rect 52846 -142350 52922 -141107
rect 53454 -142350 53530 -141107
rect 54062 -142350 54138 -141107
rect 54670 -142350 54746 -141107
rect 55278 -142350 55354 -141107
rect 55886 -142350 55962 -141107
rect 56494 -142350 56570 -141107
rect 57102 -142350 57178 -141107
rect 57710 -142350 57786 -141107
rect 58318 -142350 58394 -141107
rect 58926 -142350 59002 -141107
rect 59534 -142350 59610 -141107
rect 60142 -142350 60218 -141107
rect 60750 -142350 60826 -141107
rect 61358 -142350 61434 -141107
rect 61966 -142350 62042 -141107
rect 62574 -142350 62650 -141107
rect 63182 -142350 63258 -141107
rect 63790 -142350 63866 -141107
rect 64398 -142350 64474 -141107
rect 65006 -142350 65082 -141107
rect 65614 -142350 65690 -141107
rect 66222 -142350 66298 -141107
rect 66830 -142350 66906 -141107
rect 67438 -142350 67514 -141107
rect 68046 -142350 68122 -141107
rect 68654 -142350 68730 -141107
rect 69262 -142350 69338 -141107
rect 69870 -142350 69946 -141107
rect 70478 -142350 70554 -141107
rect 71086 -142350 71162 -141107
rect 71694 -142350 71770 -141107
rect 72302 -142350 72378 -141107
rect 75744 -162352 75978 -141107
rect 76510 -142350 76586 -141107
rect 77118 -142350 77194 -141107
rect 77726 -142350 77802 -141107
rect 78334 -142350 78410 -141107
rect 78942 -142350 79018 -141107
rect 79550 -142350 79626 -141107
rect 80158 -142350 80234 -141107
rect 80766 -142350 80842 -141107
rect 81374 -142350 81450 -141107
rect 81982 -142350 82058 -141107
rect 82590 -142350 82666 -141107
rect 83198 -142350 83274 -141107
rect 83806 -142350 83882 -141107
rect 84414 -142350 84490 -141107
rect 85022 -142350 85098 -141107
rect 85630 -142350 85706 -141107
rect 86238 -142350 86314 -141107
rect 86846 -142350 86922 -141107
rect 87454 -142350 87530 -141107
rect 88062 -142350 88138 -141107
rect 88670 -142350 88746 -141107
rect 89278 -142350 89354 -141107
rect 89886 -142350 89962 -141107
rect 90494 -142350 90570 -141107
rect 91102 -142350 91178 -141107
rect 91710 -142350 91786 -141107
rect 92318 -142350 92394 -141107
rect 92926 -142350 93002 -141107
rect 93534 -142350 93610 -141107
rect 94142 -142350 94218 -141107
rect 94750 -142350 94826 -141107
rect 95358 -142350 95434 -141107
rect 95966 -142350 96042 -141107
rect 96574 -142350 96650 -141107
rect 97182 -142350 97258 -141107
rect 97790 -142350 97866 -141107
rect 98398 -142350 98474 -141107
rect 99006 -142350 99082 -141107
rect 99614 -142350 99690 -141107
rect 100222 -142350 100298 -141107
rect 100830 -142350 100906 -141107
rect 101438 -142350 101514 -141107
rect 102046 -142350 102122 -141107
rect 102654 -142350 102730 -141107
rect 103262 -142350 103338 -141107
rect 103870 -142350 103946 -141107
rect 104478 -142350 104554 -141107
rect 105086 -142350 105162 -141107
rect 105694 -142350 105770 -141107
rect 106302 -142350 106378 -141107
rect 109744 -162352 109978 -141107
rect 110510 -142350 110586 -141107
rect 111118 -142350 111194 -141107
rect 111726 -142350 111802 -141107
rect 112334 -142350 112410 -141107
rect 112942 -142350 113018 -141107
rect 113550 -142350 113626 -141107
rect 114158 -142350 114234 -141107
rect 114766 -142350 114842 -141107
rect 115374 -142350 115450 -141107
rect 115982 -142350 116058 -141107
rect 116590 -142350 116666 -141107
rect 117198 -142350 117274 -141107
rect 117806 -142350 117882 -141107
rect 118414 -142350 118490 -141107
rect 119022 -142350 119098 -141107
rect 119630 -142350 119706 -141107
rect 120238 -142350 120314 -141107
rect 120846 -142350 120922 -141107
rect 121454 -142350 121530 -141107
rect 122062 -142350 122138 -141107
rect 122670 -142350 122746 -141107
rect 123278 -142350 123354 -141107
rect 123886 -142350 123962 -141107
rect 124494 -142350 124570 -141107
rect 125102 -142350 125178 -141107
rect 125710 -142350 125786 -141107
rect 126318 -142350 126394 -141107
rect 126926 -142350 127002 -141107
rect 127534 -142350 127610 -141107
rect 128142 -142350 128218 -141107
rect 128750 -142350 128826 -141107
rect 129358 -142350 129434 -141107
rect 129966 -142350 130042 -141107
rect 130574 -142350 130650 -141107
rect 131182 -142350 131258 -141107
rect 131790 -142350 131866 -141107
rect 132398 -142350 132474 -141107
rect 133006 -142350 133082 -141107
rect 133614 -142350 133690 -141107
rect 134222 -142350 134298 -141107
rect 134830 -142350 134906 -141107
rect 135438 -142350 135514 -141107
rect 136046 -142350 136122 -141107
rect 136654 -142350 136730 -141107
rect 137262 -142350 137338 -141107
rect 137870 -142350 137946 -141107
rect 138478 -142350 138554 -141107
rect 139086 -142350 139162 -141107
rect 139694 -142350 139770 -141107
rect 140302 -142350 140378 -141107
rect 143744 -162352 143978 -141107
rect 144510 -142350 144586 -141107
rect 145118 -142350 145194 -141107
rect 145726 -142350 145802 -141107
rect 146334 -142350 146410 -141107
rect 146942 -142350 147018 -141107
rect 147550 -142350 147626 -141107
rect 148158 -142350 148234 -141107
rect 148766 -142350 148842 -141107
rect 149374 -142350 149450 -141107
rect 149982 -142350 150058 -141107
rect 150590 -142350 150666 -141107
rect 151198 -142350 151274 -141107
rect 151806 -142350 151882 -141107
rect 152414 -142350 152490 -141107
rect 153022 -142350 153098 -141107
rect 153630 -142350 153706 -141107
rect 154238 -142350 154314 -141107
rect 154846 -142350 154922 -141107
rect 155454 -142350 155530 -141107
rect 156062 -142350 156138 -141107
rect 156670 -142350 156746 -141107
rect 157278 -142350 157354 -141107
rect 157886 -142350 157962 -141107
rect 158494 -142350 158570 -141107
rect 159102 -142350 159178 -141107
rect 159710 -142350 159786 -141107
rect 160318 -142350 160394 -141107
rect 160926 -142350 161002 -141107
rect 161534 -142350 161610 -141107
rect 162142 -142350 162218 -141107
rect 162750 -142350 162826 -141107
rect 163358 -142350 163434 -141107
rect 163966 -142350 164042 -141107
rect 164574 -142350 164650 -141107
rect 165182 -142350 165258 -141107
rect 165790 -142350 165866 -141107
rect 166398 -142350 166474 -141107
rect 167006 -142350 167082 -141107
rect 167614 -142350 167690 -141107
rect 168222 -142350 168298 -141107
rect 168830 -142350 168906 -141107
rect 169438 -142350 169514 -141107
rect 170046 -142350 170122 -141107
rect 170654 -142350 170730 -141107
rect 171262 -142350 171338 -141107
rect 171870 -142350 171946 -141107
rect 172478 -142350 172554 -141107
rect 173086 -142350 173162 -141107
rect 173694 -142350 173770 -141107
rect 174302 -142350 174378 -141107
rect -97672 -164600 -72506 -163392
rect -59794 -163597 -59718 -162354
rect -59186 -163597 -59110 -162354
rect -58578 -163597 -58502 -162354
rect -57970 -163597 -57894 -162354
rect -57362 -163597 -57286 -162354
rect -56754 -163597 -56678 -162354
rect -56146 -163597 -56070 -162354
rect -55538 -163597 -55462 -162354
rect -54930 -163597 -54854 -162354
rect -54322 -163597 -54246 -162354
rect -53714 -163597 -53638 -162354
rect -53106 -163597 -53030 -162354
rect -52498 -163597 -52422 -162354
rect -51890 -163597 -51814 -162354
rect -51282 -163597 -51206 -162354
rect -50674 -163597 -50598 -162354
rect -50066 -163597 -49990 -162354
rect -49458 -163597 -49382 -162354
rect -48850 -163597 -48774 -162354
rect -48242 -163597 -48166 -162354
rect -47634 -163597 -47558 -162354
rect -47026 -163597 -46950 -162354
rect -46418 -163597 -46342 -162354
rect -45810 -163597 -45734 -162354
rect -45202 -163597 -45126 -162354
rect -44594 -163597 -44518 -162354
rect -43986 -163597 -43910 -162354
rect -43378 -163597 -43302 -162354
rect -42770 -163597 -42694 -162354
rect -42162 -163597 -42086 -162354
rect -41554 -163597 -41478 -162354
rect -40946 -163597 -40870 -162354
rect -40338 -163597 -40262 -162354
rect -39730 -163597 -39654 -162354
rect -39122 -163597 -39046 -162354
rect -38514 -163597 -38438 -162354
rect -37906 -163597 -37830 -162354
rect -37298 -163597 -37222 -162354
rect -36690 -163597 -36614 -162354
rect -36082 -163597 -36006 -162354
rect -35474 -163597 -35398 -162354
rect -34866 -163597 -34790 -162354
rect -34258 -163597 -34182 -162354
rect -33650 -163597 -33574 -162354
rect -33042 -163597 -32966 -162354
rect -32434 -163597 -32358 -162354
rect -31826 -163597 -31750 -162354
rect -31218 -163597 -31142 -162354
rect -30610 -163597 -30534 -162354
rect -30002 -163597 -29926 -162354
rect -25794 -163597 -25718 -162354
rect -25186 -163597 -25110 -162354
rect -24578 -163597 -24502 -162354
rect -23970 -163597 -23894 -162354
rect -23362 -163597 -23286 -162354
rect -22754 -163597 -22678 -162354
rect -22146 -163597 -22070 -162354
rect -21538 -163597 -21462 -162354
rect -20930 -163597 -20854 -162354
rect -20322 -163597 -20246 -162354
rect -19714 -163597 -19638 -162354
rect -19106 -163597 -19030 -162354
rect -18498 -163597 -18422 -162354
rect -17890 -163597 -17814 -162354
rect -17282 -163597 -17206 -162354
rect -16674 -163597 -16598 -162354
rect -16066 -163597 -15990 -162354
rect -15458 -163597 -15382 -162354
rect -14850 -163597 -14774 -162354
rect -14242 -163597 -14166 -162354
rect -13634 -163597 -13558 -162354
rect -13026 -163597 -12950 -162354
rect -12418 -163597 -12342 -162354
rect -11810 -163597 -11734 -162354
rect -11202 -163597 -11126 -162354
rect -10594 -163597 -10518 -162354
rect -9986 -163597 -9910 -162354
rect -9378 -163597 -9302 -162354
rect -8770 -163597 -8694 -162354
rect -8162 -163597 -8086 -162354
rect -7554 -163597 -7478 -162354
rect -6946 -163597 -6870 -162354
rect -6338 -163597 -6262 -162354
rect -5730 -163597 -5654 -162354
rect -5122 -163597 -5046 -162354
rect -4514 -163597 -4438 -162354
rect -3906 -163597 -3830 -162354
rect -3298 -163597 -3222 -162354
rect -2690 -163597 -2614 -162354
rect -2082 -163597 -2006 -162354
rect -1474 -163597 -1398 -162354
rect -866 -163597 -790 -162354
rect -258 -163597 -182 -162354
rect 350 -163597 426 -162354
rect 958 -163597 1034 -162354
rect 1566 -163597 1642 -162354
rect 2174 -163597 2250 -162354
rect 2782 -163597 2858 -162354
rect 3390 -163597 3466 -162354
rect 3998 -163597 4074 -162354
rect 8206 -163597 8282 -162354
rect 8814 -163597 8890 -162354
rect 9422 -163597 9498 -162354
rect 10030 -163597 10106 -162354
rect 10638 -163597 10714 -162354
rect 11246 -163597 11322 -162354
rect 11854 -163597 11930 -162354
rect 12462 -163597 12538 -162354
rect 13070 -163597 13146 -162354
rect 13678 -163597 13754 -162354
rect 14286 -163597 14362 -162354
rect 14894 -163597 14970 -162354
rect 15502 -163597 15578 -162354
rect 16110 -163597 16186 -162354
rect 16718 -163597 16794 -162354
rect 17326 -163597 17402 -162354
rect 17934 -163597 18010 -162354
rect 18542 -163597 18618 -162354
rect 19150 -163597 19226 -162354
rect 19758 -163597 19834 -162354
rect 20366 -163597 20442 -162354
rect 20974 -163597 21050 -162354
rect 21582 -163597 21658 -162354
rect 22190 -163597 22266 -162354
rect 22798 -163597 22874 -162354
rect 23406 -163597 23482 -162354
rect 24014 -163597 24090 -162354
rect 24622 -163597 24698 -162354
rect 25230 -163597 25306 -162354
rect 25838 -163597 25914 -162354
rect 26446 -163597 26522 -162354
rect 27054 -163597 27130 -162354
rect 27662 -163597 27738 -162354
rect 28270 -163597 28346 -162354
rect 28878 -163597 28954 -162354
rect 29486 -163597 29562 -162354
rect 30094 -163597 30170 -162354
rect 30702 -163597 30778 -162354
rect 31310 -163597 31386 -162354
rect 31918 -163597 31994 -162354
rect 32526 -163597 32602 -162354
rect 33134 -163597 33210 -162354
rect 33742 -163597 33818 -162354
rect 34350 -163597 34426 -162354
rect 34958 -163597 35034 -162354
rect 35566 -163597 35642 -162354
rect 36174 -163597 36250 -162354
rect 36782 -163597 36858 -162354
rect 37390 -163597 37466 -162354
rect 37998 -163597 38074 -162354
rect 42206 -163597 42282 -162354
rect 42814 -163597 42890 -162354
rect 43422 -163597 43498 -162354
rect 44030 -163597 44106 -162354
rect 44638 -163597 44714 -162354
rect 45246 -163597 45322 -162354
rect 45854 -163597 45930 -162354
rect 46462 -163597 46538 -162354
rect 47070 -163597 47146 -162354
rect 47678 -163597 47754 -162354
rect 48286 -163597 48362 -162354
rect 48894 -163597 48970 -162354
rect 49502 -163597 49578 -162354
rect 50110 -163597 50186 -162354
rect 50718 -163597 50794 -162354
rect 51326 -163597 51402 -162354
rect 51934 -163597 52010 -162354
rect 52542 -163597 52618 -162354
rect 53150 -163597 53226 -162354
rect 53758 -163597 53834 -162354
rect 54366 -163597 54442 -162354
rect 54974 -163597 55050 -162354
rect 55582 -163597 55658 -162354
rect 56190 -163597 56266 -162354
rect 56798 -163597 56874 -162354
rect 57406 -163597 57482 -162354
rect 58014 -163597 58090 -162354
rect 58622 -163597 58698 -162354
rect 59230 -163597 59306 -162354
rect 59838 -163597 59914 -162354
rect 60446 -163597 60522 -162354
rect 61054 -163597 61130 -162354
rect 61662 -163597 61738 -162354
rect 62270 -163597 62346 -162354
rect 62878 -163597 62954 -162354
rect 63486 -163597 63562 -162354
rect 64094 -163597 64170 -162354
rect 64702 -163597 64778 -162354
rect 65310 -163597 65386 -162354
rect 65918 -163597 65994 -162354
rect 66526 -163597 66602 -162354
rect 67134 -163597 67210 -162354
rect 67742 -163597 67818 -162354
rect 68350 -163597 68426 -162354
rect 68958 -163597 69034 -162354
rect 69566 -163597 69642 -162354
rect 70174 -163597 70250 -162354
rect 70782 -163597 70858 -162354
rect 71390 -163597 71466 -162354
rect 71998 -163597 72074 -162354
rect 76206 -163597 76282 -162354
rect 76814 -163597 76890 -162354
rect 77422 -163597 77498 -162354
rect 78030 -163597 78106 -162354
rect 78638 -163597 78714 -162354
rect 79246 -163597 79322 -162354
rect 79854 -163597 79930 -162354
rect 80462 -163597 80538 -162354
rect 81070 -163597 81146 -162354
rect 81678 -163597 81754 -162354
rect 82286 -163597 82362 -162354
rect 82894 -163597 82970 -162354
rect 83502 -163597 83578 -162354
rect 84110 -163597 84186 -162354
rect 84718 -163597 84794 -162354
rect 85326 -163597 85402 -162354
rect 85934 -163597 86010 -162354
rect 86542 -163597 86618 -162354
rect 87150 -163597 87226 -162354
rect 87758 -163597 87834 -162354
rect 88366 -163597 88442 -162354
rect 88974 -163597 89050 -162354
rect 89582 -163597 89658 -162354
rect 90190 -163597 90266 -162354
rect 90798 -163597 90874 -162354
rect 91406 -163597 91482 -162354
rect 92014 -163597 92090 -162354
rect 92622 -163597 92698 -162354
rect 93230 -163597 93306 -162354
rect 93838 -163597 93914 -162354
rect 94446 -163597 94522 -162354
rect 95054 -163597 95130 -162354
rect 95662 -163597 95738 -162354
rect 96270 -163597 96346 -162354
rect 96878 -163597 96954 -162354
rect 97486 -163597 97562 -162354
rect 98094 -163597 98170 -162354
rect 98702 -163597 98778 -162354
rect 99310 -163597 99386 -162354
rect 99918 -163597 99994 -162354
rect 100526 -163597 100602 -162354
rect 101134 -163597 101210 -162354
rect 101742 -163597 101818 -162354
rect 102350 -163597 102426 -162354
rect 102958 -163597 103034 -162354
rect 103566 -163597 103642 -162354
rect 104174 -163597 104250 -162354
rect 104782 -163597 104858 -162354
rect 105390 -163597 105466 -162354
rect 105998 -163597 106074 -162354
rect 110206 -163597 110282 -162354
rect 110814 -163597 110890 -162354
rect 111422 -163597 111498 -162354
rect 112030 -163597 112106 -162354
rect 112638 -163597 112714 -162354
rect 113246 -163597 113322 -162354
rect 113854 -163597 113930 -162354
rect 114462 -163597 114538 -162354
rect 115070 -163597 115146 -162354
rect 115678 -163597 115754 -162354
rect 116286 -163597 116362 -162354
rect 116894 -163597 116970 -162354
rect 117502 -163597 117578 -162354
rect 118110 -163597 118186 -162354
rect 118718 -163597 118794 -162354
rect 119326 -163597 119402 -162354
rect 119934 -163597 120010 -162354
rect 120542 -163597 120618 -162354
rect 121150 -163597 121226 -162354
rect 121758 -163597 121834 -162354
rect 122366 -163597 122442 -162354
rect 122974 -163597 123050 -162354
rect 123582 -163597 123658 -162354
rect 124190 -163597 124266 -162354
rect 124798 -163597 124874 -162354
rect 125406 -163597 125482 -162354
rect 126014 -163597 126090 -162354
rect 126622 -163597 126698 -162354
rect 127230 -163597 127306 -162354
rect 127838 -163597 127914 -162354
rect 128446 -163597 128522 -162354
rect 129054 -163597 129130 -162354
rect 129662 -163597 129738 -162354
rect 130270 -163597 130346 -162354
rect 130878 -163597 130954 -162354
rect 131486 -163597 131562 -162354
rect 132094 -163597 132170 -162354
rect 132702 -163597 132778 -162354
rect 133310 -163597 133386 -162354
rect 133918 -163597 133994 -162354
rect 134526 -163597 134602 -162354
rect 135134 -163597 135210 -162354
rect 135742 -163597 135818 -162354
rect 136350 -163597 136426 -162354
rect 136958 -163597 137034 -162354
rect 137566 -163597 137642 -162354
rect 138174 -163597 138250 -162354
rect 138782 -163597 138858 -162354
rect 139390 -163597 139466 -162354
rect 139998 -163597 140074 -162354
rect 144206 -163597 144282 -162354
rect 144814 -163597 144890 -162354
rect 145422 -163597 145498 -162354
rect 146030 -163597 146106 -162354
rect 146638 -163597 146714 -162354
rect 147246 -163597 147322 -162354
rect 147854 -163597 147930 -162354
rect 148462 -163597 148538 -162354
rect 149070 -163597 149146 -162354
rect 149678 -163597 149754 -162354
rect 150286 -163597 150362 -162354
rect 150894 -163597 150970 -162354
rect 151502 -163597 151578 -162354
rect 152110 -163597 152186 -162354
rect 152718 -163597 152794 -162354
rect 153326 -163597 153402 -162354
rect 153934 -163597 154010 -162354
rect 154542 -163597 154618 -162354
rect 155150 -163597 155226 -162354
rect 155758 -163597 155834 -162354
rect 156366 -163597 156442 -162354
rect 156974 -163597 157050 -162354
rect 157582 -163597 157658 -162354
rect 158190 -163597 158266 -162354
rect 158798 -163597 158874 -162354
rect 159406 -163597 159482 -162354
rect 160014 -163597 160090 -162354
rect 160622 -163597 160698 -162354
rect 161230 -163597 161306 -162354
rect 161838 -163597 161914 -162354
rect 162446 -163597 162522 -162354
rect 163054 -163597 163130 -162354
rect 163662 -163597 163738 -162354
rect 164270 -163597 164346 -162354
rect 164878 -163597 164954 -162354
rect 165486 -163597 165562 -162354
rect 166094 -163597 166170 -162354
rect 166702 -163597 166778 -162354
rect 167310 -163597 167386 -162354
rect 167918 -163597 167994 -162354
rect 168526 -163597 168602 -162354
rect 169134 -163597 169210 -162354
rect 169742 -163597 169818 -162354
rect 170350 -163597 170426 -162354
rect 170958 -163597 171034 -162354
rect 171566 -163597 171642 -162354
rect 172174 -163597 172250 -162354
rect 172782 -163597 172858 -162354
rect 173390 -163597 173466 -162354
rect 173998 -163597 174074 -162354
rect -59794 -165615 174682 -163597
rect -59794 -165659 145268 -165615
rect 145312 -165659 145368 -165615
rect 145412 -165659 145468 -165615
rect 145512 -165659 145568 -165615
rect 145612 -165659 145668 -165615
rect 145712 -165659 145768 -165615
rect 145812 -165659 145868 -165615
rect 145912 -165659 145968 -165615
rect 146012 -165659 146068 -165615
rect 146112 -165659 146168 -165615
rect 146212 -165659 146268 -165615
rect 146312 -165659 146368 -165615
rect 146412 -165659 146468 -165615
rect 146512 -165659 146568 -165615
rect 146612 -165659 146668 -165615
rect 146712 -165659 146768 -165615
rect 146812 -165659 147268 -165615
rect 147312 -165659 147368 -165615
rect 147412 -165659 147468 -165615
rect 147512 -165659 147568 -165615
rect 147612 -165659 147668 -165615
rect 147712 -165659 147768 -165615
rect 147812 -165659 147868 -165615
rect 147912 -165659 147968 -165615
rect 148012 -165659 148068 -165615
rect 148112 -165659 148168 -165615
rect 148212 -165659 148268 -165615
rect 148312 -165659 148368 -165615
rect 148412 -165659 148468 -165615
rect 148512 -165659 148568 -165615
rect 148612 -165659 148668 -165615
rect 148712 -165659 148768 -165615
rect 148812 -165659 149268 -165615
rect 149312 -165659 149368 -165615
rect 149412 -165659 149468 -165615
rect 149512 -165659 149568 -165615
rect 149612 -165659 149668 -165615
rect 149712 -165659 149768 -165615
rect 149812 -165659 149868 -165615
rect 149912 -165659 149968 -165615
rect 150012 -165659 150068 -165615
rect 150112 -165659 150168 -165615
rect 150212 -165659 150268 -165615
rect 150312 -165659 150368 -165615
rect 150412 -165659 150468 -165615
rect 150512 -165659 150568 -165615
rect 150612 -165659 150668 -165615
rect 150712 -165659 150768 -165615
rect 150812 -165659 151268 -165615
rect 151312 -165659 151368 -165615
rect 151412 -165659 151468 -165615
rect 151512 -165659 151568 -165615
rect 151612 -165659 151668 -165615
rect 151712 -165659 151768 -165615
rect 151812 -165659 151868 -165615
rect 151912 -165659 151968 -165615
rect 152012 -165659 152068 -165615
rect 152112 -165659 152168 -165615
rect 152212 -165659 152268 -165615
rect 152312 -165659 152368 -165615
rect 152412 -165659 152468 -165615
rect 152512 -165659 152568 -165615
rect 152612 -165659 152668 -165615
rect 152712 -165659 152768 -165615
rect 152812 -165659 174682 -165615
rect -59794 -165715 174682 -165659
rect -59794 -165759 145268 -165715
rect 145312 -165759 145368 -165715
rect 145412 -165759 145468 -165715
rect 145512 -165759 145568 -165715
rect 145612 -165759 145668 -165715
rect 145712 -165759 145768 -165715
rect 145812 -165759 145868 -165715
rect 145912 -165759 145968 -165715
rect 146012 -165759 146068 -165715
rect 146112 -165759 146168 -165715
rect 146212 -165759 146268 -165715
rect 146312 -165759 146368 -165715
rect 146412 -165759 146468 -165715
rect 146512 -165759 146568 -165715
rect 146612 -165759 146668 -165715
rect 146712 -165759 146768 -165715
rect 146812 -165759 147268 -165715
rect 147312 -165759 147368 -165715
rect 147412 -165759 147468 -165715
rect 147512 -165759 147568 -165715
rect 147612 -165759 147668 -165715
rect 147712 -165759 147768 -165715
rect 147812 -165759 147868 -165715
rect 147912 -165759 147968 -165715
rect 148012 -165759 148068 -165715
rect 148112 -165759 148168 -165715
rect 148212 -165759 148268 -165715
rect 148312 -165759 148368 -165715
rect 148412 -165759 148468 -165715
rect 148512 -165759 148568 -165715
rect 148612 -165759 148668 -165715
rect 148712 -165759 148768 -165715
rect 148812 -165759 149268 -165715
rect 149312 -165759 149368 -165715
rect 149412 -165759 149468 -165715
rect 149512 -165759 149568 -165715
rect 149612 -165759 149668 -165715
rect 149712 -165759 149768 -165715
rect 149812 -165759 149868 -165715
rect 149912 -165759 149968 -165715
rect 150012 -165759 150068 -165715
rect 150112 -165759 150168 -165715
rect 150212 -165759 150268 -165715
rect 150312 -165759 150368 -165715
rect 150412 -165759 150468 -165715
rect 150512 -165759 150568 -165715
rect 150612 -165759 150668 -165715
rect 150712 -165759 150768 -165715
rect 150812 -165759 151268 -165715
rect 151312 -165759 151368 -165715
rect 151412 -165759 151468 -165715
rect 151512 -165759 151568 -165715
rect 151612 -165759 151668 -165715
rect 151712 -165759 151768 -165715
rect 151812 -165759 151868 -165715
rect 151912 -165759 151968 -165715
rect 152012 -165759 152068 -165715
rect 152112 -165759 152168 -165715
rect 152212 -165759 152268 -165715
rect 152312 -165759 152368 -165715
rect 152412 -165759 152468 -165715
rect 152512 -165759 152568 -165715
rect 152612 -165759 152668 -165715
rect 152712 -165759 152768 -165715
rect 152812 -165759 174682 -165715
rect -59794 -165815 174682 -165759
rect -59794 -165859 145268 -165815
rect 145312 -165859 145368 -165815
rect 145412 -165859 145468 -165815
rect 145512 -165859 145568 -165815
rect 145612 -165859 145668 -165815
rect 145712 -165859 145768 -165815
rect 145812 -165859 145868 -165815
rect 145912 -165859 145968 -165815
rect 146012 -165859 146068 -165815
rect 146112 -165859 146168 -165815
rect 146212 -165859 146268 -165815
rect 146312 -165859 146368 -165815
rect 146412 -165859 146468 -165815
rect 146512 -165859 146568 -165815
rect 146612 -165859 146668 -165815
rect 146712 -165859 146768 -165815
rect 146812 -165859 147268 -165815
rect 147312 -165859 147368 -165815
rect 147412 -165859 147468 -165815
rect 147512 -165859 147568 -165815
rect 147612 -165859 147668 -165815
rect 147712 -165859 147768 -165815
rect 147812 -165859 147868 -165815
rect 147912 -165859 147968 -165815
rect 148012 -165859 148068 -165815
rect 148112 -165859 148168 -165815
rect 148212 -165859 148268 -165815
rect 148312 -165859 148368 -165815
rect 148412 -165859 148468 -165815
rect 148512 -165859 148568 -165815
rect 148612 -165859 148668 -165815
rect 148712 -165859 148768 -165815
rect 148812 -165859 149268 -165815
rect 149312 -165859 149368 -165815
rect 149412 -165859 149468 -165815
rect 149512 -165859 149568 -165815
rect 149612 -165859 149668 -165815
rect 149712 -165859 149768 -165815
rect 149812 -165859 149868 -165815
rect 149912 -165859 149968 -165815
rect 150012 -165859 150068 -165815
rect 150112 -165859 150168 -165815
rect 150212 -165859 150268 -165815
rect 150312 -165859 150368 -165815
rect 150412 -165859 150468 -165815
rect 150512 -165859 150568 -165815
rect 150612 -165859 150668 -165815
rect 150712 -165859 150768 -165815
rect 150812 -165859 151268 -165815
rect 151312 -165859 151368 -165815
rect 151412 -165859 151468 -165815
rect 151512 -165859 151568 -165815
rect 151612 -165859 151668 -165815
rect 151712 -165859 151768 -165815
rect 151812 -165859 151868 -165815
rect 151912 -165859 151968 -165815
rect 152012 -165859 152068 -165815
rect 152112 -165859 152168 -165815
rect 152212 -165859 152268 -165815
rect 152312 -165859 152368 -165815
rect 152412 -165859 152468 -165815
rect 152512 -165859 152568 -165815
rect 152612 -165859 152668 -165815
rect 152712 -165859 152768 -165815
rect 152812 -165859 174682 -165815
rect -59794 -165915 174682 -165859
rect -59794 -165959 145268 -165915
rect 145312 -165959 145368 -165915
rect 145412 -165959 145468 -165915
rect 145512 -165959 145568 -165915
rect 145612 -165959 145668 -165915
rect 145712 -165959 145768 -165915
rect 145812 -165959 145868 -165915
rect 145912 -165959 145968 -165915
rect 146012 -165959 146068 -165915
rect 146112 -165959 146168 -165915
rect 146212 -165959 146268 -165915
rect 146312 -165959 146368 -165915
rect 146412 -165959 146468 -165915
rect 146512 -165959 146568 -165915
rect 146612 -165959 146668 -165915
rect 146712 -165959 146768 -165915
rect 146812 -165959 147268 -165915
rect 147312 -165959 147368 -165915
rect 147412 -165959 147468 -165915
rect 147512 -165959 147568 -165915
rect 147612 -165959 147668 -165915
rect 147712 -165959 147768 -165915
rect 147812 -165959 147868 -165915
rect 147912 -165959 147968 -165915
rect 148012 -165959 148068 -165915
rect 148112 -165959 148168 -165915
rect 148212 -165959 148268 -165915
rect 148312 -165959 148368 -165915
rect 148412 -165959 148468 -165915
rect 148512 -165959 148568 -165915
rect 148612 -165959 148668 -165915
rect 148712 -165959 148768 -165915
rect 148812 -165959 149268 -165915
rect 149312 -165959 149368 -165915
rect 149412 -165959 149468 -165915
rect 149512 -165959 149568 -165915
rect 149612 -165959 149668 -165915
rect 149712 -165959 149768 -165915
rect 149812 -165959 149868 -165915
rect 149912 -165959 149968 -165915
rect 150012 -165959 150068 -165915
rect 150112 -165959 150168 -165915
rect 150212 -165959 150268 -165915
rect 150312 -165959 150368 -165915
rect 150412 -165959 150468 -165915
rect 150512 -165959 150568 -165915
rect 150612 -165959 150668 -165915
rect 150712 -165959 150768 -165915
rect 150812 -165959 151268 -165915
rect 151312 -165959 151368 -165915
rect 151412 -165959 151468 -165915
rect 151512 -165959 151568 -165915
rect 151612 -165959 151668 -165915
rect 151712 -165959 151768 -165915
rect 151812 -165959 151868 -165915
rect 151912 -165959 151968 -165915
rect 152012 -165959 152068 -165915
rect 152112 -165959 152168 -165915
rect 152212 -165959 152268 -165915
rect 152312 -165959 152368 -165915
rect 152412 -165959 152468 -165915
rect 152512 -165959 152568 -165915
rect 152612 -165959 152668 -165915
rect 152712 -165959 152768 -165915
rect 152812 -165959 174682 -165915
rect -59794 -166015 174682 -165959
rect -59794 -166059 145268 -166015
rect 145312 -166059 145368 -166015
rect 145412 -166059 145468 -166015
rect 145512 -166059 145568 -166015
rect 145612 -166059 145668 -166015
rect 145712 -166059 145768 -166015
rect 145812 -166059 145868 -166015
rect 145912 -166059 145968 -166015
rect 146012 -166059 146068 -166015
rect 146112 -166059 146168 -166015
rect 146212 -166059 146268 -166015
rect 146312 -166059 146368 -166015
rect 146412 -166059 146468 -166015
rect 146512 -166059 146568 -166015
rect 146612 -166059 146668 -166015
rect 146712 -166059 146768 -166015
rect 146812 -166059 147268 -166015
rect 147312 -166059 147368 -166015
rect 147412 -166059 147468 -166015
rect 147512 -166059 147568 -166015
rect 147612 -166059 147668 -166015
rect 147712 -166059 147768 -166015
rect 147812 -166059 147868 -166015
rect 147912 -166059 147968 -166015
rect 148012 -166059 148068 -166015
rect 148112 -166059 148168 -166015
rect 148212 -166059 148268 -166015
rect 148312 -166059 148368 -166015
rect 148412 -166059 148468 -166015
rect 148512 -166059 148568 -166015
rect 148612 -166059 148668 -166015
rect 148712 -166059 148768 -166015
rect 148812 -166059 149268 -166015
rect 149312 -166059 149368 -166015
rect 149412 -166059 149468 -166015
rect 149512 -166059 149568 -166015
rect 149612 -166059 149668 -166015
rect 149712 -166059 149768 -166015
rect 149812 -166059 149868 -166015
rect 149912 -166059 149968 -166015
rect 150012 -166059 150068 -166015
rect 150112 -166059 150168 -166015
rect 150212 -166059 150268 -166015
rect 150312 -166059 150368 -166015
rect 150412 -166059 150468 -166015
rect 150512 -166059 150568 -166015
rect 150612 -166059 150668 -166015
rect 150712 -166059 150768 -166015
rect 150812 -166059 151268 -166015
rect 151312 -166059 151368 -166015
rect 151412 -166059 151468 -166015
rect 151512 -166059 151568 -166015
rect 151612 -166059 151668 -166015
rect 151712 -166059 151768 -166015
rect 151812 -166059 151868 -166015
rect 151912 -166059 151968 -166015
rect 152012 -166059 152068 -166015
rect 152112 -166059 152168 -166015
rect 152212 -166059 152268 -166015
rect 152312 -166059 152368 -166015
rect 152412 -166059 152468 -166015
rect 152512 -166059 152568 -166015
rect 152612 -166059 152668 -166015
rect 152712 -166059 152768 -166015
rect 152812 -166059 174682 -166015
rect -59794 -166115 174682 -166059
rect -59794 -166159 145268 -166115
rect 145312 -166159 145368 -166115
rect 145412 -166159 145468 -166115
rect 145512 -166159 145568 -166115
rect 145612 -166159 145668 -166115
rect 145712 -166159 145768 -166115
rect 145812 -166159 145868 -166115
rect 145912 -166159 145968 -166115
rect 146012 -166159 146068 -166115
rect 146112 -166159 146168 -166115
rect 146212 -166159 146268 -166115
rect 146312 -166159 146368 -166115
rect 146412 -166159 146468 -166115
rect 146512 -166159 146568 -166115
rect 146612 -166159 146668 -166115
rect 146712 -166159 146768 -166115
rect 146812 -166159 147268 -166115
rect 147312 -166159 147368 -166115
rect 147412 -166159 147468 -166115
rect 147512 -166159 147568 -166115
rect 147612 -166159 147668 -166115
rect 147712 -166159 147768 -166115
rect 147812 -166159 147868 -166115
rect 147912 -166159 147968 -166115
rect 148012 -166159 148068 -166115
rect 148112 -166159 148168 -166115
rect 148212 -166159 148268 -166115
rect 148312 -166159 148368 -166115
rect 148412 -166159 148468 -166115
rect 148512 -166159 148568 -166115
rect 148612 -166159 148668 -166115
rect 148712 -166159 148768 -166115
rect 148812 -166159 149268 -166115
rect 149312 -166159 149368 -166115
rect 149412 -166159 149468 -166115
rect 149512 -166159 149568 -166115
rect 149612 -166159 149668 -166115
rect 149712 -166159 149768 -166115
rect 149812 -166159 149868 -166115
rect 149912 -166159 149968 -166115
rect 150012 -166159 150068 -166115
rect 150112 -166159 150168 -166115
rect 150212 -166159 150268 -166115
rect 150312 -166159 150368 -166115
rect 150412 -166159 150468 -166115
rect 150512 -166159 150568 -166115
rect 150612 -166159 150668 -166115
rect 150712 -166159 150768 -166115
rect 150812 -166159 151268 -166115
rect 151312 -166159 151368 -166115
rect 151412 -166159 151468 -166115
rect 151512 -166159 151568 -166115
rect 151612 -166159 151668 -166115
rect 151712 -166159 151768 -166115
rect 151812 -166159 151868 -166115
rect 151912 -166159 151968 -166115
rect 152012 -166159 152068 -166115
rect 152112 -166159 152168 -166115
rect 152212 -166159 152268 -166115
rect 152312 -166159 152368 -166115
rect 152412 -166159 152468 -166115
rect 152512 -166159 152568 -166115
rect 152612 -166159 152668 -166115
rect 152712 -166159 152768 -166115
rect 152812 -166159 174682 -166115
rect -59794 -166215 174682 -166159
rect -59794 -166259 145268 -166215
rect 145312 -166259 145368 -166215
rect 145412 -166259 145468 -166215
rect 145512 -166259 145568 -166215
rect 145612 -166259 145668 -166215
rect 145712 -166259 145768 -166215
rect 145812 -166259 145868 -166215
rect 145912 -166259 145968 -166215
rect 146012 -166259 146068 -166215
rect 146112 -166259 146168 -166215
rect 146212 -166259 146268 -166215
rect 146312 -166259 146368 -166215
rect 146412 -166259 146468 -166215
rect 146512 -166259 146568 -166215
rect 146612 -166259 146668 -166215
rect 146712 -166259 146768 -166215
rect 146812 -166259 147268 -166215
rect 147312 -166259 147368 -166215
rect 147412 -166259 147468 -166215
rect 147512 -166259 147568 -166215
rect 147612 -166259 147668 -166215
rect 147712 -166259 147768 -166215
rect 147812 -166259 147868 -166215
rect 147912 -166259 147968 -166215
rect 148012 -166259 148068 -166215
rect 148112 -166259 148168 -166215
rect 148212 -166259 148268 -166215
rect 148312 -166259 148368 -166215
rect 148412 -166259 148468 -166215
rect 148512 -166259 148568 -166215
rect 148612 -166259 148668 -166215
rect 148712 -166259 148768 -166215
rect 148812 -166259 149268 -166215
rect 149312 -166259 149368 -166215
rect 149412 -166259 149468 -166215
rect 149512 -166259 149568 -166215
rect 149612 -166259 149668 -166215
rect 149712 -166259 149768 -166215
rect 149812 -166259 149868 -166215
rect 149912 -166259 149968 -166215
rect 150012 -166259 150068 -166215
rect 150112 -166259 150168 -166215
rect 150212 -166259 150268 -166215
rect 150312 -166259 150368 -166215
rect 150412 -166259 150468 -166215
rect 150512 -166259 150568 -166215
rect 150612 -166259 150668 -166215
rect 150712 -166259 150768 -166215
rect 150812 -166259 151268 -166215
rect 151312 -166259 151368 -166215
rect 151412 -166259 151468 -166215
rect 151512 -166259 151568 -166215
rect 151612 -166259 151668 -166215
rect 151712 -166259 151768 -166215
rect 151812 -166259 151868 -166215
rect 151912 -166259 151968 -166215
rect 152012 -166259 152068 -166215
rect 152112 -166259 152168 -166215
rect 152212 -166259 152268 -166215
rect 152312 -166259 152368 -166215
rect 152412 -166259 152468 -166215
rect 152512 -166259 152568 -166215
rect 152612 -166259 152668 -166215
rect 152712 -166259 152768 -166215
rect 152812 -166259 174682 -166215
rect -59794 -166315 174682 -166259
rect -59794 -166359 145268 -166315
rect 145312 -166359 145368 -166315
rect 145412 -166359 145468 -166315
rect 145512 -166359 145568 -166315
rect 145612 -166359 145668 -166315
rect 145712 -166359 145768 -166315
rect 145812 -166359 145868 -166315
rect 145912 -166359 145968 -166315
rect 146012 -166359 146068 -166315
rect 146112 -166359 146168 -166315
rect 146212 -166359 146268 -166315
rect 146312 -166359 146368 -166315
rect 146412 -166359 146468 -166315
rect 146512 -166359 146568 -166315
rect 146612 -166359 146668 -166315
rect 146712 -166359 146768 -166315
rect 146812 -166359 147268 -166315
rect 147312 -166359 147368 -166315
rect 147412 -166359 147468 -166315
rect 147512 -166359 147568 -166315
rect 147612 -166359 147668 -166315
rect 147712 -166359 147768 -166315
rect 147812 -166359 147868 -166315
rect 147912 -166359 147968 -166315
rect 148012 -166359 148068 -166315
rect 148112 -166359 148168 -166315
rect 148212 -166359 148268 -166315
rect 148312 -166359 148368 -166315
rect 148412 -166359 148468 -166315
rect 148512 -166359 148568 -166315
rect 148612 -166359 148668 -166315
rect 148712 -166359 148768 -166315
rect 148812 -166359 149268 -166315
rect 149312 -166359 149368 -166315
rect 149412 -166359 149468 -166315
rect 149512 -166359 149568 -166315
rect 149612 -166359 149668 -166315
rect 149712 -166359 149768 -166315
rect 149812 -166359 149868 -166315
rect 149912 -166359 149968 -166315
rect 150012 -166359 150068 -166315
rect 150112 -166359 150168 -166315
rect 150212 -166359 150268 -166315
rect 150312 -166359 150368 -166315
rect 150412 -166359 150468 -166315
rect 150512 -166359 150568 -166315
rect 150612 -166359 150668 -166315
rect 150712 -166359 150768 -166315
rect 150812 -166359 151268 -166315
rect 151312 -166359 151368 -166315
rect 151412 -166359 151468 -166315
rect 151512 -166359 151568 -166315
rect 151612 -166359 151668 -166315
rect 151712 -166359 151768 -166315
rect 151812 -166359 151868 -166315
rect 151912 -166359 151968 -166315
rect 152012 -166359 152068 -166315
rect 152112 -166359 152168 -166315
rect 152212 -166359 152268 -166315
rect 152312 -166359 152368 -166315
rect 152412 -166359 152468 -166315
rect 152512 -166359 152568 -166315
rect 152612 -166359 152668 -166315
rect 152712 -166359 152768 -166315
rect 152812 -166359 174682 -166315
rect -59794 -166415 174682 -166359
rect -59794 -166459 145268 -166415
rect 145312 -166459 145368 -166415
rect 145412 -166459 145468 -166415
rect 145512 -166459 145568 -166415
rect 145612 -166459 145668 -166415
rect 145712 -166459 145768 -166415
rect 145812 -166459 145868 -166415
rect 145912 -166459 145968 -166415
rect 146012 -166459 146068 -166415
rect 146112 -166459 146168 -166415
rect 146212 -166459 146268 -166415
rect 146312 -166459 146368 -166415
rect 146412 -166459 146468 -166415
rect 146512 -166459 146568 -166415
rect 146612 -166459 146668 -166415
rect 146712 -166459 146768 -166415
rect 146812 -166459 147268 -166415
rect 147312 -166459 147368 -166415
rect 147412 -166459 147468 -166415
rect 147512 -166459 147568 -166415
rect 147612 -166459 147668 -166415
rect 147712 -166459 147768 -166415
rect 147812 -166459 147868 -166415
rect 147912 -166459 147968 -166415
rect 148012 -166459 148068 -166415
rect 148112 -166459 148168 -166415
rect 148212 -166459 148268 -166415
rect 148312 -166459 148368 -166415
rect 148412 -166459 148468 -166415
rect 148512 -166459 148568 -166415
rect 148612 -166459 148668 -166415
rect 148712 -166459 148768 -166415
rect 148812 -166459 149268 -166415
rect 149312 -166459 149368 -166415
rect 149412 -166459 149468 -166415
rect 149512 -166459 149568 -166415
rect 149612 -166459 149668 -166415
rect 149712 -166459 149768 -166415
rect 149812 -166459 149868 -166415
rect 149912 -166459 149968 -166415
rect 150012 -166459 150068 -166415
rect 150112 -166459 150168 -166415
rect 150212 -166459 150268 -166415
rect 150312 -166459 150368 -166415
rect 150412 -166459 150468 -166415
rect 150512 -166459 150568 -166415
rect 150612 -166459 150668 -166415
rect 150712 -166459 150768 -166415
rect 150812 -166459 151268 -166415
rect 151312 -166459 151368 -166415
rect 151412 -166459 151468 -166415
rect 151512 -166459 151568 -166415
rect 151612 -166459 151668 -166415
rect 151712 -166459 151768 -166415
rect 151812 -166459 151868 -166415
rect 151912 -166459 151968 -166415
rect 152012 -166459 152068 -166415
rect 152112 -166459 152168 -166415
rect 152212 -166459 152268 -166415
rect 152312 -166459 152368 -166415
rect 152412 -166459 152468 -166415
rect 152512 -166459 152568 -166415
rect 152612 -166459 152668 -166415
rect 152712 -166459 152768 -166415
rect 152812 -166459 174682 -166415
rect -59794 -166515 174682 -166459
rect -59794 -166559 145268 -166515
rect 145312 -166559 145368 -166515
rect 145412 -166559 145468 -166515
rect 145512 -166559 145568 -166515
rect 145612 -166559 145668 -166515
rect 145712 -166559 145768 -166515
rect 145812 -166559 145868 -166515
rect 145912 -166559 145968 -166515
rect 146012 -166559 146068 -166515
rect 146112 -166559 146168 -166515
rect 146212 -166559 146268 -166515
rect 146312 -166559 146368 -166515
rect 146412 -166559 146468 -166515
rect 146512 -166559 146568 -166515
rect 146612 -166559 146668 -166515
rect 146712 -166559 146768 -166515
rect 146812 -166559 147268 -166515
rect 147312 -166559 147368 -166515
rect 147412 -166559 147468 -166515
rect 147512 -166559 147568 -166515
rect 147612 -166559 147668 -166515
rect 147712 -166559 147768 -166515
rect 147812 -166559 147868 -166515
rect 147912 -166559 147968 -166515
rect 148012 -166559 148068 -166515
rect 148112 -166559 148168 -166515
rect 148212 -166559 148268 -166515
rect 148312 -166559 148368 -166515
rect 148412 -166559 148468 -166515
rect 148512 -166559 148568 -166515
rect 148612 -166559 148668 -166515
rect 148712 -166559 148768 -166515
rect 148812 -166559 149268 -166515
rect 149312 -166559 149368 -166515
rect 149412 -166559 149468 -166515
rect 149512 -166559 149568 -166515
rect 149612 -166559 149668 -166515
rect 149712 -166559 149768 -166515
rect 149812 -166559 149868 -166515
rect 149912 -166559 149968 -166515
rect 150012 -166559 150068 -166515
rect 150112 -166559 150168 -166515
rect 150212 -166559 150268 -166515
rect 150312 -166559 150368 -166515
rect 150412 -166559 150468 -166515
rect 150512 -166559 150568 -166515
rect 150612 -166559 150668 -166515
rect 150712 -166559 150768 -166515
rect 150812 -166559 151268 -166515
rect 151312 -166559 151368 -166515
rect 151412 -166559 151468 -166515
rect 151512 -166559 151568 -166515
rect 151612 -166559 151668 -166515
rect 151712 -166559 151768 -166515
rect 151812 -166559 151868 -166515
rect 151912 -166559 151968 -166515
rect 152012 -166559 152068 -166515
rect 152112 -166559 152168 -166515
rect 152212 -166559 152268 -166515
rect 152312 -166559 152368 -166515
rect 152412 -166559 152468 -166515
rect 152512 -166559 152568 -166515
rect 152612 -166559 152668 -166515
rect 152712 -166559 152768 -166515
rect 152812 -166559 174682 -166515
rect -59794 -166615 174682 -166559
rect -59794 -166659 145268 -166615
rect 145312 -166659 145368 -166615
rect 145412 -166659 145468 -166615
rect 145512 -166659 145568 -166615
rect 145612 -166659 145668 -166615
rect 145712 -166659 145768 -166615
rect 145812 -166659 145868 -166615
rect 145912 -166659 145968 -166615
rect 146012 -166659 146068 -166615
rect 146112 -166659 146168 -166615
rect 146212 -166659 146268 -166615
rect 146312 -166659 146368 -166615
rect 146412 -166659 146468 -166615
rect 146512 -166659 146568 -166615
rect 146612 -166659 146668 -166615
rect 146712 -166659 146768 -166615
rect 146812 -166659 147268 -166615
rect 147312 -166659 147368 -166615
rect 147412 -166659 147468 -166615
rect 147512 -166659 147568 -166615
rect 147612 -166659 147668 -166615
rect 147712 -166659 147768 -166615
rect 147812 -166659 147868 -166615
rect 147912 -166659 147968 -166615
rect 148012 -166659 148068 -166615
rect 148112 -166659 148168 -166615
rect 148212 -166659 148268 -166615
rect 148312 -166659 148368 -166615
rect 148412 -166659 148468 -166615
rect 148512 -166659 148568 -166615
rect 148612 -166659 148668 -166615
rect 148712 -166659 148768 -166615
rect 148812 -166659 149268 -166615
rect 149312 -166659 149368 -166615
rect 149412 -166659 149468 -166615
rect 149512 -166659 149568 -166615
rect 149612 -166659 149668 -166615
rect 149712 -166659 149768 -166615
rect 149812 -166659 149868 -166615
rect 149912 -166659 149968 -166615
rect 150012 -166659 150068 -166615
rect 150112 -166659 150168 -166615
rect 150212 -166659 150268 -166615
rect 150312 -166659 150368 -166615
rect 150412 -166659 150468 -166615
rect 150512 -166659 150568 -166615
rect 150612 -166659 150668 -166615
rect 150712 -166659 150768 -166615
rect 150812 -166659 151268 -166615
rect 151312 -166659 151368 -166615
rect 151412 -166659 151468 -166615
rect 151512 -166659 151568 -166615
rect 151612 -166659 151668 -166615
rect 151712 -166659 151768 -166615
rect 151812 -166659 151868 -166615
rect 151912 -166659 151968 -166615
rect 152012 -166659 152068 -166615
rect 152112 -166659 152168 -166615
rect 152212 -166659 152268 -166615
rect 152312 -166659 152368 -166615
rect 152412 -166659 152468 -166615
rect 152512 -166659 152568 -166615
rect 152612 -166659 152668 -166615
rect 152712 -166659 152768 -166615
rect 152812 -166659 174682 -166615
rect -59794 -166715 174682 -166659
rect -59794 -166759 145268 -166715
rect 145312 -166759 145368 -166715
rect 145412 -166759 145468 -166715
rect 145512 -166759 145568 -166715
rect 145612 -166759 145668 -166715
rect 145712 -166759 145768 -166715
rect 145812 -166759 145868 -166715
rect 145912 -166759 145968 -166715
rect 146012 -166759 146068 -166715
rect 146112 -166759 146168 -166715
rect 146212 -166759 146268 -166715
rect 146312 -166759 146368 -166715
rect 146412 -166759 146468 -166715
rect 146512 -166759 146568 -166715
rect 146612 -166759 146668 -166715
rect 146712 -166759 146768 -166715
rect 146812 -166759 147268 -166715
rect 147312 -166759 147368 -166715
rect 147412 -166759 147468 -166715
rect 147512 -166759 147568 -166715
rect 147612 -166759 147668 -166715
rect 147712 -166759 147768 -166715
rect 147812 -166759 147868 -166715
rect 147912 -166759 147968 -166715
rect 148012 -166759 148068 -166715
rect 148112 -166759 148168 -166715
rect 148212 -166759 148268 -166715
rect 148312 -166759 148368 -166715
rect 148412 -166759 148468 -166715
rect 148512 -166759 148568 -166715
rect 148612 -166759 148668 -166715
rect 148712 -166759 148768 -166715
rect 148812 -166759 149268 -166715
rect 149312 -166759 149368 -166715
rect 149412 -166759 149468 -166715
rect 149512 -166759 149568 -166715
rect 149612 -166759 149668 -166715
rect 149712 -166759 149768 -166715
rect 149812 -166759 149868 -166715
rect 149912 -166759 149968 -166715
rect 150012 -166759 150068 -166715
rect 150112 -166759 150168 -166715
rect 150212 -166759 150268 -166715
rect 150312 -166759 150368 -166715
rect 150412 -166759 150468 -166715
rect 150512 -166759 150568 -166715
rect 150612 -166759 150668 -166715
rect 150712 -166759 150768 -166715
rect 150812 -166759 151268 -166715
rect 151312 -166759 151368 -166715
rect 151412 -166759 151468 -166715
rect 151512 -166759 151568 -166715
rect 151612 -166759 151668 -166715
rect 151712 -166759 151768 -166715
rect 151812 -166759 151868 -166715
rect 151912 -166759 151968 -166715
rect 152012 -166759 152068 -166715
rect 152112 -166759 152168 -166715
rect 152212 -166759 152268 -166715
rect 152312 -166759 152368 -166715
rect 152412 -166759 152468 -166715
rect 152512 -166759 152568 -166715
rect 152612 -166759 152668 -166715
rect 152712 -166759 152768 -166715
rect 152812 -166759 174682 -166715
rect -59794 -166815 174682 -166759
rect -59794 -166859 145268 -166815
rect 145312 -166859 145368 -166815
rect 145412 -166859 145468 -166815
rect 145512 -166859 145568 -166815
rect 145612 -166859 145668 -166815
rect 145712 -166859 145768 -166815
rect 145812 -166859 145868 -166815
rect 145912 -166859 145968 -166815
rect 146012 -166859 146068 -166815
rect 146112 -166859 146168 -166815
rect 146212 -166859 146268 -166815
rect 146312 -166859 146368 -166815
rect 146412 -166859 146468 -166815
rect 146512 -166859 146568 -166815
rect 146612 -166859 146668 -166815
rect 146712 -166859 146768 -166815
rect 146812 -166859 147268 -166815
rect 147312 -166859 147368 -166815
rect 147412 -166859 147468 -166815
rect 147512 -166859 147568 -166815
rect 147612 -166859 147668 -166815
rect 147712 -166859 147768 -166815
rect 147812 -166859 147868 -166815
rect 147912 -166859 147968 -166815
rect 148012 -166859 148068 -166815
rect 148112 -166859 148168 -166815
rect 148212 -166859 148268 -166815
rect 148312 -166859 148368 -166815
rect 148412 -166859 148468 -166815
rect 148512 -166859 148568 -166815
rect 148612 -166859 148668 -166815
rect 148712 -166859 148768 -166815
rect 148812 -166859 149268 -166815
rect 149312 -166859 149368 -166815
rect 149412 -166859 149468 -166815
rect 149512 -166859 149568 -166815
rect 149612 -166859 149668 -166815
rect 149712 -166859 149768 -166815
rect 149812 -166859 149868 -166815
rect 149912 -166859 149968 -166815
rect 150012 -166859 150068 -166815
rect 150112 -166859 150168 -166815
rect 150212 -166859 150268 -166815
rect 150312 -166859 150368 -166815
rect 150412 -166859 150468 -166815
rect 150512 -166859 150568 -166815
rect 150612 -166859 150668 -166815
rect 150712 -166859 150768 -166815
rect 150812 -166859 151268 -166815
rect 151312 -166859 151368 -166815
rect 151412 -166859 151468 -166815
rect 151512 -166859 151568 -166815
rect 151612 -166859 151668 -166815
rect 151712 -166859 151768 -166815
rect 151812 -166859 151868 -166815
rect 151912 -166859 151968 -166815
rect 152012 -166859 152068 -166815
rect 152112 -166859 152168 -166815
rect 152212 -166859 152268 -166815
rect 152312 -166859 152368 -166815
rect 152412 -166859 152468 -166815
rect 152512 -166859 152568 -166815
rect 152612 -166859 152668 -166815
rect 152712 -166859 152768 -166815
rect 152812 -166859 174682 -166815
rect -59794 -166915 174682 -166859
rect -59794 -166959 145268 -166915
rect 145312 -166959 145368 -166915
rect 145412 -166959 145468 -166915
rect 145512 -166959 145568 -166915
rect 145612 -166959 145668 -166915
rect 145712 -166959 145768 -166915
rect 145812 -166959 145868 -166915
rect 145912 -166959 145968 -166915
rect 146012 -166959 146068 -166915
rect 146112 -166959 146168 -166915
rect 146212 -166959 146268 -166915
rect 146312 -166959 146368 -166915
rect 146412 -166959 146468 -166915
rect 146512 -166959 146568 -166915
rect 146612 -166959 146668 -166915
rect 146712 -166959 146768 -166915
rect 146812 -166959 147268 -166915
rect 147312 -166959 147368 -166915
rect 147412 -166959 147468 -166915
rect 147512 -166959 147568 -166915
rect 147612 -166959 147668 -166915
rect 147712 -166959 147768 -166915
rect 147812 -166959 147868 -166915
rect 147912 -166959 147968 -166915
rect 148012 -166959 148068 -166915
rect 148112 -166959 148168 -166915
rect 148212 -166959 148268 -166915
rect 148312 -166959 148368 -166915
rect 148412 -166959 148468 -166915
rect 148512 -166959 148568 -166915
rect 148612 -166959 148668 -166915
rect 148712 -166959 148768 -166915
rect 148812 -166959 149268 -166915
rect 149312 -166959 149368 -166915
rect 149412 -166959 149468 -166915
rect 149512 -166959 149568 -166915
rect 149612 -166959 149668 -166915
rect 149712 -166959 149768 -166915
rect 149812 -166959 149868 -166915
rect 149912 -166959 149968 -166915
rect 150012 -166959 150068 -166915
rect 150112 -166959 150168 -166915
rect 150212 -166959 150268 -166915
rect 150312 -166959 150368 -166915
rect 150412 -166959 150468 -166915
rect 150512 -166959 150568 -166915
rect 150612 -166959 150668 -166915
rect 150712 -166959 150768 -166915
rect 150812 -166959 151268 -166915
rect 151312 -166959 151368 -166915
rect 151412 -166959 151468 -166915
rect 151512 -166959 151568 -166915
rect 151612 -166959 151668 -166915
rect 151712 -166959 151768 -166915
rect 151812 -166959 151868 -166915
rect 151912 -166959 151968 -166915
rect 152012 -166959 152068 -166915
rect 152112 -166959 152168 -166915
rect 152212 -166959 152268 -166915
rect 152312 -166959 152368 -166915
rect 152412 -166959 152468 -166915
rect 152512 -166959 152568 -166915
rect 152612 -166959 152668 -166915
rect 152712 -166959 152768 -166915
rect 152812 -166959 174682 -166915
rect -59794 -167015 174682 -166959
rect -59794 -167059 145268 -167015
rect 145312 -167059 145368 -167015
rect 145412 -167059 145468 -167015
rect 145512 -167059 145568 -167015
rect 145612 -167059 145668 -167015
rect 145712 -167059 145768 -167015
rect 145812 -167059 145868 -167015
rect 145912 -167059 145968 -167015
rect 146012 -167059 146068 -167015
rect 146112 -167059 146168 -167015
rect 146212 -167059 146268 -167015
rect 146312 -167059 146368 -167015
rect 146412 -167059 146468 -167015
rect 146512 -167059 146568 -167015
rect 146612 -167059 146668 -167015
rect 146712 -167059 146768 -167015
rect 146812 -167059 147268 -167015
rect 147312 -167059 147368 -167015
rect 147412 -167059 147468 -167015
rect 147512 -167059 147568 -167015
rect 147612 -167059 147668 -167015
rect 147712 -167059 147768 -167015
rect 147812 -167059 147868 -167015
rect 147912 -167059 147968 -167015
rect 148012 -167059 148068 -167015
rect 148112 -167059 148168 -167015
rect 148212 -167059 148268 -167015
rect 148312 -167059 148368 -167015
rect 148412 -167059 148468 -167015
rect 148512 -167059 148568 -167015
rect 148612 -167059 148668 -167015
rect 148712 -167059 148768 -167015
rect 148812 -167059 149268 -167015
rect 149312 -167059 149368 -167015
rect 149412 -167059 149468 -167015
rect 149512 -167059 149568 -167015
rect 149612 -167059 149668 -167015
rect 149712 -167059 149768 -167015
rect 149812 -167059 149868 -167015
rect 149912 -167059 149968 -167015
rect 150012 -167059 150068 -167015
rect 150112 -167059 150168 -167015
rect 150212 -167059 150268 -167015
rect 150312 -167059 150368 -167015
rect 150412 -167059 150468 -167015
rect 150512 -167059 150568 -167015
rect 150612 -167059 150668 -167015
rect 150712 -167059 150768 -167015
rect 150812 -167059 151268 -167015
rect 151312 -167059 151368 -167015
rect 151412 -167059 151468 -167015
rect 151512 -167059 151568 -167015
rect 151612 -167059 151668 -167015
rect 151712 -167059 151768 -167015
rect 151812 -167059 151868 -167015
rect 151912 -167059 151968 -167015
rect 152012 -167059 152068 -167015
rect 152112 -167059 152168 -167015
rect 152212 -167059 152268 -167015
rect 152312 -167059 152368 -167015
rect 152412 -167059 152468 -167015
rect 152512 -167059 152568 -167015
rect 152612 -167059 152668 -167015
rect 152712 -167059 152768 -167015
rect 152812 -167059 174682 -167015
rect -59794 -167115 174682 -167059
rect -59794 -167159 145268 -167115
rect 145312 -167159 145368 -167115
rect 145412 -167159 145468 -167115
rect 145512 -167159 145568 -167115
rect 145612 -167159 145668 -167115
rect 145712 -167159 145768 -167115
rect 145812 -167159 145868 -167115
rect 145912 -167159 145968 -167115
rect 146012 -167159 146068 -167115
rect 146112 -167159 146168 -167115
rect 146212 -167159 146268 -167115
rect 146312 -167159 146368 -167115
rect 146412 -167159 146468 -167115
rect 146512 -167159 146568 -167115
rect 146612 -167159 146668 -167115
rect 146712 -167159 146768 -167115
rect 146812 -167159 147268 -167115
rect 147312 -167159 147368 -167115
rect 147412 -167159 147468 -167115
rect 147512 -167159 147568 -167115
rect 147612 -167159 147668 -167115
rect 147712 -167159 147768 -167115
rect 147812 -167159 147868 -167115
rect 147912 -167159 147968 -167115
rect 148012 -167159 148068 -167115
rect 148112 -167159 148168 -167115
rect 148212 -167159 148268 -167115
rect 148312 -167159 148368 -167115
rect 148412 -167159 148468 -167115
rect 148512 -167159 148568 -167115
rect 148612 -167159 148668 -167115
rect 148712 -167159 148768 -167115
rect 148812 -167159 149268 -167115
rect 149312 -167159 149368 -167115
rect 149412 -167159 149468 -167115
rect 149512 -167159 149568 -167115
rect 149612 -167159 149668 -167115
rect 149712 -167159 149768 -167115
rect 149812 -167159 149868 -167115
rect 149912 -167159 149968 -167115
rect 150012 -167159 150068 -167115
rect 150112 -167159 150168 -167115
rect 150212 -167159 150268 -167115
rect 150312 -167159 150368 -167115
rect 150412 -167159 150468 -167115
rect 150512 -167159 150568 -167115
rect 150612 -167159 150668 -167115
rect 150712 -167159 150768 -167115
rect 150812 -167159 151268 -167115
rect 151312 -167159 151368 -167115
rect 151412 -167159 151468 -167115
rect 151512 -167159 151568 -167115
rect 151612 -167159 151668 -167115
rect 151712 -167159 151768 -167115
rect 151812 -167159 151868 -167115
rect 151912 -167159 151968 -167115
rect 152012 -167159 152068 -167115
rect 152112 -167159 152168 -167115
rect 152212 -167159 152268 -167115
rect 152312 -167159 152368 -167115
rect 152412 -167159 152468 -167115
rect 152512 -167159 152568 -167115
rect 152612 -167159 152668 -167115
rect 152712 -167159 152768 -167115
rect 152812 -167159 174682 -167115
rect -59794 -168689 174682 -167159
rect -114442 -172989 178472 -171279
rect -114442 -173033 165525 -172989
rect 165569 -173033 165625 -172989
rect 165669 -173033 165725 -172989
rect 165769 -173033 165825 -172989
rect 165869 -173033 165925 -172989
rect 165969 -173033 166025 -172989
rect 166069 -173033 166125 -172989
rect 166169 -173033 166225 -172989
rect 166269 -173033 166325 -172989
rect 166369 -173033 166425 -172989
rect 166469 -173033 166525 -172989
rect 166569 -173033 166625 -172989
rect 166669 -173033 166725 -172989
rect 166769 -173033 166825 -172989
rect 166869 -173033 166925 -172989
rect 166969 -173033 167025 -172989
rect 167069 -173033 167525 -172989
rect 167569 -173033 167625 -172989
rect 167669 -173033 167725 -172989
rect 167769 -173033 167825 -172989
rect 167869 -173033 167925 -172989
rect 167969 -173033 168025 -172989
rect 168069 -173033 168125 -172989
rect 168169 -173033 168225 -172989
rect 168269 -173033 168325 -172989
rect 168369 -173033 168425 -172989
rect 168469 -173033 168525 -172989
rect 168569 -173033 168625 -172989
rect 168669 -173033 168725 -172989
rect 168769 -173033 168825 -172989
rect 168869 -173033 168925 -172989
rect 168969 -173033 169025 -172989
rect 169069 -173033 169525 -172989
rect 169569 -173033 169625 -172989
rect 169669 -173033 169725 -172989
rect 169769 -173033 169825 -172989
rect 169869 -173033 169925 -172989
rect 169969 -173033 170025 -172989
rect 170069 -173033 170125 -172989
rect 170169 -173033 170225 -172989
rect 170269 -173033 170325 -172989
rect 170369 -173033 170425 -172989
rect 170469 -173033 170525 -172989
rect 170569 -173033 170625 -172989
rect 170669 -173033 170725 -172989
rect 170769 -173033 170825 -172989
rect 170869 -173033 170925 -172989
rect 170969 -173033 171025 -172989
rect 171069 -173033 171525 -172989
rect 171569 -173033 171625 -172989
rect 171669 -173033 171725 -172989
rect 171769 -173033 171825 -172989
rect 171869 -173033 171925 -172989
rect 171969 -173033 172025 -172989
rect 172069 -173033 172125 -172989
rect 172169 -173033 172225 -172989
rect 172269 -173033 172325 -172989
rect 172369 -173033 172425 -172989
rect 172469 -173033 172525 -172989
rect 172569 -173033 172625 -172989
rect 172669 -173033 172725 -172989
rect 172769 -173033 172825 -172989
rect 172869 -173033 172925 -172989
rect 172969 -173033 173025 -172989
rect 173069 -173033 178472 -172989
rect -114442 -173049 178472 -173033
rect -114442 -173093 81627 -173049
rect 81671 -173093 81727 -173049
rect 81771 -173093 81827 -173049
rect 81871 -173093 81927 -173049
rect 81971 -173093 82027 -173049
rect 82071 -173093 82127 -173049
rect 82171 -173093 82227 -173049
rect 82271 -173093 82327 -173049
rect 82371 -173093 82427 -173049
rect 82471 -173093 82527 -173049
rect 82571 -173093 82627 -173049
rect 82671 -173093 82727 -173049
rect 82771 -173093 82827 -173049
rect 82871 -173093 82927 -173049
rect 82971 -173093 83027 -173049
rect 83071 -173093 83127 -173049
rect 83171 -173093 83627 -173049
rect 83671 -173093 83727 -173049
rect 83771 -173093 83827 -173049
rect 83871 -173093 83927 -173049
rect 83971 -173093 84027 -173049
rect 84071 -173093 84127 -173049
rect 84171 -173093 84227 -173049
rect 84271 -173093 84327 -173049
rect 84371 -173093 84427 -173049
rect 84471 -173093 84527 -173049
rect 84571 -173093 84627 -173049
rect 84671 -173093 84727 -173049
rect 84771 -173093 84827 -173049
rect 84871 -173093 84927 -173049
rect 84971 -173093 85027 -173049
rect 85071 -173093 85127 -173049
rect 85171 -173093 85627 -173049
rect 85671 -173093 85727 -173049
rect 85771 -173093 85827 -173049
rect 85871 -173093 85927 -173049
rect 85971 -173093 86027 -173049
rect 86071 -173093 86127 -173049
rect 86171 -173093 86227 -173049
rect 86271 -173093 86327 -173049
rect 86371 -173093 86427 -173049
rect 86471 -173093 86527 -173049
rect 86571 -173093 86627 -173049
rect 86671 -173093 86727 -173049
rect 86771 -173093 86827 -173049
rect 86871 -173093 86927 -173049
rect 86971 -173093 87027 -173049
rect 87071 -173093 87127 -173049
rect 87171 -173093 87627 -173049
rect 87671 -173093 87727 -173049
rect 87771 -173093 87827 -173049
rect 87871 -173093 87927 -173049
rect 87971 -173093 88027 -173049
rect 88071 -173093 88127 -173049
rect 88171 -173093 88227 -173049
rect 88271 -173093 88327 -173049
rect 88371 -173093 88427 -173049
rect 88471 -173093 88527 -173049
rect 88571 -173093 88627 -173049
rect 88671 -173093 88727 -173049
rect 88771 -173093 88827 -173049
rect 88871 -173093 88927 -173049
rect 88971 -173093 89027 -173049
rect 89071 -173093 89127 -173049
rect 89171 -173089 178472 -173049
rect 89171 -173093 165525 -173089
rect -114442 -173133 165525 -173093
rect 165569 -173133 165625 -173089
rect 165669 -173133 165725 -173089
rect 165769 -173133 165825 -173089
rect 165869 -173133 165925 -173089
rect 165969 -173133 166025 -173089
rect 166069 -173133 166125 -173089
rect 166169 -173133 166225 -173089
rect 166269 -173133 166325 -173089
rect 166369 -173133 166425 -173089
rect 166469 -173133 166525 -173089
rect 166569 -173133 166625 -173089
rect 166669 -173133 166725 -173089
rect 166769 -173133 166825 -173089
rect 166869 -173133 166925 -173089
rect 166969 -173133 167025 -173089
rect 167069 -173133 167525 -173089
rect 167569 -173133 167625 -173089
rect 167669 -173133 167725 -173089
rect 167769 -173133 167825 -173089
rect 167869 -173133 167925 -173089
rect 167969 -173133 168025 -173089
rect 168069 -173133 168125 -173089
rect 168169 -173133 168225 -173089
rect 168269 -173133 168325 -173089
rect 168369 -173133 168425 -173089
rect 168469 -173133 168525 -173089
rect 168569 -173133 168625 -173089
rect 168669 -173133 168725 -173089
rect 168769 -173133 168825 -173089
rect 168869 -173133 168925 -173089
rect 168969 -173133 169025 -173089
rect 169069 -173133 169525 -173089
rect 169569 -173133 169625 -173089
rect 169669 -173133 169725 -173089
rect 169769 -173133 169825 -173089
rect 169869 -173133 169925 -173089
rect 169969 -173133 170025 -173089
rect 170069 -173133 170125 -173089
rect 170169 -173133 170225 -173089
rect 170269 -173133 170325 -173089
rect 170369 -173133 170425 -173089
rect 170469 -173133 170525 -173089
rect 170569 -173133 170625 -173089
rect 170669 -173133 170725 -173089
rect 170769 -173133 170825 -173089
rect 170869 -173133 170925 -173089
rect 170969 -173133 171025 -173089
rect 171069 -173133 171525 -173089
rect 171569 -173133 171625 -173089
rect 171669 -173133 171725 -173089
rect 171769 -173133 171825 -173089
rect 171869 -173133 171925 -173089
rect 171969 -173133 172025 -173089
rect 172069 -173133 172125 -173089
rect 172169 -173133 172225 -173089
rect 172269 -173133 172325 -173089
rect 172369 -173133 172425 -173089
rect 172469 -173133 172525 -173089
rect 172569 -173133 172625 -173089
rect 172669 -173133 172725 -173089
rect 172769 -173133 172825 -173089
rect 172869 -173133 172925 -173089
rect 172969 -173133 173025 -173089
rect 173069 -173133 178472 -173089
rect -114442 -173149 178472 -173133
rect -114442 -173193 81627 -173149
rect 81671 -173193 81727 -173149
rect 81771 -173193 81827 -173149
rect 81871 -173193 81927 -173149
rect 81971 -173193 82027 -173149
rect 82071 -173193 82127 -173149
rect 82171 -173193 82227 -173149
rect 82271 -173193 82327 -173149
rect 82371 -173193 82427 -173149
rect 82471 -173193 82527 -173149
rect 82571 -173193 82627 -173149
rect 82671 -173193 82727 -173149
rect 82771 -173193 82827 -173149
rect 82871 -173193 82927 -173149
rect 82971 -173193 83027 -173149
rect 83071 -173193 83127 -173149
rect 83171 -173193 83627 -173149
rect 83671 -173193 83727 -173149
rect 83771 -173193 83827 -173149
rect 83871 -173193 83927 -173149
rect 83971 -173193 84027 -173149
rect 84071 -173193 84127 -173149
rect 84171 -173193 84227 -173149
rect 84271 -173193 84327 -173149
rect 84371 -173193 84427 -173149
rect 84471 -173193 84527 -173149
rect 84571 -173193 84627 -173149
rect 84671 -173193 84727 -173149
rect 84771 -173193 84827 -173149
rect 84871 -173193 84927 -173149
rect 84971 -173193 85027 -173149
rect 85071 -173193 85127 -173149
rect 85171 -173193 85627 -173149
rect 85671 -173193 85727 -173149
rect 85771 -173193 85827 -173149
rect 85871 -173193 85927 -173149
rect 85971 -173193 86027 -173149
rect 86071 -173193 86127 -173149
rect 86171 -173193 86227 -173149
rect 86271 -173193 86327 -173149
rect 86371 -173193 86427 -173149
rect 86471 -173193 86527 -173149
rect 86571 -173193 86627 -173149
rect 86671 -173193 86727 -173149
rect 86771 -173193 86827 -173149
rect 86871 -173193 86927 -173149
rect 86971 -173193 87027 -173149
rect 87071 -173193 87127 -173149
rect 87171 -173193 87627 -173149
rect 87671 -173193 87727 -173149
rect 87771 -173193 87827 -173149
rect 87871 -173193 87927 -173149
rect 87971 -173193 88027 -173149
rect 88071 -173193 88127 -173149
rect 88171 -173193 88227 -173149
rect 88271 -173193 88327 -173149
rect 88371 -173193 88427 -173149
rect 88471 -173193 88527 -173149
rect 88571 -173193 88627 -173149
rect 88671 -173193 88727 -173149
rect 88771 -173193 88827 -173149
rect 88871 -173193 88927 -173149
rect 88971 -173193 89027 -173149
rect 89071 -173193 89127 -173149
rect 89171 -173189 178472 -173149
rect 89171 -173193 165525 -173189
rect -114442 -173233 165525 -173193
rect 165569 -173233 165625 -173189
rect 165669 -173233 165725 -173189
rect 165769 -173233 165825 -173189
rect 165869 -173233 165925 -173189
rect 165969 -173233 166025 -173189
rect 166069 -173233 166125 -173189
rect 166169 -173233 166225 -173189
rect 166269 -173233 166325 -173189
rect 166369 -173233 166425 -173189
rect 166469 -173233 166525 -173189
rect 166569 -173233 166625 -173189
rect 166669 -173233 166725 -173189
rect 166769 -173233 166825 -173189
rect 166869 -173233 166925 -173189
rect 166969 -173233 167025 -173189
rect 167069 -173233 167525 -173189
rect 167569 -173233 167625 -173189
rect 167669 -173233 167725 -173189
rect 167769 -173233 167825 -173189
rect 167869 -173233 167925 -173189
rect 167969 -173233 168025 -173189
rect 168069 -173233 168125 -173189
rect 168169 -173233 168225 -173189
rect 168269 -173233 168325 -173189
rect 168369 -173233 168425 -173189
rect 168469 -173233 168525 -173189
rect 168569 -173233 168625 -173189
rect 168669 -173233 168725 -173189
rect 168769 -173233 168825 -173189
rect 168869 -173233 168925 -173189
rect 168969 -173233 169025 -173189
rect 169069 -173233 169525 -173189
rect 169569 -173233 169625 -173189
rect 169669 -173233 169725 -173189
rect 169769 -173233 169825 -173189
rect 169869 -173233 169925 -173189
rect 169969 -173233 170025 -173189
rect 170069 -173233 170125 -173189
rect 170169 -173233 170225 -173189
rect 170269 -173233 170325 -173189
rect 170369 -173233 170425 -173189
rect 170469 -173233 170525 -173189
rect 170569 -173233 170625 -173189
rect 170669 -173233 170725 -173189
rect 170769 -173233 170825 -173189
rect 170869 -173233 170925 -173189
rect 170969 -173233 171025 -173189
rect 171069 -173233 171525 -173189
rect 171569 -173233 171625 -173189
rect 171669 -173233 171725 -173189
rect 171769 -173233 171825 -173189
rect 171869 -173233 171925 -173189
rect 171969 -173233 172025 -173189
rect 172069 -173233 172125 -173189
rect 172169 -173233 172225 -173189
rect 172269 -173233 172325 -173189
rect 172369 -173233 172425 -173189
rect 172469 -173233 172525 -173189
rect 172569 -173233 172625 -173189
rect 172669 -173233 172725 -173189
rect 172769 -173233 172825 -173189
rect 172869 -173233 172925 -173189
rect 172969 -173233 173025 -173189
rect 173069 -173233 178472 -173189
rect -114442 -173249 178472 -173233
rect -114442 -173293 81627 -173249
rect 81671 -173293 81727 -173249
rect 81771 -173293 81827 -173249
rect 81871 -173293 81927 -173249
rect 81971 -173293 82027 -173249
rect 82071 -173293 82127 -173249
rect 82171 -173293 82227 -173249
rect 82271 -173293 82327 -173249
rect 82371 -173293 82427 -173249
rect 82471 -173293 82527 -173249
rect 82571 -173293 82627 -173249
rect 82671 -173293 82727 -173249
rect 82771 -173293 82827 -173249
rect 82871 -173293 82927 -173249
rect 82971 -173293 83027 -173249
rect 83071 -173293 83127 -173249
rect 83171 -173293 83627 -173249
rect 83671 -173293 83727 -173249
rect 83771 -173293 83827 -173249
rect 83871 -173293 83927 -173249
rect 83971 -173293 84027 -173249
rect 84071 -173293 84127 -173249
rect 84171 -173293 84227 -173249
rect 84271 -173293 84327 -173249
rect 84371 -173293 84427 -173249
rect 84471 -173293 84527 -173249
rect 84571 -173293 84627 -173249
rect 84671 -173293 84727 -173249
rect 84771 -173293 84827 -173249
rect 84871 -173293 84927 -173249
rect 84971 -173293 85027 -173249
rect 85071 -173293 85127 -173249
rect 85171 -173293 85627 -173249
rect 85671 -173293 85727 -173249
rect 85771 -173293 85827 -173249
rect 85871 -173293 85927 -173249
rect 85971 -173293 86027 -173249
rect 86071 -173293 86127 -173249
rect 86171 -173293 86227 -173249
rect 86271 -173293 86327 -173249
rect 86371 -173293 86427 -173249
rect 86471 -173293 86527 -173249
rect 86571 -173293 86627 -173249
rect 86671 -173293 86727 -173249
rect 86771 -173293 86827 -173249
rect 86871 -173293 86927 -173249
rect 86971 -173293 87027 -173249
rect 87071 -173293 87127 -173249
rect 87171 -173293 87627 -173249
rect 87671 -173293 87727 -173249
rect 87771 -173293 87827 -173249
rect 87871 -173293 87927 -173249
rect 87971 -173293 88027 -173249
rect 88071 -173293 88127 -173249
rect 88171 -173293 88227 -173249
rect 88271 -173293 88327 -173249
rect 88371 -173293 88427 -173249
rect 88471 -173293 88527 -173249
rect 88571 -173293 88627 -173249
rect 88671 -173293 88727 -173249
rect 88771 -173293 88827 -173249
rect 88871 -173293 88927 -173249
rect 88971 -173293 89027 -173249
rect 89071 -173293 89127 -173249
rect 89171 -173289 178472 -173249
rect 89171 -173293 165525 -173289
rect -114442 -173333 165525 -173293
rect 165569 -173333 165625 -173289
rect 165669 -173333 165725 -173289
rect 165769 -173333 165825 -173289
rect 165869 -173333 165925 -173289
rect 165969 -173333 166025 -173289
rect 166069 -173333 166125 -173289
rect 166169 -173333 166225 -173289
rect 166269 -173333 166325 -173289
rect 166369 -173333 166425 -173289
rect 166469 -173333 166525 -173289
rect 166569 -173333 166625 -173289
rect 166669 -173333 166725 -173289
rect 166769 -173333 166825 -173289
rect 166869 -173333 166925 -173289
rect 166969 -173333 167025 -173289
rect 167069 -173333 167525 -173289
rect 167569 -173333 167625 -173289
rect 167669 -173333 167725 -173289
rect 167769 -173333 167825 -173289
rect 167869 -173333 167925 -173289
rect 167969 -173333 168025 -173289
rect 168069 -173333 168125 -173289
rect 168169 -173333 168225 -173289
rect 168269 -173333 168325 -173289
rect 168369 -173333 168425 -173289
rect 168469 -173333 168525 -173289
rect 168569 -173333 168625 -173289
rect 168669 -173333 168725 -173289
rect 168769 -173333 168825 -173289
rect 168869 -173333 168925 -173289
rect 168969 -173333 169025 -173289
rect 169069 -173333 169525 -173289
rect 169569 -173333 169625 -173289
rect 169669 -173333 169725 -173289
rect 169769 -173333 169825 -173289
rect 169869 -173333 169925 -173289
rect 169969 -173333 170025 -173289
rect 170069 -173333 170125 -173289
rect 170169 -173333 170225 -173289
rect 170269 -173333 170325 -173289
rect 170369 -173333 170425 -173289
rect 170469 -173333 170525 -173289
rect 170569 -173333 170625 -173289
rect 170669 -173333 170725 -173289
rect 170769 -173333 170825 -173289
rect 170869 -173333 170925 -173289
rect 170969 -173333 171025 -173289
rect 171069 -173333 171525 -173289
rect 171569 -173333 171625 -173289
rect 171669 -173333 171725 -173289
rect 171769 -173333 171825 -173289
rect 171869 -173333 171925 -173289
rect 171969 -173333 172025 -173289
rect 172069 -173333 172125 -173289
rect 172169 -173333 172225 -173289
rect 172269 -173333 172325 -173289
rect 172369 -173333 172425 -173289
rect 172469 -173333 172525 -173289
rect 172569 -173333 172625 -173289
rect 172669 -173333 172725 -173289
rect 172769 -173333 172825 -173289
rect 172869 -173333 172925 -173289
rect 172969 -173333 173025 -173289
rect 173069 -173333 178472 -173289
rect -114442 -173349 178472 -173333
rect -114442 -173393 81627 -173349
rect 81671 -173393 81727 -173349
rect 81771 -173393 81827 -173349
rect 81871 -173393 81927 -173349
rect 81971 -173393 82027 -173349
rect 82071 -173393 82127 -173349
rect 82171 -173393 82227 -173349
rect 82271 -173393 82327 -173349
rect 82371 -173393 82427 -173349
rect 82471 -173393 82527 -173349
rect 82571 -173393 82627 -173349
rect 82671 -173393 82727 -173349
rect 82771 -173393 82827 -173349
rect 82871 -173393 82927 -173349
rect 82971 -173393 83027 -173349
rect 83071 -173393 83127 -173349
rect 83171 -173393 83627 -173349
rect 83671 -173393 83727 -173349
rect 83771 -173393 83827 -173349
rect 83871 -173393 83927 -173349
rect 83971 -173393 84027 -173349
rect 84071 -173393 84127 -173349
rect 84171 -173393 84227 -173349
rect 84271 -173393 84327 -173349
rect 84371 -173393 84427 -173349
rect 84471 -173393 84527 -173349
rect 84571 -173393 84627 -173349
rect 84671 -173393 84727 -173349
rect 84771 -173393 84827 -173349
rect 84871 -173393 84927 -173349
rect 84971 -173393 85027 -173349
rect 85071 -173393 85127 -173349
rect 85171 -173393 85627 -173349
rect 85671 -173393 85727 -173349
rect 85771 -173393 85827 -173349
rect 85871 -173393 85927 -173349
rect 85971 -173393 86027 -173349
rect 86071 -173393 86127 -173349
rect 86171 -173393 86227 -173349
rect 86271 -173393 86327 -173349
rect 86371 -173393 86427 -173349
rect 86471 -173393 86527 -173349
rect 86571 -173393 86627 -173349
rect 86671 -173393 86727 -173349
rect 86771 -173393 86827 -173349
rect 86871 -173393 86927 -173349
rect 86971 -173393 87027 -173349
rect 87071 -173393 87127 -173349
rect 87171 -173393 87627 -173349
rect 87671 -173393 87727 -173349
rect 87771 -173393 87827 -173349
rect 87871 -173393 87927 -173349
rect 87971 -173393 88027 -173349
rect 88071 -173393 88127 -173349
rect 88171 -173393 88227 -173349
rect 88271 -173393 88327 -173349
rect 88371 -173393 88427 -173349
rect 88471 -173393 88527 -173349
rect 88571 -173393 88627 -173349
rect 88671 -173393 88727 -173349
rect 88771 -173393 88827 -173349
rect 88871 -173393 88927 -173349
rect 88971 -173393 89027 -173349
rect 89071 -173393 89127 -173349
rect 89171 -173389 178472 -173349
rect 89171 -173393 165525 -173389
rect -114442 -173433 165525 -173393
rect 165569 -173433 165625 -173389
rect 165669 -173433 165725 -173389
rect 165769 -173433 165825 -173389
rect 165869 -173433 165925 -173389
rect 165969 -173433 166025 -173389
rect 166069 -173433 166125 -173389
rect 166169 -173433 166225 -173389
rect 166269 -173433 166325 -173389
rect 166369 -173433 166425 -173389
rect 166469 -173433 166525 -173389
rect 166569 -173433 166625 -173389
rect 166669 -173433 166725 -173389
rect 166769 -173433 166825 -173389
rect 166869 -173433 166925 -173389
rect 166969 -173433 167025 -173389
rect 167069 -173433 167525 -173389
rect 167569 -173433 167625 -173389
rect 167669 -173433 167725 -173389
rect 167769 -173433 167825 -173389
rect 167869 -173433 167925 -173389
rect 167969 -173433 168025 -173389
rect 168069 -173433 168125 -173389
rect 168169 -173433 168225 -173389
rect 168269 -173433 168325 -173389
rect 168369 -173433 168425 -173389
rect 168469 -173433 168525 -173389
rect 168569 -173433 168625 -173389
rect 168669 -173433 168725 -173389
rect 168769 -173433 168825 -173389
rect 168869 -173433 168925 -173389
rect 168969 -173433 169025 -173389
rect 169069 -173433 169525 -173389
rect 169569 -173433 169625 -173389
rect 169669 -173433 169725 -173389
rect 169769 -173433 169825 -173389
rect 169869 -173433 169925 -173389
rect 169969 -173433 170025 -173389
rect 170069 -173433 170125 -173389
rect 170169 -173433 170225 -173389
rect 170269 -173433 170325 -173389
rect 170369 -173433 170425 -173389
rect 170469 -173433 170525 -173389
rect 170569 -173433 170625 -173389
rect 170669 -173433 170725 -173389
rect 170769 -173433 170825 -173389
rect 170869 -173433 170925 -173389
rect 170969 -173433 171025 -173389
rect 171069 -173433 171525 -173389
rect 171569 -173433 171625 -173389
rect 171669 -173433 171725 -173389
rect 171769 -173433 171825 -173389
rect 171869 -173433 171925 -173389
rect 171969 -173433 172025 -173389
rect 172069 -173433 172125 -173389
rect 172169 -173433 172225 -173389
rect 172269 -173433 172325 -173389
rect 172369 -173433 172425 -173389
rect 172469 -173433 172525 -173389
rect 172569 -173433 172625 -173389
rect 172669 -173433 172725 -173389
rect 172769 -173433 172825 -173389
rect 172869 -173433 172925 -173389
rect 172969 -173433 173025 -173389
rect 173069 -173433 178472 -173389
rect -114442 -173449 178472 -173433
rect -114442 -173493 81627 -173449
rect 81671 -173493 81727 -173449
rect 81771 -173493 81827 -173449
rect 81871 -173493 81927 -173449
rect 81971 -173493 82027 -173449
rect 82071 -173493 82127 -173449
rect 82171 -173493 82227 -173449
rect 82271 -173493 82327 -173449
rect 82371 -173493 82427 -173449
rect 82471 -173493 82527 -173449
rect 82571 -173493 82627 -173449
rect 82671 -173493 82727 -173449
rect 82771 -173493 82827 -173449
rect 82871 -173493 82927 -173449
rect 82971 -173493 83027 -173449
rect 83071 -173493 83127 -173449
rect 83171 -173493 83627 -173449
rect 83671 -173493 83727 -173449
rect 83771 -173493 83827 -173449
rect 83871 -173493 83927 -173449
rect 83971 -173493 84027 -173449
rect 84071 -173493 84127 -173449
rect 84171 -173493 84227 -173449
rect 84271 -173493 84327 -173449
rect 84371 -173493 84427 -173449
rect 84471 -173493 84527 -173449
rect 84571 -173493 84627 -173449
rect 84671 -173493 84727 -173449
rect 84771 -173493 84827 -173449
rect 84871 -173493 84927 -173449
rect 84971 -173493 85027 -173449
rect 85071 -173493 85127 -173449
rect 85171 -173493 85627 -173449
rect 85671 -173493 85727 -173449
rect 85771 -173493 85827 -173449
rect 85871 -173493 85927 -173449
rect 85971 -173493 86027 -173449
rect 86071 -173493 86127 -173449
rect 86171 -173493 86227 -173449
rect 86271 -173493 86327 -173449
rect 86371 -173493 86427 -173449
rect 86471 -173493 86527 -173449
rect 86571 -173493 86627 -173449
rect 86671 -173493 86727 -173449
rect 86771 -173493 86827 -173449
rect 86871 -173493 86927 -173449
rect 86971 -173493 87027 -173449
rect 87071 -173493 87127 -173449
rect 87171 -173493 87627 -173449
rect 87671 -173493 87727 -173449
rect 87771 -173493 87827 -173449
rect 87871 -173493 87927 -173449
rect 87971 -173493 88027 -173449
rect 88071 -173493 88127 -173449
rect 88171 -173493 88227 -173449
rect 88271 -173493 88327 -173449
rect 88371 -173493 88427 -173449
rect 88471 -173493 88527 -173449
rect 88571 -173493 88627 -173449
rect 88671 -173493 88727 -173449
rect 88771 -173493 88827 -173449
rect 88871 -173493 88927 -173449
rect 88971 -173493 89027 -173449
rect 89071 -173493 89127 -173449
rect 89171 -173489 178472 -173449
rect 89171 -173493 165525 -173489
rect -114442 -173533 165525 -173493
rect 165569 -173533 165625 -173489
rect 165669 -173533 165725 -173489
rect 165769 -173533 165825 -173489
rect 165869 -173533 165925 -173489
rect 165969 -173533 166025 -173489
rect 166069 -173533 166125 -173489
rect 166169 -173533 166225 -173489
rect 166269 -173533 166325 -173489
rect 166369 -173533 166425 -173489
rect 166469 -173533 166525 -173489
rect 166569 -173533 166625 -173489
rect 166669 -173533 166725 -173489
rect 166769 -173533 166825 -173489
rect 166869 -173533 166925 -173489
rect 166969 -173533 167025 -173489
rect 167069 -173533 167525 -173489
rect 167569 -173533 167625 -173489
rect 167669 -173533 167725 -173489
rect 167769 -173533 167825 -173489
rect 167869 -173533 167925 -173489
rect 167969 -173533 168025 -173489
rect 168069 -173533 168125 -173489
rect 168169 -173533 168225 -173489
rect 168269 -173533 168325 -173489
rect 168369 -173533 168425 -173489
rect 168469 -173533 168525 -173489
rect 168569 -173533 168625 -173489
rect 168669 -173533 168725 -173489
rect 168769 -173533 168825 -173489
rect 168869 -173533 168925 -173489
rect 168969 -173533 169025 -173489
rect 169069 -173533 169525 -173489
rect 169569 -173533 169625 -173489
rect 169669 -173533 169725 -173489
rect 169769 -173533 169825 -173489
rect 169869 -173533 169925 -173489
rect 169969 -173533 170025 -173489
rect 170069 -173533 170125 -173489
rect 170169 -173533 170225 -173489
rect 170269 -173533 170325 -173489
rect 170369 -173533 170425 -173489
rect 170469 -173533 170525 -173489
rect 170569 -173533 170625 -173489
rect 170669 -173533 170725 -173489
rect 170769 -173533 170825 -173489
rect 170869 -173533 170925 -173489
rect 170969 -173533 171025 -173489
rect 171069 -173533 171525 -173489
rect 171569 -173533 171625 -173489
rect 171669 -173533 171725 -173489
rect 171769 -173533 171825 -173489
rect 171869 -173533 171925 -173489
rect 171969 -173533 172025 -173489
rect 172069 -173533 172125 -173489
rect 172169 -173533 172225 -173489
rect 172269 -173533 172325 -173489
rect 172369 -173533 172425 -173489
rect 172469 -173533 172525 -173489
rect 172569 -173533 172625 -173489
rect 172669 -173533 172725 -173489
rect 172769 -173533 172825 -173489
rect 172869 -173533 172925 -173489
rect 172969 -173533 173025 -173489
rect 173069 -173533 178472 -173489
rect -114442 -173549 178472 -173533
rect -114442 -173593 81627 -173549
rect 81671 -173593 81727 -173549
rect 81771 -173593 81827 -173549
rect 81871 -173593 81927 -173549
rect 81971 -173593 82027 -173549
rect 82071 -173593 82127 -173549
rect 82171 -173593 82227 -173549
rect 82271 -173593 82327 -173549
rect 82371 -173593 82427 -173549
rect 82471 -173593 82527 -173549
rect 82571 -173593 82627 -173549
rect 82671 -173593 82727 -173549
rect 82771 -173593 82827 -173549
rect 82871 -173593 82927 -173549
rect 82971 -173593 83027 -173549
rect 83071 -173593 83127 -173549
rect 83171 -173593 83627 -173549
rect 83671 -173593 83727 -173549
rect 83771 -173593 83827 -173549
rect 83871 -173593 83927 -173549
rect 83971 -173593 84027 -173549
rect 84071 -173593 84127 -173549
rect 84171 -173593 84227 -173549
rect 84271 -173593 84327 -173549
rect 84371 -173593 84427 -173549
rect 84471 -173593 84527 -173549
rect 84571 -173593 84627 -173549
rect 84671 -173593 84727 -173549
rect 84771 -173593 84827 -173549
rect 84871 -173593 84927 -173549
rect 84971 -173593 85027 -173549
rect 85071 -173593 85127 -173549
rect 85171 -173593 85627 -173549
rect 85671 -173593 85727 -173549
rect 85771 -173593 85827 -173549
rect 85871 -173593 85927 -173549
rect 85971 -173593 86027 -173549
rect 86071 -173593 86127 -173549
rect 86171 -173593 86227 -173549
rect 86271 -173593 86327 -173549
rect 86371 -173593 86427 -173549
rect 86471 -173593 86527 -173549
rect 86571 -173593 86627 -173549
rect 86671 -173593 86727 -173549
rect 86771 -173593 86827 -173549
rect 86871 -173593 86927 -173549
rect 86971 -173593 87027 -173549
rect 87071 -173593 87127 -173549
rect 87171 -173593 87627 -173549
rect 87671 -173593 87727 -173549
rect 87771 -173593 87827 -173549
rect 87871 -173593 87927 -173549
rect 87971 -173593 88027 -173549
rect 88071 -173593 88127 -173549
rect 88171 -173593 88227 -173549
rect 88271 -173593 88327 -173549
rect 88371 -173593 88427 -173549
rect 88471 -173593 88527 -173549
rect 88571 -173593 88627 -173549
rect 88671 -173593 88727 -173549
rect 88771 -173593 88827 -173549
rect 88871 -173593 88927 -173549
rect 88971 -173593 89027 -173549
rect 89071 -173593 89127 -173549
rect 89171 -173589 178472 -173549
rect 89171 -173593 165525 -173589
rect -114442 -173633 165525 -173593
rect 165569 -173633 165625 -173589
rect 165669 -173633 165725 -173589
rect 165769 -173633 165825 -173589
rect 165869 -173633 165925 -173589
rect 165969 -173633 166025 -173589
rect 166069 -173633 166125 -173589
rect 166169 -173633 166225 -173589
rect 166269 -173633 166325 -173589
rect 166369 -173633 166425 -173589
rect 166469 -173633 166525 -173589
rect 166569 -173633 166625 -173589
rect 166669 -173633 166725 -173589
rect 166769 -173633 166825 -173589
rect 166869 -173633 166925 -173589
rect 166969 -173633 167025 -173589
rect 167069 -173633 167525 -173589
rect 167569 -173633 167625 -173589
rect 167669 -173633 167725 -173589
rect 167769 -173633 167825 -173589
rect 167869 -173633 167925 -173589
rect 167969 -173633 168025 -173589
rect 168069 -173633 168125 -173589
rect 168169 -173633 168225 -173589
rect 168269 -173633 168325 -173589
rect 168369 -173633 168425 -173589
rect 168469 -173633 168525 -173589
rect 168569 -173633 168625 -173589
rect 168669 -173633 168725 -173589
rect 168769 -173633 168825 -173589
rect 168869 -173633 168925 -173589
rect 168969 -173633 169025 -173589
rect 169069 -173633 169525 -173589
rect 169569 -173633 169625 -173589
rect 169669 -173633 169725 -173589
rect 169769 -173633 169825 -173589
rect 169869 -173633 169925 -173589
rect 169969 -173633 170025 -173589
rect 170069 -173633 170125 -173589
rect 170169 -173633 170225 -173589
rect 170269 -173633 170325 -173589
rect 170369 -173633 170425 -173589
rect 170469 -173633 170525 -173589
rect 170569 -173633 170625 -173589
rect 170669 -173633 170725 -173589
rect 170769 -173633 170825 -173589
rect 170869 -173633 170925 -173589
rect 170969 -173633 171025 -173589
rect 171069 -173633 171525 -173589
rect 171569 -173633 171625 -173589
rect 171669 -173633 171725 -173589
rect 171769 -173633 171825 -173589
rect 171869 -173633 171925 -173589
rect 171969 -173633 172025 -173589
rect 172069 -173633 172125 -173589
rect 172169 -173633 172225 -173589
rect 172269 -173633 172325 -173589
rect 172369 -173633 172425 -173589
rect 172469 -173633 172525 -173589
rect 172569 -173633 172625 -173589
rect 172669 -173633 172725 -173589
rect 172769 -173633 172825 -173589
rect 172869 -173633 172925 -173589
rect 172969 -173633 173025 -173589
rect 173069 -173633 178472 -173589
rect -114442 -173649 178472 -173633
rect -114442 -173693 81627 -173649
rect 81671 -173693 81727 -173649
rect 81771 -173693 81827 -173649
rect 81871 -173693 81927 -173649
rect 81971 -173693 82027 -173649
rect 82071 -173693 82127 -173649
rect 82171 -173693 82227 -173649
rect 82271 -173693 82327 -173649
rect 82371 -173693 82427 -173649
rect 82471 -173693 82527 -173649
rect 82571 -173693 82627 -173649
rect 82671 -173693 82727 -173649
rect 82771 -173693 82827 -173649
rect 82871 -173693 82927 -173649
rect 82971 -173693 83027 -173649
rect 83071 -173693 83127 -173649
rect 83171 -173693 83627 -173649
rect 83671 -173693 83727 -173649
rect 83771 -173693 83827 -173649
rect 83871 -173693 83927 -173649
rect 83971 -173693 84027 -173649
rect 84071 -173693 84127 -173649
rect 84171 -173693 84227 -173649
rect 84271 -173693 84327 -173649
rect 84371 -173693 84427 -173649
rect 84471 -173693 84527 -173649
rect 84571 -173693 84627 -173649
rect 84671 -173693 84727 -173649
rect 84771 -173693 84827 -173649
rect 84871 -173693 84927 -173649
rect 84971 -173693 85027 -173649
rect 85071 -173693 85127 -173649
rect 85171 -173693 85627 -173649
rect 85671 -173693 85727 -173649
rect 85771 -173693 85827 -173649
rect 85871 -173693 85927 -173649
rect 85971 -173693 86027 -173649
rect 86071 -173693 86127 -173649
rect 86171 -173693 86227 -173649
rect 86271 -173693 86327 -173649
rect 86371 -173693 86427 -173649
rect 86471 -173693 86527 -173649
rect 86571 -173693 86627 -173649
rect 86671 -173693 86727 -173649
rect 86771 -173693 86827 -173649
rect 86871 -173693 86927 -173649
rect 86971 -173693 87027 -173649
rect 87071 -173693 87127 -173649
rect 87171 -173693 87627 -173649
rect 87671 -173693 87727 -173649
rect 87771 -173693 87827 -173649
rect 87871 -173693 87927 -173649
rect 87971 -173693 88027 -173649
rect 88071 -173693 88127 -173649
rect 88171 -173693 88227 -173649
rect 88271 -173693 88327 -173649
rect 88371 -173693 88427 -173649
rect 88471 -173693 88527 -173649
rect 88571 -173693 88627 -173649
rect 88671 -173693 88727 -173649
rect 88771 -173693 88827 -173649
rect 88871 -173693 88927 -173649
rect 88971 -173693 89027 -173649
rect 89071 -173693 89127 -173649
rect 89171 -173689 178472 -173649
rect 89171 -173693 165525 -173689
rect -114442 -173733 165525 -173693
rect 165569 -173733 165625 -173689
rect 165669 -173733 165725 -173689
rect 165769 -173733 165825 -173689
rect 165869 -173733 165925 -173689
rect 165969 -173733 166025 -173689
rect 166069 -173733 166125 -173689
rect 166169 -173733 166225 -173689
rect 166269 -173733 166325 -173689
rect 166369 -173733 166425 -173689
rect 166469 -173733 166525 -173689
rect 166569 -173733 166625 -173689
rect 166669 -173733 166725 -173689
rect 166769 -173733 166825 -173689
rect 166869 -173733 166925 -173689
rect 166969 -173733 167025 -173689
rect 167069 -173733 167525 -173689
rect 167569 -173733 167625 -173689
rect 167669 -173733 167725 -173689
rect 167769 -173733 167825 -173689
rect 167869 -173733 167925 -173689
rect 167969 -173733 168025 -173689
rect 168069 -173733 168125 -173689
rect 168169 -173733 168225 -173689
rect 168269 -173733 168325 -173689
rect 168369 -173733 168425 -173689
rect 168469 -173733 168525 -173689
rect 168569 -173733 168625 -173689
rect 168669 -173733 168725 -173689
rect 168769 -173733 168825 -173689
rect 168869 -173733 168925 -173689
rect 168969 -173733 169025 -173689
rect 169069 -173733 169525 -173689
rect 169569 -173733 169625 -173689
rect 169669 -173733 169725 -173689
rect 169769 -173733 169825 -173689
rect 169869 -173733 169925 -173689
rect 169969 -173733 170025 -173689
rect 170069 -173733 170125 -173689
rect 170169 -173733 170225 -173689
rect 170269 -173733 170325 -173689
rect 170369 -173733 170425 -173689
rect 170469 -173733 170525 -173689
rect 170569 -173733 170625 -173689
rect 170669 -173733 170725 -173689
rect 170769 -173733 170825 -173689
rect 170869 -173733 170925 -173689
rect 170969 -173733 171025 -173689
rect 171069 -173733 171525 -173689
rect 171569 -173733 171625 -173689
rect 171669 -173733 171725 -173689
rect 171769 -173733 171825 -173689
rect 171869 -173733 171925 -173689
rect 171969 -173733 172025 -173689
rect 172069 -173733 172125 -173689
rect 172169 -173733 172225 -173689
rect 172269 -173733 172325 -173689
rect 172369 -173733 172425 -173689
rect 172469 -173733 172525 -173689
rect 172569 -173733 172625 -173689
rect 172669 -173733 172725 -173689
rect 172769 -173733 172825 -173689
rect 172869 -173733 172925 -173689
rect 172969 -173733 173025 -173689
rect 173069 -173733 178472 -173689
rect -114442 -173749 178472 -173733
rect -114442 -173793 81627 -173749
rect 81671 -173793 81727 -173749
rect 81771 -173793 81827 -173749
rect 81871 -173793 81927 -173749
rect 81971 -173793 82027 -173749
rect 82071 -173793 82127 -173749
rect 82171 -173793 82227 -173749
rect 82271 -173793 82327 -173749
rect 82371 -173793 82427 -173749
rect 82471 -173793 82527 -173749
rect 82571 -173793 82627 -173749
rect 82671 -173793 82727 -173749
rect 82771 -173793 82827 -173749
rect 82871 -173793 82927 -173749
rect 82971 -173793 83027 -173749
rect 83071 -173793 83127 -173749
rect 83171 -173793 83627 -173749
rect 83671 -173793 83727 -173749
rect 83771 -173793 83827 -173749
rect 83871 -173793 83927 -173749
rect 83971 -173793 84027 -173749
rect 84071 -173793 84127 -173749
rect 84171 -173793 84227 -173749
rect 84271 -173793 84327 -173749
rect 84371 -173793 84427 -173749
rect 84471 -173793 84527 -173749
rect 84571 -173793 84627 -173749
rect 84671 -173793 84727 -173749
rect 84771 -173793 84827 -173749
rect 84871 -173793 84927 -173749
rect 84971 -173793 85027 -173749
rect 85071 -173793 85127 -173749
rect 85171 -173793 85627 -173749
rect 85671 -173793 85727 -173749
rect 85771 -173793 85827 -173749
rect 85871 -173793 85927 -173749
rect 85971 -173793 86027 -173749
rect 86071 -173793 86127 -173749
rect 86171 -173793 86227 -173749
rect 86271 -173793 86327 -173749
rect 86371 -173793 86427 -173749
rect 86471 -173793 86527 -173749
rect 86571 -173793 86627 -173749
rect 86671 -173793 86727 -173749
rect 86771 -173793 86827 -173749
rect 86871 -173793 86927 -173749
rect 86971 -173793 87027 -173749
rect 87071 -173793 87127 -173749
rect 87171 -173793 87627 -173749
rect 87671 -173793 87727 -173749
rect 87771 -173793 87827 -173749
rect 87871 -173793 87927 -173749
rect 87971 -173793 88027 -173749
rect 88071 -173793 88127 -173749
rect 88171 -173793 88227 -173749
rect 88271 -173793 88327 -173749
rect 88371 -173793 88427 -173749
rect 88471 -173793 88527 -173749
rect 88571 -173793 88627 -173749
rect 88671 -173793 88727 -173749
rect 88771 -173793 88827 -173749
rect 88871 -173793 88927 -173749
rect 88971 -173793 89027 -173749
rect 89071 -173793 89127 -173749
rect 89171 -173789 178472 -173749
rect 89171 -173793 165525 -173789
rect -114442 -173833 165525 -173793
rect 165569 -173833 165625 -173789
rect 165669 -173833 165725 -173789
rect 165769 -173833 165825 -173789
rect 165869 -173833 165925 -173789
rect 165969 -173833 166025 -173789
rect 166069 -173833 166125 -173789
rect 166169 -173833 166225 -173789
rect 166269 -173833 166325 -173789
rect 166369 -173833 166425 -173789
rect 166469 -173833 166525 -173789
rect 166569 -173833 166625 -173789
rect 166669 -173833 166725 -173789
rect 166769 -173833 166825 -173789
rect 166869 -173833 166925 -173789
rect 166969 -173833 167025 -173789
rect 167069 -173833 167525 -173789
rect 167569 -173833 167625 -173789
rect 167669 -173833 167725 -173789
rect 167769 -173833 167825 -173789
rect 167869 -173833 167925 -173789
rect 167969 -173833 168025 -173789
rect 168069 -173833 168125 -173789
rect 168169 -173833 168225 -173789
rect 168269 -173833 168325 -173789
rect 168369 -173833 168425 -173789
rect 168469 -173833 168525 -173789
rect 168569 -173833 168625 -173789
rect 168669 -173833 168725 -173789
rect 168769 -173833 168825 -173789
rect 168869 -173833 168925 -173789
rect 168969 -173833 169025 -173789
rect 169069 -173833 169525 -173789
rect 169569 -173833 169625 -173789
rect 169669 -173833 169725 -173789
rect 169769 -173833 169825 -173789
rect 169869 -173833 169925 -173789
rect 169969 -173833 170025 -173789
rect 170069 -173833 170125 -173789
rect 170169 -173833 170225 -173789
rect 170269 -173833 170325 -173789
rect 170369 -173833 170425 -173789
rect 170469 -173833 170525 -173789
rect 170569 -173833 170625 -173789
rect 170669 -173833 170725 -173789
rect 170769 -173833 170825 -173789
rect 170869 -173833 170925 -173789
rect 170969 -173833 171025 -173789
rect 171069 -173833 171525 -173789
rect 171569 -173833 171625 -173789
rect 171669 -173833 171725 -173789
rect 171769 -173833 171825 -173789
rect 171869 -173833 171925 -173789
rect 171969 -173833 172025 -173789
rect 172069 -173833 172125 -173789
rect 172169 -173833 172225 -173789
rect 172269 -173833 172325 -173789
rect 172369 -173833 172425 -173789
rect 172469 -173833 172525 -173789
rect 172569 -173833 172625 -173789
rect 172669 -173833 172725 -173789
rect 172769 -173833 172825 -173789
rect 172869 -173833 172925 -173789
rect 172969 -173833 173025 -173789
rect 173069 -173833 178472 -173789
rect -114442 -173849 178472 -173833
rect -114442 -173893 81627 -173849
rect 81671 -173893 81727 -173849
rect 81771 -173893 81827 -173849
rect 81871 -173893 81927 -173849
rect 81971 -173893 82027 -173849
rect 82071 -173893 82127 -173849
rect 82171 -173893 82227 -173849
rect 82271 -173893 82327 -173849
rect 82371 -173893 82427 -173849
rect 82471 -173893 82527 -173849
rect 82571 -173893 82627 -173849
rect 82671 -173893 82727 -173849
rect 82771 -173893 82827 -173849
rect 82871 -173893 82927 -173849
rect 82971 -173893 83027 -173849
rect 83071 -173893 83127 -173849
rect 83171 -173893 83627 -173849
rect 83671 -173893 83727 -173849
rect 83771 -173893 83827 -173849
rect 83871 -173893 83927 -173849
rect 83971 -173893 84027 -173849
rect 84071 -173893 84127 -173849
rect 84171 -173893 84227 -173849
rect 84271 -173893 84327 -173849
rect 84371 -173893 84427 -173849
rect 84471 -173893 84527 -173849
rect 84571 -173893 84627 -173849
rect 84671 -173893 84727 -173849
rect 84771 -173893 84827 -173849
rect 84871 -173893 84927 -173849
rect 84971 -173893 85027 -173849
rect 85071 -173893 85127 -173849
rect 85171 -173893 85627 -173849
rect 85671 -173893 85727 -173849
rect 85771 -173893 85827 -173849
rect 85871 -173893 85927 -173849
rect 85971 -173893 86027 -173849
rect 86071 -173893 86127 -173849
rect 86171 -173893 86227 -173849
rect 86271 -173893 86327 -173849
rect 86371 -173893 86427 -173849
rect 86471 -173893 86527 -173849
rect 86571 -173893 86627 -173849
rect 86671 -173893 86727 -173849
rect 86771 -173893 86827 -173849
rect 86871 -173893 86927 -173849
rect 86971 -173893 87027 -173849
rect 87071 -173893 87127 -173849
rect 87171 -173893 87627 -173849
rect 87671 -173893 87727 -173849
rect 87771 -173893 87827 -173849
rect 87871 -173893 87927 -173849
rect 87971 -173893 88027 -173849
rect 88071 -173893 88127 -173849
rect 88171 -173893 88227 -173849
rect 88271 -173893 88327 -173849
rect 88371 -173893 88427 -173849
rect 88471 -173893 88527 -173849
rect 88571 -173893 88627 -173849
rect 88671 -173893 88727 -173849
rect 88771 -173893 88827 -173849
rect 88871 -173893 88927 -173849
rect 88971 -173893 89027 -173849
rect 89071 -173893 89127 -173849
rect 89171 -173889 178472 -173849
rect 89171 -173893 165525 -173889
rect -114442 -173933 165525 -173893
rect 165569 -173933 165625 -173889
rect 165669 -173933 165725 -173889
rect 165769 -173933 165825 -173889
rect 165869 -173933 165925 -173889
rect 165969 -173933 166025 -173889
rect 166069 -173933 166125 -173889
rect 166169 -173933 166225 -173889
rect 166269 -173933 166325 -173889
rect 166369 -173933 166425 -173889
rect 166469 -173933 166525 -173889
rect 166569 -173933 166625 -173889
rect 166669 -173933 166725 -173889
rect 166769 -173933 166825 -173889
rect 166869 -173933 166925 -173889
rect 166969 -173933 167025 -173889
rect 167069 -173933 167525 -173889
rect 167569 -173933 167625 -173889
rect 167669 -173933 167725 -173889
rect 167769 -173933 167825 -173889
rect 167869 -173933 167925 -173889
rect 167969 -173933 168025 -173889
rect 168069 -173933 168125 -173889
rect 168169 -173933 168225 -173889
rect 168269 -173933 168325 -173889
rect 168369 -173933 168425 -173889
rect 168469 -173933 168525 -173889
rect 168569 -173933 168625 -173889
rect 168669 -173933 168725 -173889
rect 168769 -173933 168825 -173889
rect 168869 -173933 168925 -173889
rect 168969 -173933 169025 -173889
rect 169069 -173933 169525 -173889
rect 169569 -173933 169625 -173889
rect 169669 -173933 169725 -173889
rect 169769 -173933 169825 -173889
rect 169869 -173933 169925 -173889
rect 169969 -173933 170025 -173889
rect 170069 -173933 170125 -173889
rect 170169 -173933 170225 -173889
rect 170269 -173933 170325 -173889
rect 170369 -173933 170425 -173889
rect 170469 -173933 170525 -173889
rect 170569 -173933 170625 -173889
rect 170669 -173933 170725 -173889
rect 170769 -173933 170825 -173889
rect 170869 -173933 170925 -173889
rect 170969 -173933 171025 -173889
rect 171069 -173933 171525 -173889
rect 171569 -173933 171625 -173889
rect 171669 -173933 171725 -173889
rect 171769 -173933 171825 -173889
rect 171869 -173933 171925 -173889
rect 171969 -173933 172025 -173889
rect 172069 -173933 172125 -173889
rect 172169 -173933 172225 -173889
rect 172269 -173933 172325 -173889
rect 172369 -173933 172425 -173889
rect 172469 -173933 172525 -173889
rect 172569 -173933 172625 -173889
rect 172669 -173933 172725 -173889
rect 172769 -173933 172825 -173889
rect 172869 -173933 172925 -173889
rect 172969 -173933 173025 -173889
rect 173069 -173933 178472 -173889
rect -114442 -173949 178472 -173933
rect -114442 -173993 81627 -173949
rect 81671 -173993 81727 -173949
rect 81771 -173993 81827 -173949
rect 81871 -173993 81927 -173949
rect 81971 -173993 82027 -173949
rect 82071 -173993 82127 -173949
rect 82171 -173993 82227 -173949
rect 82271 -173993 82327 -173949
rect 82371 -173993 82427 -173949
rect 82471 -173993 82527 -173949
rect 82571 -173993 82627 -173949
rect 82671 -173993 82727 -173949
rect 82771 -173993 82827 -173949
rect 82871 -173993 82927 -173949
rect 82971 -173993 83027 -173949
rect 83071 -173993 83127 -173949
rect 83171 -173993 83627 -173949
rect 83671 -173993 83727 -173949
rect 83771 -173993 83827 -173949
rect 83871 -173993 83927 -173949
rect 83971 -173993 84027 -173949
rect 84071 -173993 84127 -173949
rect 84171 -173993 84227 -173949
rect 84271 -173993 84327 -173949
rect 84371 -173993 84427 -173949
rect 84471 -173993 84527 -173949
rect 84571 -173993 84627 -173949
rect 84671 -173993 84727 -173949
rect 84771 -173993 84827 -173949
rect 84871 -173993 84927 -173949
rect 84971 -173993 85027 -173949
rect 85071 -173993 85127 -173949
rect 85171 -173993 85627 -173949
rect 85671 -173993 85727 -173949
rect 85771 -173993 85827 -173949
rect 85871 -173993 85927 -173949
rect 85971 -173993 86027 -173949
rect 86071 -173993 86127 -173949
rect 86171 -173993 86227 -173949
rect 86271 -173993 86327 -173949
rect 86371 -173993 86427 -173949
rect 86471 -173993 86527 -173949
rect 86571 -173993 86627 -173949
rect 86671 -173993 86727 -173949
rect 86771 -173993 86827 -173949
rect 86871 -173993 86927 -173949
rect 86971 -173993 87027 -173949
rect 87071 -173993 87127 -173949
rect 87171 -173993 87627 -173949
rect 87671 -173993 87727 -173949
rect 87771 -173993 87827 -173949
rect 87871 -173993 87927 -173949
rect 87971 -173993 88027 -173949
rect 88071 -173993 88127 -173949
rect 88171 -173993 88227 -173949
rect 88271 -173993 88327 -173949
rect 88371 -173993 88427 -173949
rect 88471 -173993 88527 -173949
rect 88571 -173993 88627 -173949
rect 88671 -173993 88727 -173949
rect 88771 -173993 88827 -173949
rect 88871 -173993 88927 -173949
rect 88971 -173993 89027 -173949
rect 89071 -173993 89127 -173949
rect 89171 -173989 178472 -173949
rect 89171 -173993 165525 -173989
rect -114442 -174033 165525 -173993
rect 165569 -174033 165625 -173989
rect 165669 -174033 165725 -173989
rect 165769 -174033 165825 -173989
rect 165869 -174033 165925 -173989
rect 165969 -174033 166025 -173989
rect 166069 -174033 166125 -173989
rect 166169 -174033 166225 -173989
rect 166269 -174033 166325 -173989
rect 166369 -174033 166425 -173989
rect 166469 -174033 166525 -173989
rect 166569 -174033 166625 -173989
rect 166669 -174033 166725 -173989
rect 166769 -174033 166825 -173989
rect 166869 -174033 166925 -173989
rect 166969 -174033 167025 -173989
rect 167069 -174033 167525 -173989
rect 167569 -174033 167625 -173989
rect 167669 -174033 167725 -173989
rect 167769 -174033 167825 -173989
rect 167869 -174033 167925 -173989
rect 167969 -174033 168025 -173989
rect 168069 -174033 168125 -173989
rect 168169 -174033 168225 -173989
rect 168269 -174033 168325 -173989
rect 168369 -174033 168425 -173989
rect 168469 -174033 168525 -173989
rect 168569 -174033 168625 -173989
rect 168669 -174033 168725 -173989
rect 168769 -174033 168825 -173989
rect 168869 -174033 168925 -173989
rect 168969 -174033 169025 -173989
rect 169069 -174033 169525 -173989
rect 169569 -174033 169625 -173989
rect 169669 -174033 169725 -173989
rect 169769 -174033 169825 -173989
rect 169869 -174033 169925 -173989
rect 169969 -174033 170025 -173989
rect 170069 -174033 170125 -173989
rect 170169 -174033 170225 -173989
rect 170269 -174033 170325 -173989
rect 170369 -174033 170425 -173989
rect 170469 -174033 170525 -173989
rect 170569 -174033 170625 -173989
rect 170669 -174033 170725 -173989
rect 170769 -174033 170825 -173989
rect 170869 -174033 170925 -173989
rect 170969 -174033 171025 -173989
rect 171069 -174033 171525 -173989
rect 171569 -174033 171625 -173989
rect 171669 -174033 171725 -173989
rect 171769 -174033 171825 -173989
rect 171869 -174033 171925 -173989
rect 171969 -174033 172025 -173989
rect 172069 -174033 172125 -173989
rect 172169 -174033 172225 -173989
rect 172269 -174033 172325 -173989
rect 172369 -174033 172425 -173989
rect 172469 -174033 172525 -173989
rect 172569 -174033 172625 -173989
rect 172669 -174033 172725 -173989
rect 172769 -174033 172825 -173989
rect 172869 -174033 172925 -173989
rect 172969 -174033 173025 -173989
rect 173069 -174033 178472 -173989
rect -114442 -174049 178472 -174033
rect -114442 -174093 81627 -174049
rect 81671 -174093 81727 -174049
rect 81771 -174093 81827 -174049
rect 81871 -174093 81927 -174049
rect 81971 -174093 82027 -174049
rect 82071 -174093 82127 -174049
rect 82171 -174093 82227 -174049
rect 82271 -174093 82327 -174049
rect 82371 -174093 82427 -174049
rect 82471 -174093 82527 -174049
rect 82571 -174093 82627 -174049
rect 82671 -174093 82727 -174049
rect 82771 -174093 82827 -174049
rect 82871 -174093 82927 -174049
rect 82971 -174093 83027 -174049
rect 83071 -174093 83127 -174049
rect 83171 -174093 83627 -174049
rect 83671 -174093 83727 -174049
rect 83771 -174093 83827 -174049
rect 83871 -174093 83927 -174049
rect 83971 -174093 84027 -174049
rect 84071 -174093 84127 -174049
rect 84171 -174093 84227 -174049
rect 84271 -174093 84327 -174049
rect 84371 -174093 84427 -174049
rect 84471 -174093 84527 -174049
rect 84571 -174093 84627 -174049
rect 84671 -174093 84727 -174049
rect 84771 -174093 84827 -174049
rect 84871 -174093 84927 -174049
rect 84971 -174093 85027 -174049
rect 85071 -174093 85127 -174049
rect 85171 -174093 85627 -174049
rect 85671 -174093 85727 -174049
rect 85771 -174093 85827 -174049
rect 85871 -174093 85927 -174049
rect 85971 -174093 86027 -174049
rect 86071 -174093 86127 -174049
rect 86171 -174093 86227 -174049
rect 86271 -174093 86327 -174049
rect 86371 -174093 86427 -174049
rect 86471 -174093 86527 -174049
rect 86571 -174093 86627 -174049
rect 86671 -174093 86727 -174049
rect 86771 -174093 86827 -174049
rect 86871 -174093 86927 -174049
rect 86971 -174093 87027 -174049
rect 87071 -174093 87127 -174049
rect 87171 -174093 87627 -174049
rect 87671 -174093 87727 -174049
rect 87771 -174093 87827 -174049
rect 87871 -174093 87927 -174049
rect 87971 -174093 88027 -174049
rect 88071 -174093 88127 -174049
rect 88171 -174093 88227 -174049
rect 88271 -174093 88327 -174049
rect 88371 -174093 88427 -174049
rect 88471 -174093 88527 -174049
rect 88571 -174093 88627 -174049
rect 88671 -174093 88727 -174049
rect 88771 -174093 88827 -174049
rect 88871 -174093 88927 -174049
rect 88971 -174093 89027 -174049
rect 89071 -174093 89127 -174049
rect 89171 -174089 178472 -174049
rect 89171 -174093 165525 -174089
rect -114442 -174133 165525 -174093
rect 165569 -174133 165625 -174089
rect 165669 -174133 165725 -174089
rect 165769 -174133 165825 -174089
rect 165869 -174133 165925 -174089
rect 165969 -174133 166025 -174089
rect 166069 -174133 166125 -174089
rect 166169 -174133 166225 -174089
rect 166269 -174133 166325 -174089
rect 166369 -174133 166425 -174089
rect 166469 -174133 166525 -174089
rect 166569 -174133 166625 -174089
rect 166669 -174133 166725 -174089
rect 166769 -174133 166825 -174089
rect 166869 -174133 166925 -174089
rect 166969 -174133 167025 -174089
rect 167069 -174133 167525 -174089
rect 167569 -174133 167625 -174089
rect 167669 -174133 167725 -174089
rect 167769 -174133 167825 -174089
rect 167869 -174133 167925 -174089
rect 167969 -174133 168025 -174089
rect 168069 -174133 168125 -174089
rect 168169 -174133 168225 -174089
rect 168269 -174133 168325 -174089
rect 168369 -174133 168425 -174089
rect 168469 -174133 168525 -174089
rect 168569 -174133 168625 -174089
rect 168669 -174133 168725 -174089
rect 168769 -174133 168825 -174089
rect 168869 -174133 168925 -174089
rect 168969 -174133 169025 -174089
rect 169069 -174133 169525 -174089
rect 169569 -174133 169625 -174089
rect 169669 -174133 169725 -174089
rect 169769 -174133 169825 -174089
rect 169869 -174133 169925 -174089
rect 169969 -174133 170025 -174089
rect 170069 -174133 170125 -174089
rect 170169 -174133 170225 -174089
rect 170269 -174133 170325 -174089
rect 170369 -174133 170425 -174089
rect 170469 -174133 170525 -174089
rect 170569 -174133 170625 -174089
rect 170669 -174133 170725 -174089
rect 170769 -174133 170825 -174089
rect 170869 -174133 170925 -174089
rect 170969 -174133 171025 -174089
rect 171069 -174133 171525 -174089
rect 171569 -174133 171625 -174089
rect 171669 -174133 171725 -174089
rect 171769 -174133 171825 -174089
rect 171869 -174133 171925 -174089
rect 171969 -174133 172025 -174089
rect 172069 -174133 172125 -174089
rect 172169 -174133 172225 -174089
rect 172269 -174133 172325 -174089
rect 172369 -174133 172425 -174089
rect 172469 -174133 172525 -174089
rect 172569 -174133 172625 -174089
rect 172669 -174133 172725 -174089
rect 172769 -174133 172825 -174089
rect 172869 -174133 172925 -174089
rect 172969 -174133 173025 -174089
rect 173069 -174133 178472 -174089
rect -114442 -174149 178472 -174133
rect -114442 -174193 81627 -174149
rect 81671 -174193 81727 -174149
rect 81771 -174193 81827 -174149
rect 81871 -174193 81927 -174149
rect 81971 -174193 82027 -174149
rect 82071 -174193 82127 -174149
rect 82171 -174193 82227 -174149
rect 82271 -174193 82327 -174149
rect 82371 -174193 82427 -174149
rect 82471 -174193 82527 -174149
rect 82571 -174193 82627 -174149
rect 82671 -174193 82727 -174149
rect 82771 -174193 82827 -174149
rect 82871 -174193 82927 -174149
rect 82971 -174193 83027 -174149
rect 83071 -174193 83127 -174149
rect 83171 -174193 83627 -174149
rect 83671 -174193 83727 -174149
rect 83771 -174193 83827 -174149
rect 83871 -174193 83927 -174149
rect 83971 -174193 84027 -174149
rect 84071 -174193 84127 -174149
rect 84171 -174193 84227 -174149
rect 84271 -174193 84327 -174149
rect 84371 -174193 84427 -174149
rect 84471 -174193 84527 -174149
rect 84571 -174193 84627 -174149
rect 84671 -174193 84727 -174149
rect 84771 -174193 84827 -174149
rect 84871 -174193 84927 -174149
rect 84971 -174193 85027 -174149
rect 85071 -174193 85127 -174149
rect 85171 -174193 85627 -174149
rect 85671 -174193 85727 -174149
rect 85771 -174193 85827 -174149
rect 85871 -174193 85927 -174149
rect 85971 -174193 86027 -174149
rect 86071 -174193 86127 -174149
rect 86171 -174193 86227 -174149
rect 86271 -174193 86327 -174149
rect 86371 -174193 86427 -174149
rect 86471 -174193 86527 -174149
rect 86571 -174193 86627 -174149
rect 86671 -174193 86727 -174149
rect 86771 -174193 86827 -174149
rect 86871 -174193 86927 -174149
rect 86971 -174193 87027 -174149
rect 87071 -174193 87127 -174149
rect 87171 -174193 87627 -174149
rect 87671 -174193 87727 -174149
rect 87771 -174193 87827 -174149
rect 87871 -174193 87927 -174149
rect 87971 -174193 88027 -174149
rect 88071 -174193 88127 -174149
rect 88171 -174193 88227 -174149
rect 88271 -174193 88327 -174149
rect 88371 -174193 88427 -174149
rect 88471 -174193 88527 -174149
rect 88571 -174193 88627 -174149
rect 88671 -174193 88727 -174149
rect 88771 -174193 88827 -174149
rect 88871 -174193 88927 -174149
rect 88971 -174193 89027 -174149
rect 89071 -174193 89127 -174149
rect 89171 -174189 178472 -174149
rect 89171 -174193 165525 -174189
rect -114442 -174233 165525 -174193
rect 165569 -174233 165625 -174189
rect 165669 -174233 165725 -174189
rect 165769 -174233 165825 -174189
rect 165869 -174233 165925 -174189
rect 165969 -174233 166025 -174189
rect 166069 -174233 166125 -174189
rect 166169 -174233 166225 -174189
rect 166269 -174233 166325 -174189
rect 166369 -174233 166425 -174189
rect 166469 -174233 166525 -174189
rect 166569 -174233 166625 -174189
rect 166669 -174233 166725 -174189
rect 166769 -174233 166825 -174189
rect 166869 -174233 166925 -174189
rect 166969 -174233 167025 -174189
rect 167069 -174233 167525 -174189
rect 167569 -174233 167625 -174189
rect 167669 -174233 167725 -174189
rect 167769 -174233 167825 -174189
rect 167869 -174233 167925 -174189
rect 167969 -174233 168025 -174189
rect 168069 -174233 168125 -174189
rect 168169 -174233 168225 -174189
rect 168269 -174233 168325 -174189
rect 168369 -174233 168425 -174189
rect 168469 -174233 168525 -174189
rect 168569 -174233 168625 -174189
rect 168669 -174233 168725 -174189
rect 168769 -174233 168825 -174189
rect 168869 -174233 168925 -174189
rect 168969 -174233 169025 -174189
rect 169069 -174233 169525 -174189
rect 169569 -174233 169625 -174189
rect 169669 -174233 169725 -174189
rect 169769 -174233 169825 -174189
rect 169869 -174233 169925 -174189
rect 169969 -174233 170025 -174189
rect 170069 -174233 170125 -174189
rect 170169 -174233 170225 -174189
rect 170269 -174233 170325 -174189
rect 170369 -174233 170425 -174189
rect 170469 -174233 170525 -174189
rect 170569 -174233 170625 -174189
rect 170669 -174233 170725 -174189
rect 170769 -174233 170825 -174189
rect 170869 -174233 170925 -174189
rect 170969 -174233 171025 -174189
rect 171069 -174233 171525 -174189
rect 171569 -174233 171625 -174189
rect 171669 -174233 171725 -174189
rect 171769 -174233 171825 -174189
rect 171869 -174233 171925 -174189
rect 171969 -174233 172025 -174189
rect 172069 -174233 172125 -174189
rect 172169 -174233 172225 -174189
rect 172269 -174233 172325 -174189
rect 172369 -174233 172425 -174189
rect 172469 -174233 172525 -174189
rect 172569 -174233 172625 -174189
rect 172669 -174233 172725 -174189
rect 172769 -174233 172825 -174189
rect 172869 -174233 172925 -174189
rect 172969 -174233 173025 -174189
rect 173069 -174233 178472 -174189
rect -114442 -174249 178472 -174233
rect -114442 -174293 81627 -174249
rect 81671 -174293 81727 -174249
rect 81771 -174293 81827 -174249
rect 81871 -174293 81927 -174249
rect 81971 -174293 82027 -174249
rect 82071 -174293 82127 -174249
rect 82171 -174293 82227 -174249
rect 82271 -174293 82327 -174249
rect 82371 -174293 82427 -174249
rect 82471 -174293 82527 -174249
rect 82571 -174293 82627 -174249
rect 82671 -174293 82727 -174249
rect 82771 -174293 82827 -174249
rect 82871 -174293 82927 -174249
rect 82971 -174293 83027 -174249
rect 83071 -174293 83127 -174249
rect 83171 -174293 83627 -174249
rect 83671 -174293 83727 -174249
rect 83771 -174293 83827 -174249
rect 83871 -174293 83927 -174249
rect 83971 -174293 84027 -174249
rect 84071 -174293 84127 -174249
rect 84171 -174293 84227 -174249
rect 84271 -174293 84327 -174249
rect 84371 -174293 84427 -174249
rect 84471 -174293 84527 -174249
rect 84571 -174293 84627 -174249
rect 84671 -174293 84727 -174249
rect 84771 -174293 84827 -174249
rect 84871 -174293 84927 -174249
rect 84971 -174293 85027 -174249
rect 85071 -174293 85127 -174249
rect 85171 -174293 85627 -174249
rect 85671 -174293 85727 -174249
rect 85771 -174293 85827 -174249
rect 85871 -174293 85927 -174249
rect 85971 -174293 86027 -174249
rect 86071 -174293 86127 -174249
rect 86171 -174293 86227 -174249
rect 86271 -174293 86327 -174249
rect 86371 -174293 86427 -174249
rect 86471 -174293 86527 -174249
rect 86571 -174293 86627 -174249
rect 86671 -174293 86727 -174249
rect 86771 -174293 86827 -174249
rect 86871 -174293 86927 -174249
rect 86971 -174293 87027 -174249
rect 87071 -174293 87127 -174249
rect 87171 -174293 87627 -174249
rect 87671 -174293 87727 -174249
rect 87771 -174293 87827 -174249
rect 87871 -174293 87927 -174249
rect 87971 -174293 88027 -174249
rect 88071 -174293 88127 -174249
rect 88171 -174293 88227 -174249
rect 88271 -174293 88327 -174249
rect 88371 -174293 88427 -174249
rect 88471 -174293 88527 -174249
rect 88571 -174293 88627 -174249
rect 88671 -174293 88727 -174249
rect 88771 -174293 88827 -174249
rect 88871 -174293 88927 -174249
rect 88971 -174293 89027 -174249
rect 89071 -174293 89127 -174249
rect 89171 -174289 178472 -174249
rect 89171 -174293 165525 -174289
rect -114442 -174333 165525 -174293
rect 165569 -174333 165625 -174289
rect 165669 -174333 165725 -174289
rect 165769 -174333 165825 -174289
rect 165869 -174333 165925 -174289
rect 165969 -174333 166025 -174289
rect 166069 -174333 166125 -174289
rect 166169 -174333 166225 -174289
rect 166269 -174333 166325 -174289
rect 166369 -174333 166425 -174289
rect 166469 -174333 166525 -174289
rect 166569 -174333 166625 -174289
rect 166669 -174333 166725 -174289
rect 166769 -174333 166825 -174289
rect 166869 -174333 166925 -174289
rect 166969 -174333 167025 -174289
rect 167069 -174333 167525 -174289
rect 167569 -174333 167625 -174289
rect 167669 -174333 167725 -174289
rect 167769 -174333 167825 -174289
rect 167869 -174333 167925 -174289
rect 167969 -174333 168025 -174289
rect 168069 -174333 168125 -174289
rect 168169 -174333 168225 -174289
rect 168269 -174333 168325 -174289
rect 168369 -174333 168425 -174289
rect 168469 -174333 168525 -174289
rect 168569 -174333 168625 -174289
rect 168669 -174333 168725 -174289
rect 168769 -174333 168825 -174289
rect 168869 -174333 168925 -174289
rect 168969 -174333 169025 -174289
rect 169069 -174333 169525 -174289
rect 169569 -174333 169625 -174289
rect 169669 -174333 169725 -174289
rect 169769 -174333 169825 -174289
rect 169869 -174333 169925 -174289
rect 169969 -174333 170025 -174289
rect 170069 -174333 170125 -174289
rect 170169 -174333 170225 -174289
rect 170269 -174333 170325 -174289
rect 170369 -174333 170425 -174289
rect 170469 -174333 170525 -174289
rect 170569 -174333 170625 -174289
rect 170669 -174333 170725 -174289
rect 170769 -174333 170825 -174289
rect 170869 -174333 170925 -174289
rect 170969 -174333 171025 -174289
rect 171069 -174333 171525 -174289
rect 171569 -174333 171625 -174289
rect 171669 -174333 171725 -174289
rect 171769 -174333 171825 -174289
rect 171869 -174333 171925 -174289
rect 171969 -174333 172025 -174289
rect 172069 -174333 172125 -174289
rect 172169 -174333 172225 -174289
rect 172269 -174333 172325 -174289
rect 172369 -174333 172425 -174289
rect 172469 -174333 172525 -174289
rect 172569 -174333 172625 -174289
rect 172669 -174333 172725 -174289
rect 172769 -174333 172825 -174289
rect 172869 -174333 172925 -174289
rect 172969 -174333 173025 -174289
rect 173069 -174333 178472 -174289
rect -114442 -174349 178472 -174333
rect -114442 -174393 81627 -174349
rect 81671 -174393 81727 -174349
rect 81771 -174393 81827 -174349
rect 81871 -174393 81927 -174349
rect 81971 -174393 82027 -174349
rect 82071 -174393 82127 -174349
rect 82171 -174393 82227 -174349
rect 82271 -174393 82327 -174349
rect 82371 -174393 82427 -174349
rect 82471 -174393 82527 -174349
rect 82571 -174393 82627 -174349
rect 82671 -174393 82727 -174349
rect 82771 -174393 82827 -174349
rect 82871 -174393 82927 -174349
rect 82971 -174393 83027 -174349
rect 83071 -174393 83127 -174349
rect 83171 -174393 83627 -174349
rect 83671 -174393 83727 -174349
rect 83771 -174393 83827 -174349
rect 83871 -174393 83927 -174349
rect 83971 -174393 84027 -174349
rect 84071 -174393 84127 -174349
rect 84171 -174393 84227 -174349
rect 84271 -174393 84327 -174349
rect 84371 -174393 84427 -174349
rect 84471 -174393 84527 -174349
rect 84571 -174393 84627 -174349
rect 84671 -174393 84727 -174349
rect 84771 -174393 84827 -174349
rect 84871 -174393 84927 -174349
rect 84971 -174393 85027 -174349
rect 85071 -174393 85127 -174349
rect 85171 -174393 85627 -174349
rect 85671 -174393 85727 -174349
rect 85771 -174393 85827 -174349
rect 85871 -174393 85927 -174349
rect 85971 -174393 86027 -174349
rect 86071 -174393 86127 -174349
rect 86171 -174393 86227 -174349
rect 86271 -174393 86327 -174349
rect 86371 -174393 86427 -174349
rect 86471 -174393 86527 -174349
rect 86571 -174393 86627 -174349
rect 86671 -174393 86727 -174349
rect 86771 -174393 86827 -174349
rect 86871 -174393 86927 -174349
rect 86971 -174393 87027 -174349
rect 87071 -174393 87127 -174349
rect 87171 -174393 87627 -174349
rect 87671 -174393 87727 -174349
rect 87771 -174393 87827 -174349
rect 87871 -174393 87927 -174349
rect 87971 -174393 88027 -174349
rect 88071 -174393 88127 -174349
rect 88171 -174393 88227 -174349
rect 88271 -174393 88327 -174349
rect 88371 -174393 88427 -174349
rect 88471 -174393 88527 -174349
rect 88571 -174393 88627 -174349
rect 88671 -174393 88727 -174349
rect 88771 -174393 88827 -174349
rect 88871 -174393 88927 -174349
rect 88971 -174393 89027 -174349
rect 89071 -174393 89127 -174349
rect 89171 -174389 178472 -174349
rect 89171 -174393 165525 -174389
rect -114442 -174433 165525 -174393
rect 165569 -174433 165625 -174389
rect 165669 -174433 165725 -174389
rect 165769 -174433 165825 -174389
rect 165869 -174433 165925 -174389
rect 165969 -174433 166025 -174389
rect 166069 -174433 166125 -174389
rect 166169 -174433 166225 -174389
rect 166269 -174433 166325 -174389
rect 166369 -174433 166425 -174389
rect 166469 -174433 166525 -174389
rect 166569 -174433 166625 -174389
rect 166669 -174433 166725 -174389
rect 166769 -174433 166825 -174389
rect 166869 -174433 166925 -174389
rect 166969 -174433 167025 -174389
rect 167069 -174433 167525 -174389
rect 167569 -174433 167625 -174389
rect 167669 -174433 167725 -174389
rect 167769 -174433 167825 -174389
rect 167869 -174433 167925 -174389
rect 167969 -174433 168025 -174389
rect 168069 -174433 168125 -174389
rect 168169 -174433 168225 -174389
rect 168269 -174433 168325 -174389
rect 168369 -174433 168425 -174389
rect 168469 -174433 168525 -174389
rect 168569 -174433 168625 -174389
rect 168669 -174433 168725 -174389
rect 168769 -174433 168825 -174389
rect 168869 -174433 168925 -174389
rect 168969 -174433 169025 -174389
rect 169069 -174433 169525 -174389
rect 169569 -174433 169625 -174389
rect 169669 -174433 169725 -174389
rect 169769 -174433 169825 -174389
rect 169869 -174433 169925 -174389
rect 169969 -174433 170025 -174389
rect 170069 -174433 170125 -174389
rect 170169 -174433 170225 -174389
rect 170269 -174433 170325 -174389
rect 170369 -174433 170425 -174389
rect 170469 -174433 170525 -174389
rect 170569 -174433 170625 -174389
rect 170669 -174433 170725 -174389
rect 170769 -174433 170825 -174389
rect 170869 -174433 170925 -174389
rect 170969 -174433 171025 -174389
rect 171069 -174433 171525 -174389
rect 171569 -174433 171625 -174389
rect 171669 -174433 171725 -174389
rect 171769 -174433 171825 -174389
rect 171869 -174433 171925 -174389
rect 171969 -174433 172025 -174389
rect 172069 -174433 172125 -174389
rect 172169 -174433 172225 -174389
rect 172269 -174433 172325 -174389
rect 172369 -174433 172425 -174389
rect 172469 -174433 172525 -174389
rect 172569 -174433 172625 -174389
rect 172669 -174433 172725 -174389
rect 172769 -174433 172825 -174389
rect 172869 -174433 172925 -174389
rect 172969 -174433 173025 -174389
rect 173069 -174433 178472 -174389
rect -114442 -174449 178472 -174433
rect -114442 -174493 81627 -174449
rect 81671 -174493 81727 -174449
rect 81771 -174493 81827 -174449
rect 81871 -174493 81927 -174449
rect 81971 -174493 82027 -174449
rect 82071 -174493 82127 -174449
rect 82171 -174493 82227 -174449
rect 82271 -174493 82327 -174449
rect 82371 -174493 82427 -174449
rect 82471 -174493 82527 -174449
rect 82571 -174493 82627 -174449
rect 82671 -174493 82727 -174449
rect 82771 -174493 82827 -174449
rect 82871 -174493 82927 -174449
rect 82971 -174493 83027 -174449
rect 83071 -174493 83127 -174449
rect 83171 -174493 83627 -174449
rect 83671 -174493 83727 -174449
rect 83771 -174493 83827 -174449
rect 83871 -174493 83927 -174449
rect 83971 -174493 84027 -174449
rect 84071 -174493 84127 -174449
rect 84171 -174493 84227 -174449
rect 84271 -174493 84327 -174449
rect 84371 -174493 84427 -174449
rect 84471 -174493 84527 -174449
rect 84571 -174493 84627 -174449
rect 84671 -174493 84727 -174449
rect 84771 -174493 84827 -174449
rect 84871 -174493 84927 -174449
rect 84971 -174493 85027 -174449
rect 85071 -174493 85127 -174449
rect 85171 -174493 85627 -174449
rect 85671 -174493 85727 -174449
rect 85771 -174493 85827 -174449
rect 85871 -174493 85927 -174449
rect 85971 -174493 86027 -174449
rect 86071 -174493 86127 -174449
rect 86171 -174493 86227 -174449
rect 86271 -174493 86327 -174449
rect 86371 -174493 86427 -174449
rect 86471 -174493 86527 -174449
rect 86571 -174493 86627 -174449
rect 86671 -174493 86727 -174449
rect 86771 -174493 86827 -174449
rect 86871 -174493 86927 -174449
rect 86971 -174493 87027 -174449
rect 87071 -174493 87127 -174449
rect 87171 -174493 87627 -174449
rect 87671 -174493 87727 -174449
rect 87771 -174493 87827 -174449
rect 87871 -174493 87927 -174449
rect 87971 -174493 88027 -174449
rect 88071 -174493 88127 -174449
rect 88171 -174493 88227 -174449
rect 88271 -174493 88327 -174449
rect 88371 -174493 88427 -174449
rect 88471 -174493 88527 -174449
rect 88571 -174493 88627 -174449
rect 88671 -174493 88727 -174449
rect 88771 -174493 88827 -174449
rect 88871 -174493 88927 -174449
rect 88971 -174493 89027 -174449
rect 89071 -174493 89127 -174449
rect 89171 -174489 178472 -174449
rect 89171 -174493 165525 -174489
rect -114442 -174533 165525 -174493
rect 165569 -174533 165625 -174489
rect 165669 -174533 165725 -174489
rect 165769 -174533 165825 -174489
rect 165869 -174533 165925 -174489
rect 165969 -174533 166025 -174489
rect 166069 -174533 166125 -174489
rect 166169 -174533 166225 -174489
rect 166269 -174533 166325 -174489
rect 166369 -174533 166425 -174489
rect 166469 -174533 166525 -174489
rect 166569 -174533 166625 -174489
rect 166669 -174533 166725 -174489
rect 166769 -174533 166825 -174489
rect 166869 -174533 166925 -174489
rect 166969 -174533 167025 -174489
rect 167069 -174533 167525 -174489
rect 167569 -174533 167625 -174489
rect 167669 -174533 167725 -174489
rect 167769 -174533 167825 -174489
rect 167869 -174533 167925 -174489
rect 167969 -174533 168025 -174489
rect 168069 -174533 168125 -174489
rect 168169 -174533 168225 -174489
rect 168269 -174533 168325 -174489
rect 168369 -174533 168425 -174489
rect 168469 -174533 168525 -174489
rect 168569 -174533 168625 -174489
rect 168669 -174533 168725 -174489
rect 168769 -174533 168825 -174489
rect 168869 -174533 168925 -174489
rect 168969 -174533 169025 -174489
rect 169069 -174533 169525 -174489
rect 169569 -174533 169625 -174489
rect 169669 -174533 169725 -174489
rect 169769 -174533 169825 -174489
rect 169869 -174533 169925 -174489
rect 169969 -174533 170025 -174489
rect 170069 -174533 170125 -174489
rect 170169 -174533 170225 -174489
rect 170269 -174533 170325 -174489
rect 170369 -174533 170425 -174489
rect 170469 -174533 170525 -174489
rect 170569 -174533 170625 -174489
rect 170669 -174533 170725 -174489
rect 170769 -174533 170825 -174489
rect 170869 -174533 170925 -174489
rect 170969 -174533 171025 -174489
rect 171069 -174533 171525 -174489
rect 171569 -174533 171625 -174489
rect 171669 -174533 171725 -174489
rect 171769 -174533 171825 -174489
rect 171869 -174533 171925 -174489
rect 171969 -174533 172025 -174489
rect 172069 -174533 172125 -174489
rect 172169 -174533 172225 -174489
rect 172269 -174533 172325 -174489
rect 172369 -174533 172425 -174489
rect 172469 -174533 172525 -174489
rect 172569 -174533 172625 -174489
rect 172669 -174533 172725 -174489
rect 172769 -174533 172825 -174489
rect 172869 -174533 172925 -174489
rect 172969 -174533 173025 -174489
rect 173069 -174533 178472 -174489
rect -114442 -174549 178472 -174533
rect -114442 -174593 81627 -174549
rect 81671 -174593 81727 -174549
rect 81771 -174593 81827 -174549
rect 81871 -174593 81927 -174549
rect 81971 -174593 82027 -174549
rect 82071 -174593 82127 -174549
rect 82171 -174593 82227 -174549
rect 82271 -174593 82327 -174549
rect 82371 -174593 82427 -174549
rect 82471 -174593 82527 -174549
rect 82571 -174593 82627 -174549
rect 82671 -174593 82727 -174549
rect 82771 -174593 82827 -174549
rect 82871 -174593 82927 -174549
rect 82971 -174593 83027 -174549
rect 83071 -174593 83127 -174549
rect 83171 -174593 83627 -174549
rect 83671 -174593 83727 -174549
rect 83771 -174593 83827 -174549
rect 83871 -174593 83927 -174549
rect 83971 -174593 84027 -174549
rect 84071 -174593 84127 -174549
rect 84171 -174593 84227 -174549
rect 84271 -174593 84327 -174549
rect 84371 -174593 84427 -174549
rect 84471 -174593 84527 -174549
rect 84571 -174593 84627 -174549
rect 84671 -174593 84727 -174549
rect 84771 -174593 84827 -174549
rect 84871 -174593 84927 -174549
rect 84971 -174593 85027 -174549
rect 85071 -174593 85127 -174549
rect 85171 -174593 85627 -174549
rect 85671 -174593 85727 -174549
rect 85771 -174593 85827 -174549
rect 85871 -174593 85927 -174549
rect 85971 -174593 86027 -174549
rect 86071 -174593 86127 -174549
rect 86171 -174593 86227 -174549
rect 86271 -174593 86327 -174549
rect 86371 -174593 86427 -174549
rect 86471 -174593 86527 -174549
rect 86571 -174593 86627 -174549
rect 86671 -174593 86727 -174549
rect 86771 -174593 86827 -174549
rect 86871 -174593 86927 -174549
rect 86971 -174593 87027 -174549
rect 87071 -174593 87127 -174549
rect 87171 -174593 87627 -174549
rect 87671 -174593 87727 -174549
rect 87771 -174593 87827 -174549
rect 87871 -174593 87927 -174549
rect 87971 -174593 88027 -174549
rect 88071 -174593 88127 -174549
rect 88171 -174593 88227 -174549
rect 88271 -174593 88327 -174549
rect 88371 -174593 88427 -174549
rect 88471 -174593 88527 -174549
rect 88571 -174593 88627 -174549
rect 88671 -174593 88727 -174549
rect 88771 -174593 88827 -174549
rect 88871 -174593 88927 -174549
rect 88971 -174593 89027 -174549
rect 89071 -174593 89127 -174549
rect 89171 -174593 178472 -174549
rect -114442 -176471 178472 -174593
<< via1 >>
rect -27407 3511 -27363 3555
rect -27307 3511 -27263 3555
rect -27207 3511 -27163 3555
rect -27107 3511 -27063 3555
rect -27007 3511 -26963 3555
rect -26907 3511 -26863 3555
rect -26807 3511 -26763 3555
rect -26707 3511 -26663 3555
rect -26607 3511 -26563 3555
rect -26507 3511 -26463 3555
rect -26407 3511 -26363 3555
rect -26307 3511 -26263 3555
rect -26207 3511 -26163 3555
rect -26107 3511 -26063 3555
rect -26007 3511 -25963 3555
rect -25907 3511 -25863 3555
rect -25407 3511 -25363 3555
rect -25307 3511 -25263 3555
rect -25207 3511 -25163 3555
rect -25107 3511 -25063 3555
rect -25007 3511 -24963 3555
rect -24907 3511 -24863 3555
rect -24807 3511 -24763 3555
rect -24707 3511 -24663 3555
rect -24607 3511 -24563 3555
rect -24507 3511 -24463 3555
rect -24407 3511 -24363 3555
rect -24307 3511 -24263 3555
rect -24207 3511 -24163 3555
rect -24107 3511 -24063 3555
rect -24007 3511 -23963 3555
rect -23907 3511 -23863 3555
rect -23407 3511 -23363 3555
rect -23307 3511 -23263 3555
rect -23207 3511 -23163 3555
rect -23107 3511 -23063 3555
rect -23007 3511 -22963 3555
rect -22907 3511 -22863 3555
rect -22807 3511 -22763 3555
rect -22707 3511 -22663 3555
rect -22607 3511 -22563 3555
rect -22507 3511 -22463 3555
rect -22407 3511 -22363 3555
rect -22307 3511 -22263 3555
rect -22207 3511 -22163 3555
rect -22107 3511 -22063 3555
rect -22007 3511 -21963 3555
rect -21907 3511 -21863 3555
rect -21407 3511 -21363 3555
rect -21307 3511 -21263 3555
rect -21207 3511 -21163 3555
rect -21107 3511 -21063 3555
rect -21007 3511 -20963 3555
rect -20907 3511 -20863 3555
rect -20807 3511 -20763 3555
rect -20707 3511 -20663 3555
rect -20607 3511 -20563 3555
rect -20507 3511 -20463 3555
rect -20407 3511 -20363 3555
rect -20307 3511 -20263 3555
rect -20207 3511 -20163 3555
rect -20107 3511 -20063 3555
rect -20007 3511 -19963 3555
rect -19907 3511 -19863 3555
rect -27407 3411 -27363 3455
rect -27307 3411 -27263 3455
rect -27207 3411 -27163 3455
rect -27107 3411 -27063 3455
rect -27007 3411 -26963 3455
rect -26907 3411 -26863 3455
rect -26807 3411 -26763 3455
rect -26707 3411 -26663 3455
rect -26607 3411 -26563 3455
rect -26507 3411 -26463 3455
rect -26407 3411 -26363 3455
rect -26307 3411 -26263 3455
rect -26207 3411 -26163 3455
rect -26107 3411 -26063 3455
rect -26007 3411 -25963 3455
rect -25907 3411 -25863 3455
rect -25407 3411 -25363 3455
rect -25307 3411 -25263 3455
rect -25207 3411 -25163 3455
rect -25107 3411 -25063 3455
rect -25007 3411 -24963 3455
rect -24907 3411 -24863 3455
rect -24807 3411 -24763 3455
rect -24707 3411 -24663 3455
rect -24607 3411 -24563 3455
rect -24507 3411 -24463 3455
rect -24407 3411 -24363 3455
rect -24307 3411 -24263 3455
rect -24207 3411 -24163 3455
rect -24107 3411 -24063 3455
rect -24007 3411 -23963 3455
rect -23907 3411 -23863 3455
rect -23407 3411 -23363 3455
rect -23307 3411 -23263 3455
rect -23207 3411 -23163 3455
rect -23107 3411 -23063 3455
rect -23007 3411 -22963 3455
rect -22907 3411 -22863 3455
rect -22807 3411 -22763 3455
rect -22707 3411 -22663 3455
rect -22607 3411 -22563 3455
rect -22507 3411 -22463 3455
rect -22407 3411 -22363 3455
rect -22307 3411 -22263 3455
rect -22207 3411 -22163 3455
rect -22107 3411 -22063 3455
rect -22007 3411 -21963 3455
rect -21907 3411 -21863 3455
rect -21407 3411 -21363 3455
rect -21307 3411 -21263 3455
rect -21207 3411 -21163 3455
rect -21107 3411 -21063 3455
rect -21007 3411 -20963 3455
rect -20907 3411 -20863 3455
rect -20807 3411 -20763 3455
rect -20707 3411 -20663 3455
rect -20607 3411 -20563 3455
rect -20507 3411 -20463 3455
rect -20407 3411 -20363 3455
rect -20307 3411 -20263 3455
rect -20207 3411 -20163 3455
rect -20107 3411 -20063 3455
rect -20007 3411 -19963 3455
rect -19907 3411 -19863 3455
rect -27407 3311 -27363 3355
rect -27307 3311 -27263 3355
rect -27207 3311 -27163 3355
rect -27107 3311 -27063 3355
rect -27007 3311 -26963 3355
rect -26907 3311 -26863 3355
rect -26807 3311 -26763 3355
rect -26707 3311 -26663 3355
rect -26607 3311 -26563 3355
rect -26507 3311 -26463 3355
rect -26407 3311 -26363 3355
rect -26307 3311 -26263 3355
rect -26207 3311 -26163 3355
rect -26107 3311 -26063 3355
rect -26007 3311 -25963 3355
rect -25907 3311 -25863 3355
rect -25407 3311 -25363 3355
rect -25307 3311 -25263 3355
rect -25207 3311 -25163 3355
rect -25107 3311 -25063 3355
rect -25007 3311 -24963 3355
rect -24907 3311 -24863 3355
rect -24807 3311 -24763 3355
rect -24707 3311 -24663 3355
rect -24607 3311 -24563 3355
rect -24507 3311 -24463 3355
rect -24407 3311 -24363 3355
rect -24307 3311 -24263 3355
rect -24207 3311 -24163 3355
rect -24107 3311 -24063 3355
rect -24007 3311 -23963 3355
rect -23907 3311 -23863 3355
rect -23407 3311 -23363 3355
rect -23307 3311 -23263 3355
rect -23207 3311 -23163 3355
rect -23107 3311 -23063 3355
rect -23007 3311 -22963 3355
rect -22907 3311 -22863 3355
rect -22807 3311 -22763 3355
rect -22707 3311 -22663 3355
rect -22607 3311 -22563 3355
rect -22507 3311 -22463 3355
rect -22407 3311 -22363 3355
rect -22307 3311 -22263 3355
rect -22207 3311 -22163 3355
rect -22107 3311 -22063 3355
rect -22007 3311 -21963 3355
rect -21907 3311 -21863 3355
rect -21407 3311 -21363 3355
rect -21307 3311 -21263 3355
rect -21207 3311 -21163 3355
rect -21107 3311 -21063 3355
rect -21007 3311 -20963 3355
rect -20907 3311 -20863 3355
rect -20807 3311 -20763 3355
rect -20707 3311 -20663 3355
rect -20607 3311 -20563 3355
rect -20507 3311 -20463 3355
rect -20407 3311 -20363 3355
rect -20307 3311 -20263 3355
rect -20207 3311 -20163 3355
rect -20107 3311 -20063 3355
rect -20007 3311 -19963 3355
rect -19907 3311 -19863 3355
rect -27407 3211 -27363 3255
rect -27307 3211 -27263 3255
rect -27207 3211 -27163 3255
rect -27107 3211 -27063 3255
rect -27007 3211 -26963 3255
rect -26907 3211 -26863 3255
rect -26807 3211 -26763 3255
rect -26707 3211 -26663 3255
rect -26607 3211 -26563 3255
rect -26507 3211 -26463 3255
rect -26407 3211 -26363 3255
rect -26307 3211 -26263 3255
rect -26207 3211 -26163 3255
rect -26107 3211 -26063 3255
rect -26007 3211 -25963 3255
rect -25907 3211 -25863 3255
rect -25407 3211 -25363 3255
rect -25307 3211 -25263 3255
rect -25207 3211 -25163 3255
rect -25107 3211 -25063 3255
rect -25007 3211 -24963 3255
rect -24907 3211 -24863 3255
rect -24807 3211 -24763 3255
rect -24707 3211 -24663 3255
rect -24607 3211 -24563 3255
rect -24507 3211 -24463 3255
rect -24407 3211 -24363 3255
rect -24307 3211 -24263 3255
rect -24207 3211 -24163 3255
rect -24107 3211 -24063 3255
rect -24007 3211 -23963 3255
rect -23907 3211 -23863 3255
rect -23407 3211 -23363 3255
rect -23307 3211 -23263 3255
rect -23207 3211 -23163 3255
rect -23107 3211 -23063 3255
rect -23007 3211 -22963 3255
rect -22907 3211 -22863 3255
rect -22807 3211 -22763 3255
rect -22707 3211 -22663 3255
rect -22607 3211 -22563 3255
rect -22507 3211 -22463 3255
rect -22407 3211 -22363 3255
rect -22307 3211 -22263 3255
rect -22207 3211 -22163 3255
rect -22107 3211 -22063 3255
rect -22007 3211 -21963 3255
rect -21907 3211 -21863 3255
rect -21407 3211 -21363 3255
rect -21307 3211 -21263 3255
rect -21207 3211 -21163 3255
rect -21107 3211 -21063 3255
rect -21007 3211 -20963 3255
rect -20907 3211 -20863 3255
rect -20807 3211 -20763 3255
rect -20707 3211 -20663 3255
rect -20607 3211 -20563 3255
rect -20507 3211 -20463 3255
rect -20407 3211 -20363 3255
rect -20307 3211 -20263 3255
rect -20207 3211 -20163 3255
rect -20107 3211 -20063 3255
rect -20007 3211 -19963 3255
rect -19907 3211 -19863 3255
rect -27407 3111 -27363 3155
rect -27307 3111 -27263 3155
rect -27207 3111 -27163 3155
rect -27107 3111 -27063 3155
rect -27007 3111 -26963 3155
rect -26907 3111 -26863 3155
rect -26807 3111 -26763 3155
rect -26707 3111 -26663 3155
rect -26607 3111 -26563 3155
rect -26507 3111 -26463 3155
rect -26407 3111 -26363 3155
rect -26307 3111 -26263 3155
rect -26207 3111 -26163 3155
rect -26107 3111 -26063 3155
rect -26007 3111 -25963 3155
rect -25907 3111 -25863 3155
rect -25407 3111 -25363 3155
rect -25307 3111 -25263 3155
rect -25207 3111 -25163 3155
rect -25107 3111 -25063 3155
rect -25007 3111 -24963 3155
rect -24907 3111 -24863 3155
rect -24807 3111 -24763 3155
rect -24707 3111 -24663 3155
rect -24607 3111 -24563 3155
rect -24507 3111 -24463 3155
rect -24407 3111 -24363 3155
rect -24307 3111 -24263 3155
rect -24207 3111 -24163 3155
rect -24107 3111 -24063 3155
rect -24007 3111 -23963 3155
rect -23907 3111 -23863 3155
rect -23407 3111 -23363 3155
rect -23307 3111 -23263 3155
rect -23207 3111 -23163 3155
rect -23107 3111 -23063 3155
rect -23007 3111 -22963 3155
rect -22907 3111 -22863 3155
rect -22807 3111 -22763 3155
rect -22707 3111 -22663 3155
rect -22607 3111 -22563 3155
rect -22507 3111 -22463 3155
rect -22407 3111 -22363 3155
rect -22307 3111 -22263 3155
rect -22207 3111 -22163 3155
rect -22107 3111 -22063 3155
rect -22007 3111 -21963 3155
rect -21907 3111 -21863 3155
rect -21407 3111 -21363 3155
rect -21307 3111 -21263 3155
rect -21207 3111 -21163 3155
rect -21107 3111 -21063 3155
rect -21007 3111 -20963 3155
rect -20907 3111 -20863 3155
rect -20807 3111 -20763 3155
rect -20707 3111 -20663 3155
rect -20607 3111 -20563 3155
rect -20507 3111 -20463 3155
rect -20407 3111 -20363 3155
rect -20307 3111 -20263 3155
rect -20207 3111 -20163 3155
rect -20107 3111 -20063 3155
rect -20007 3111 -19963 3155
rect -19907 3111 -19863 3155
rect -27407 3011 -27363 3055
rect -27307 3011 -27263 3055
rect -27207 3011 -27163 3055
rect -27107 3011 -27063 3055
rect -27007 3011 -26963 3055
rect -26907 3011 -26863 3055
rect -26807 3011 -26763 3055
rect -26707 3011 -26663 3055
rect -26607 3011 -26563 3055
rect -26507 3011 -26463 3055
rect -26407 3011 -26363 3055
rect -26307 3011 -26263 3055
rect -26207 3011 -26163 3055
rect -26107 3011 -26063 3055
rect -26007 3011 -25963 3055
rect -25907 3011 -25863 3055
rect -25407 3011 -25363 3055
rect -25307 3011 -25263 3055
rect -25207 3011 -25163 3055
rect -25107 3011 -25063 3055
rect -25007 3011 -24963 3055
rect -24907 3011 -24863 3055
rect -24807 3011 -24763 3055
rect -24707 3011 -24663 3055
rect -24607 3011 -24563 3055
rect -24507 3011 -24463 3055
rect -24407 3011 -24363 3055
rect -24307 3011 -24263 3055
rect -24207 3011 -24163 3055
rect -24107 3011 -24063 3055
rect -24007 3011 -23963 3055
rect -23907 3011 -23863 3055
rect -23407 3011 -23363 3055
rect -23307 3011 -23263 3055
rect -23207 3011 -23163 3055
rect -23107 3011 -23063 3055
rect -23007 3011 -22963 3055
rect -22907 3011 -22863 3055
rect -22807 3011 -22763 3055
rect -22707 3011 -22663 3055
rect -22607 3011 -22563 3055
rect -22507 3011 -22463 3055
rect -22407 3011 -22363 3055
rect -22307 3011 -22263 3055
rect -22207 3011 -22163 3055
rect -22107 3011 -22063 3055
rect -22007 3011 -21963 3055
rect -21907 3011 -21863 3055
rect -21407 3011 -21363 3055
rect -21307 3011 -21263 3055
rect -21207 3011 -21163 3055
rect -21107 3011 -21063 3055
rect -21007 3011 -20963 3055
rect -20907 3011 -20863 3055
rect -20807 3011 -20763 3055
rect -20707 3011 -20663 3055
rect -20607 3011 -20563 3055
rect -20507 3011 -20463 3055
rect -20407 3011 -20363 3055
rect -20307 3011 -20263 3055
rect -20207 3011 -20163 3055
rect -20107 3011 -20063 3055
rect -20007 3011 -19963 3055
rect -19907 3011 -19863 3055
rect -27407 2911 -27363 2955
rect -27307 2911 -27263 2955
rect -27207 2911 -27163 2955
rect -27107 2911 -27063 2955
rect -27007 2911 -26963 2955
rect -26907 2911 -26863 2955
rect -26807 2911 -26763 2955
rect -26707 2911 -26663 2955
rect -26607 2911 -26563 2955
rect -26507 2911 -26463 2955
rect -26407 2911 -26363 2955
rect -26307 2911 -26263 2955
rect -26207 2911 -26163 2955
rect -26107 2911 -26063 2955
rect -26007 2911 -25963 2955
rect -25907 2911 -25863 2955
rect -25407 2911 -25363 2955
rect -25307 2911 -25263 2955
rect -25207 2911 -25163 2955
rect -25107 2911 -25063 2955
rect -25007 2911 -24963 2955
rect -24907 2911 -24863 2955
rect -24807 2911 -24763 2955
rect -24707 2911 -24663 2955
rect -24607 2911 -24563 2955
rect -24507 2911 -24463 2955
rect -24407 2911 -24363 2955
rect -24307 2911 -24263 2955
rect -24207 2911 -24163 2955
rect -24107 2911 -24063 2955
rect -24007 2911 -23963 2955
rect -23907 2911 -23863 2955
rect -23407 2911 -23363 2955
rect -23307 2911 -23263 2955
rect -23207 2911 -23163 2955
rect -23107 2911 -23063 2955
rect -23007 2911 -22963 2955
rect -22907 2911 -22863 2955
rect -22807 2911 -22763 2955
rect -22707 2911 -22663 2955
rect -22607 2911 -22563 2955
rect -22507 2911 -22463 2955
rect -22407 2911 -22363 2955
rect -22307 2911 -22263 2955
rect -22207 2911 -22163 2955
rect -22107 2911 -22063 2955
rect -22007 2911 -21963 2955
rect -21907 2911 -21863 2955
rect -21407 2911 -21363 2955
rect -21307 2911 -21263 2955
rect -21207 2911 -21163 2955
rect -21107 2911 -21063 2955
rect -21007 2911 -20963 2955
rect -20907 2911 -20863 2955
rect -20807 2911 -20763 2955
rect -20707 2911 -20663 2955
rect -20607 2911 -20563 2955
rect -20507 2911 -20463 2955
rect -20407 2911 -20363 2955
rect -20307 2911 -20263 2955
rect -20207 2911 -20163 2955
rect -20107 2911 -20063 2955
rect -20007 2911 -19963 2955
rect -19907 2911 -19863 2955
rect -27407 2811 -27363 2855
rect -27307 2811 -27263 2855
rect -27207 2811 -27163 2855
rect -27107 2811 -27063 2855
rect -27007 2811 -26963 2855
rect -26907 2811 -26863 2855
rect -26807 2811 -26763 2855
rect -26707 2811 -26663 2855
rect -26607 2811 -26563 2855
rect -26507 2811 -26463 2855
rect -26407 2811 -26363 2855
rect -26307 2811 -26263 2855
rect -26207 2811 -26163 2855
rect -26107 2811 -26063 2855
rect -26007 2811 -25963 2855
rect -25907 2811 -25863 2855
rect -25407 2811 -25363 2855
rect -25307 2811 -25263 2855
rect -25207 2811 -25163 2855
rect -25107 2811 -25063 2855
rect -25007 2811 -24963 2855
rect -24907 2811 -24863 2855
rect -24807 2811 -24763 2855
rect -24707 2811 -24663 2855
rect -24607 2811 -24563 2855
rect -24507 2811 -24463 2855
rect -24407 2811 -24363 2855
rect -24307 2811 -24263 2855
rect -24207 2811 -24163 2855
rect -24107 2811 -24063 2855
rect -24007 2811 -23963 2855
rect -23907 2811 -23863 2855
rect -23407 2811 -23363 2855
rect -23307 2811 -23263 2855
rect -23207 2811 -23163 2855
rect -23107 2811 -23063 2855
rect -23007 2811 -22963 2855
rect -22907 2811 -22863 2855
rect -22807 2811 -22763 2855
rect -22707 2811 -22663 2855
rect -22607 2811 -22563 2855
rect -22507 2811 -22463 2855
rect -22407 2811 -22363 2855
rect -22307 2811 -22263 2855
rect -22207 2811 -22163 2855
rect -22107 2811 -22063 2855
rect -22007 2811 -21963 2855
rect -21907 2811 -21863 2855
rect -21407 2811 -21363 2855
rect -21307 2811 -21263 2855
rect -21207 2811 -21163 2855
rect -21107 2811 -21063 2855
rect -21007 2811 -20963 2855
rect -20907 2811 -20863 2855
rect -20807 2811 -20763 2855
rect -20707 2811 -20663 2855
rect -20607 2811 -20563 2855
rect -20507 2811 -20463 2855
rect -20407 2811 -20363 2855
rect -20307 2811 -20263 2855
rect -20207 2811 -20163 2855
rect -20107 2811 -20063 2855
rect -20007 2811 -19963 2855
rect -19907 2811 -19863 2855
rect -27407 2711 -27363 2755
rect -27307 2711 -27263 2755
rect -27207 2711 -27163 2755
rect -27107 2711 -27063 2755
rect -27007 2711 -26963 2755
rect -26907 2711 -26863 2755
rect -26807 2711 -26763 2755
rect -26707 2711 -26663 2755
rect -26607 2711 -26563 2755
rect -26507 2711 -26463 2755
rect -26407 2711 -26363 2755
rect -26307 2711 -26263 2755
rect -26207 2711 -26163 2755
rect -26107 2711 -26063 2755
rect -26007 2711 -25963 2755
rect -25907 2711 -25863 2755
rect -25407 2711 -25363 2755
rect -25307 2711 -25263 2755
rect -25207 2711 -25163 2755
rect -25107 2711 -25063 2755
rect -25007 2711 -24963 2755
rect -24907 2711 -24863 2755
rect -24807 2711 -24763 2755
rect -24707 2711 -24663 2755
rect -24607 2711 -24563 2755
rect -24507 2711 -24463 2755
rect -24407 2711 -24363 2755
rect -24307 2711 -24263 2755
rect -24207 2711 -24163 2755
rect -24107 2711 -24063 2755
rect -24007 2711 -23963 2755
rect -23907 2711 -23863 2755
rect -23407 2711 -23363 2755
rect -23307 2711 -23263 2755
rect -23207 2711 -23163 2755
rect -23107 2711 -23063 2755
rect -23007 2711 -22963 2755
rect -22907 2711 -22863 2755
rect -22807 2711 -22763 2755
rect -22707 2711 -22663 2755
rect -22607 2711 -22563 2755
rect -22507 2711 -22463 2755
rect -22407 2711 -22363 2755
rect -22307 2711 -22263 2755
rect -22207 2711 -22163 2755
rect -22107 2711 -22063 2755
rect -22007 2711 -21963 2755
rect -21907 2711 -21863 2755
rect -21407 2711 -21363 2755
rect -21307 2711 -21263 2755
rect -21207 2711 -21163 2755
rect -21107 2711 -21063 2755
rect -21007 2711 -20963 2755
rect -20907 2711 -20863 2755
rect -20807 2711 -20763 2755
rect -20707 2711 -20663 2755
rect -20607 2711 -20563 2755
rect -20507 2711 -20463 2755
rect -20407 2711 -20363 2755
rect -20307 2711 -20263 2755
rect -20207 2711 -20163 2755
rect -20107 2711 -20063 2755
rect -20007 2711 -19963 2755
rect -19907 2711 -19863 2755
rect -27407 2611 -27363 2655
rect -27307 2611 -27263 2655
rect -27207 2611 -27163 2655
rect -27107 2611 -27063 2655
rect -27007 2611 -26963 2655
rect -26907 2611 -26863 2655
rect -26807 2611 -26763 2655
rect -26707 2611 -26663 2655
rect -26607 2611 -26563 2655
rect -26507 2611 -26463 2655
rect -26407 2611 -26363 2655
rect -26307 2611 -26263 2655
rect -26207 2611 -26163 2655
rect -26107 2611 -26063 2655
rect -26007 2611 -25963 2655
rect -25907 2611 -25863 2655
rect -25407 2611 -25363 2655
rect -25307 2611 -25263 2655
rect -25207 2611 -25163 2655
rect -25107 2611 -25063 2655
rect -25007 2611 -24963 2655
rect -24907 2611 -24863 2655
rect -24807 2611 -24763 2655
rect -24707 2611 -24663 2655
rect -24607 2611 -24563 2655
rect -24507 2611 -24463 2655
rect -24407 2611 -24363 2655
rect -24307 2611 -24263 2655
rect -24207 2611 -24163 2655
rect -24107 2611 -24063 2655
rect -24007 2611 -23963 2655
rect -23907 2611 -23863 2655
rect -23407 2611 -23363 2655
rect -23307 2611 -23263 2655
rect -23207 2611 -23163 2655
rect -23107 2611 -23063 2655
rect -23007 2611 -22963 2655
rect -22907 2611 -22863 2655
rect -22807 2611 -22763 2655
rect -22707 2611 -22663 2655
rect -22607 2611 -22563 2655
rect -22507 2611 -22463 2655
rect -22407 2611 -22363 2655
rect -22307 2611 -22263 2655
rect -22207 2611 -22163 2655
rect -22107 2611 -22063 2655
rect -22007 2611 -21963 2655
rect -21907 2611 -21863 2655
rect -21407 2611 -21363 2655
rect -21307 2611 -21263 2655
rect -21207 2611 -21163 2655
rect -21107 2611 -21063 2655
rect -21007 2611 -20963 2655
rect -20907 2611 -20863 2655
rect -20807 2611 -20763 2655
rect -20707 2611 -20663 2655
rect -20607 2611 -20563 2655
rect -20507 2611 -20463 2655
rect -20407 2611 -20363 2655
rect -20307 2611 -20263 2655
rect -20207 2611 -20163 2655
rect -20107 2611 -20063 2655
rect -20007 2611 -19963 2655
rect -19907 2611 -19863 2655
rect -27407 2511 -27363 2555
rect -27307 2511 -27263 2555
rect -27207 2511 -27163 2555
rect -27107 2511 -27063 2555
rect -27007 2511 -26963 2555
rect -26907 2511 -26863 2555
rect -26807 2511 -26763 2555
rect -26707 2511 -26663 2555
rect -26607 2511 -26563 2555
rect -26507 2511 -26463 2555
rect -26407 2511 -26363 2555
rect -26307 2511 -26263 2555
rect -26207 2511 -26163 2555
rect -26107 2511 -26063 2555
rect -26007 2511 -25963 2555
rect -25907 2511 -25863 2555
rect -25407 2511 -25363 2555
rect -25307 2511 -25263 2555
rect -25207 2511 -25163 2555
rect -25107 2511 -25063 2555
rect -25007 2511 -24963 2555
rect -24907 2511 -24863 2555
rect -24807 2511 -24763 2555
rect -24707 2511 -24663 2555
rect -24607 2511 -24563 2555
rect -24507 2511 -24463 2555
rect -24407 2511 -24363 2555
rect -24307 2511 -24263 2555
rect -24207 2511 -24163 2555
rect -24107 2511 -24063 2555
rect -24007 2511 -23963 2555
rect -23907 2511 -23863 2555
rect -23407 2511 -23363 2555
rect -23307 2511 -23263 2555
rect -23207 2511 -23163 2555
rect -23107 2511 -23063 2555
rect -23007 2511 -22963 2555
rect -22907 2511 -22863 2555
rect -22807 2511 -22763 2555
rect -22707 2511 -22663 2555
rect -22607 2511 -22563 2555
rect -22507 2511 -22463 2555
rect -22407 2511 -22363 2555
rect -22307 2511 -22263 2555
rect -22207 2511 -22163 2555
rect -22107 2511 -22063 2555
rect -22007 2511 -21963 2555
rect -21907 2511 -21863 2555
rect -21407 2511 -21363 2555
rect -21307 2511 -21263 2555
rect -21207 2511 -21163 2555
rect -21107 2511 -21063 2555
rect -21007 2511 -20963 2555
rect -20907 2511 -20863 2555
rect -20807 2511 -20763 2555
rect -20707 2511 -20663 2555
rect -20607 2511 -20563 2555
rect -20507 2511 -20463 2555
rect -20407 2511 -20363 2555
rect -20307 2511 -20263 2555
rect -20207 2511 -20163 2555
rect -20107 2511 -20063 2555
rect -20007 2511 -19963 2555
rect -19907 2511 -19863 2555
rect -27407 2411 -27363 2455
rect -27307 2411 -27263 2455
rect -27207 2411 -27163 2455
rect -27107 2411 -27063 2455
rect -27007 2411 -26963 2455
rect -26907 2411 -26863 2455
rect -26807 2411 -26763 2455
rect -26707 2411 -26663 2455
rect -26607 2411 -26563 2455
rect -26507 2411 -26463 2455
rect -26407 2411 -26363 2455
rect -26307 2411 -26263 2455
rect -26207 2411 -26163 2455
rect -26107 2411 -26063 2455
rect -26007 2411 -25963 2455
rect -25907 2411 -25863 2455
rect -25407 2411 -25363 2455
rect -25307 2411 -25263 2455
rect -25207 2411 -25163 2455
rect -25107 2411 -25063 2455
rect -25007 2411 -24963 2455
rect -24907 2411 -24863 2455
rect -24807 2411 -24763 2455
rect -24707 2411 -24663 2455
rect -24607 2411 -24563 2455
rect -24507 2411 -24463 2455
rect -24407 2411 -24363 2455
rect -24307 2411 -24263 2455
rect -24207 2411 -24163 2455
rect -24107 2411 -24063 2455
rect -24007 2411 -23963 2455
rect -23907 2411 -23863 2455
rect -23407 2411 -23363 2455
rect -23307 2411 -23263 2455
rect -23207 2411 -23163 2455
rect -23107 2411 -23063 2455
rect -23007 2411 -22963 2455
rect -22907 2411 -22863 2455
rect -22807 2411 -22763 2455
rect -22707 2411 -22663 2455
rect -22607 2411 -22563 2455
rect -22507 2411 -22463 2455
rect -22407 2411 -22363 2455
rect -22307 2411 -22263 2455
rect -22207 2411 -22163 2455
rect -22107 2411 -22063 2455
rect -22007 2411 -21963 2455
rect -21907 2411 -21863 2455
rect -21407 2411 -21363 2455
rect -21307 2411 -21263 2455
rect -21207 2411 -21163 2455
rect -21107 2411 -21063 2455
rect -21007 2411 -20963 2455
rect -20907 2411 -20863 2455
rect -20807 2411 -20763 2455
rect -20707 2411 -20663 2455
rect -20607 2411 -20563 2455
rect -20507 2411 -20463 2455
rect -20407 2411 -20363 2455
rect -20307 2411 -20263 2455
rect -20207 2411 -20163 2455
rect -20107 2411 -20063 2455
rect -20007 2411 -19963 2455
rect -19907 2411 -19863 2455
rect -27407 2311 -27363 2355
rect -27307 2311 -27263 2355
rect -27207 2311 -27163 2355
rect -27107 2311 -27063 2355
rect -27007 2311 -26963 2355
rect -26907 2311 -26863 2355
rect -26807 2311 -26763 2355
rect -26707 2311 -26663 2355
rect -26607 2311 -26563 2355
rect -26507 2311 -26463 2355
rect -26407 2311 -26363 2355
rect -26307 2311 -26263 2355
rect -26207 2311 -26163 2355
rect -26107 2311 -26063 2355
rect -26007 2311 -25963 2355
rect -25907 2311 -25863 2355
rect -25407 2311 -25363 2355
rect -25307 2311 -25263 2355
rect -25207 2311 -25163 2355
rect -25107 2311 -25063 2355
rect -25007 2311 -24963 2355
rect -24907 2311 -24863 2355
rect -24807 2311 -24763 2355
rect -24707 2311 -24663 2355
rect -24607 2311 -24563 2355
rect -24507 2311 -24463 2355
rect -24407 2311 -24363 2355
rect -24307 2311 -24263 2355
rect -24207 2311 -24163 2355
rect -24107 2311 -24063 2355
rect -24007 2311 -23963 2355
rect -23907 2311 -23863 2355
rect -23407 2311 -23363 2355
rect -23307 2311 -23263 2355
rect -23207 2311 -23163 2355
rect -23107 2311 -23063 2355
rect -23007 2311 -22963 2355
rect -22907 2311 -22863 2355
rect -22807 2311 -22763 2355
rect -22707 2311 -22663 2355
rect -22607 2311 -22563 2355
rect -22507 2311 -22463 2355
rect -22407 2311 -22363 2355
rect -22307 2311 -22263 2355
rect -22207 2311 -22163 2355
rect -22107 2311 -22063 2355
rect -22007 2311 -21963 2355
rect -21907 2311 -21863 2355
rect -21407 2311 -21363 2355
rect -21307 2311 -21263 2355
rect -21207 2311 -21163 2355
rect -21107 2311 -21063 2355
rect -21007 2311 -20963 2355
rect -20907 2311 -20863 2355
rect -20807 2311 -20763 2355
rect -20707 2311 -20663 2355
rect -20607 2311 -20563 2355
rect -20507 2311 -20463 2355
rect -20407 2311 -20363 2355
rect -20307 2311 -20263 2355
rect -20207 2311 -20163 2355
rect -20107 2311 -20063 2355
rect -20007 2311 -19963 2355
rect -19907 2311 -19863 2355
rect -27407 2211 -27363 2255
rect -27307 2211 -27263 2255
rect -27207 2211 -27163 2255
rect -27107 2211 -27063 2255
rect -27007 2211 -26963 2255
rect -26907 2211 -26863 2255
rect -26807 2211 -26763 2255
rect -26707 2211 -26663 2255
rect -26607 2211 -26563 2255
rect -26507 2211 -26463 2255
rect -26407 2211 -26363 2255
rect -26307 2211 -26263 2255
rect -26207 2211 -26163 2255
rect -26107 2211 -26063 2255
rect -26007 2211 -25963 2255
rect -25907 2211 -25863 2255
rect -25407 2211 -25363 2255
rect -25307 2211 -25263 2255
rect -25207 2211 -25163 2255
rect -25107 2211 -25063 2255
rect -25007 2211 -24963 2255
rect -24907 2211 -24863 2255
rect -24807 2211 -24763 2255
rect -24707 2211 -24663 2255
rect -24607 2211 -24563 2255
rect -24507 2211 -24463 2255
rect -24407 2211 -24363 2255
rect -24307 2211 -24263 2255
rect -24207 2211 -24163 2255
rect -24107 2211 -24063 2255
rect -24007 2211 -23963 2255
rect -23907 2211 -23863 2255
rect -23407 2211 -23363 2255
rect -23307 2211 -23263 2255
rect -23207 2211 -23163 2255
rect -23107 2211 -23063 2255
rect -23007 2211 -22963 2255
rect -22907 2211 -22863 2255
rect -22807 2211 -22763 2255
rect -22707 2211 -22663 2255
rect -22607 2211 -22563 2255
rect -22507 2211 -22463 2255
rect -22407 2211 -22363 2255
rect -22307 2211 -22263 2255
rect -22207 2211 -22163 2255
rect -22107 2211 -22063 2255
rect -22007 2211 -21963 2255
rect -21907 2211 -21863 2255
rect -21407 2211 -21363 2255
rect -21307 2211 -21263 2255
rect -21207 2211 -21163 2255
rect -21107 2211 -21063 2255
rect -21007 2211 -20963 2255
rect -20907 2211 -20863 2255
rect -20807 2211 -20763 2255
rect -20707 2211 -20663 2255
rect -20607 2211 -20563 2255
rect -20507 2211 -20463 2255
rect -20407 2211 -20363 2255
rect -20307 2211 -20263 2255
rect -20207 2211 -20163 2255
rect -20107 2211 -20063 2255
rect -20007 2211 -19963 2255
rect -19907 2211 -19863 2255
rect -27407 2111 -27363 2155
rect -27307 2111 -27263 2155
rect -27207 2111 -27163 2155
rect -27107 2111 -27063 2155
rect -27007 2111 -26963 2155
rect -26907 2111 -26863 2155
rect -26807 2111 -26763 2155
rect -26707 2111 -26663 2155
rect -26607 2111 -26563 2155
rect -26507 2111 -26463 2155
rect -26407 2111 -26363 2155
rect -26307 2111 -26263 2155
rect -26207 2111 -26163 2155
rect -26107 2111 -26063 2155
rect -26007 2111 -25963 2155
rect -25907 2111 -25863 2155
rect -25407 2111 -25363 2155
rect -25307 2111 -25263 2155
rect -25207 2111 -25163 2155
rect -25107 2111 -25063 2155
rect -25007 2111 -24963 2155
rect -24907 2111 -24863 2155
rect -24807 2111 -24763 2155
rect -24707 2111 -24663 2155
rect -24607 2111 -24563 2155
rect -24507 2111 -24463 2155
rect -24407 2111 -24363 2155
rect -24307 2111 -24263 2155
rect -24207 2111 -24163 2155
rect -24107 2111 -24063 2155
rect -24007 2111 -23963 2155
rect -23907 2111 -23863 2155
rect -23407 2111 -23363 2155
rect -23307 2111 -23263 2155
rect -23207 2111 -23163 2155
rect -23107 2111 -23063 2155
rect -23007 2111 -22963 2155
rect -22907 2111 -22863 2155
rect -22807 2111 -22763 2155
rect -22707 2111 -22663 2155
rect -22607 2111 -22563 2155
rect -22507 2111 -22463 2155
rect -22407 2111 -22363 2155
rect -22307 2111 -22263 2155
rect -22207 2111 -22163 2155
rect -22107 2111 -22063 2155
rect -22007 2111 -21963 2155
rect -21907 2111 -21863 2155
rect -21407 2111 -21363 2155
rect -21307 2111 -21263 2155
rect -21207 2111 -21163 2155
rect -21107 2111 -21063 2155
rect -21007 2111 -20963 2155
rect -20907 2111 -20863 2155
rect -20807 2111 -20763 2155
rect -20707 2111 -20663 2155
rect -20607 2111 -20563 2155
rect -20507 2111 -20463 2155
rect -20407 2111 -20363 2155
rect -20307 2111 -20263 2155
rect -20207 2111 -20163 2155
rect -20107 2111 -20063 2155
rect -20007 2111 -19963 2155
rect -19907 2111 -19863 2155
rect -27407 2011 -27363 2055
rect -27307 2011 -27263 2055
rect -27207 2011 -27163 2055
rect -27107 2011 -27063 2055
rect -27007 2011 -26963 2055
rect -26907 2011 -26863 2055
rect -26807 2011 -26763 2055
rect -26707 2011 -26663 2055
rect -26607 2011 -26563 2055
rect -26507 2011 -26463 2055
rect -26407 2011 -26363 2055
rect -26307 2011 -26263 2055
rect -26207 2011 -26163 2055
rect -26107 2011 -26063 2055
rect -26007 2011 -25963 2055
rect -25907 2011 -25863 2055
rect -25407 2011 -25363 2055
rect -25307 2011 -25263 2055
rect -25207 2011 -25163 2055
rect -25107 2011 -25063 2055
rect -25007 2011 -24963 2055
rect -24907 2011 -24863 2055
rect -24807 2011 -24763 2055
rect -24707 2011 -24663 2055
rect -24607 2011 -24563 2055
rect -24507 2011 -24463 2055
rect -24407 2011 -24363 2055
rect -24307 2011 -24263 2055
rect -24207 2011 -24163 2055
rect -24107 2011 -24063 2055
rect -24007 2011 -23963 2055
rect -23907 2011 -23863 2055
rect -23407 2011 -23363 2055
rect -23307 2011 -23263 2055
rect -23207 2011 -23163 2055
rect -23107 2011 -23063 2055
rect -23007 2011 -22963 2055
rect -22907 2011 -22863 2055
rect -22807 2011 -22763 2055
rect -22707 2011 -22663 2055
rect -22607 2011 -22563 2055
rect -22507 2011 -22463 2055
rect -22407 2011 -22363 2055
rect -22307 2011 -22263 2055
rect -22207 2011 -22163 2055
rect -22107 2011 -22063 2055
rect -22007 2011 -21963 2055
rect -21907 2011 -21863 2055
rect -21407 2011 -21363 2055
rect -21307 2011 -21263 2055
rect -21207 2011 -21163 2055
rect -21107 2011 -21063 2055
rect -21007 2011 -20963 2055
rect -20907 2011 -20863 2055
rect -20807 2011 -20763 2055
rect -20707 2011 -20663 2055
rect -20607 2011 -20563 2055
rect -20507 2011 -20463 2055
rect -20407 2011 -20363 2055
rect -20307 2011 -20263 2055
rect -20207 2011 -20163 2055
rect -20107 2011 -20063 2055
rect -20007 2011 -19963 2055
rect -19907 2011 -19863 2055
rect -12772 -7374 -12552 -7154
rect -12302 -7374 -12082 -7154
rect -11832 -7374 -11612 -7154
rect -11362 -7374 -11142 -7154
rect -10892 -7374 -10672 -7154
rect -10422 -7374 -10202 -7154
rect -9952 -7374 -9732 -7154
rect -9482 -7374 -9262 -7154
rect -9012 -7374 -8792 -7154
rect -8542 -7374 -8322 -7154
rect -8072 -7374 -7852 -7154
rect -7602 -7374 -7382 -7154
rect -7132 -7374 -6912 -7154
rect -6662 -7374 -6442 -7154
rect -12784 -13656 -12564 -13436
rect -12314 -13656 -12094 -13436
rect -11844 -13656 -11624 -13436
rect -11374 -13656 -11154 -13436
rect -10904 -13656 -10684 -13436
rect -10434 -13656 -10214 -13436
rect -9964 -13656 -9744 -13436
rect -9494 -13656 -9274 -13436
rect -9024 -13656 -8804 -13436
rect -8554 -13656 -8334 -13436
rect -8084 -13656 -7864 -13436
rect -7614 -13656 -7394 -13436
rect -7144 -13656 -6924 -13436
rect -6674 -13656 -6454 -13436
rect 9195 -9800 9239 -9756
rect 9295 -9800 9339 -9756
rect 9395 -9800 9439 -9756
rect 9495 -9800 9539 -9756
rect 9595 -9800 9639 -9756
rect 9695 -9800 9739 -9756
rect 9795 -9800 9839 -9756
rect 9895 -9800 9939 -9756
rect 9995 -9800 10039 -9756
rect 10095 -9800 10139 -9756
rect 10195 -9800 10239 -9756
rect 10295 -9800 10339 -9756
rect 10395 -9800 10439 -9756
rect 10495 -9800 10539 -9756
rect 10595 -9800 10639 -9756
rect 10695 -9800 10739 -9756
rect 11195 -9800 11239 -9756
rect 11295 -9800 11339 -9756
rect 11395 -9800 11439 -9756
rect 11495 -9800 11539 -9756
rect 11595 -9800 11639 -9756
rect 11695 -9800 11739 -9756
rect 11795 -9800 11839 -9756
rect 11895 -9800 11939 -9756
rect 11995 -9800 12039 -9756
rect 12095 -9800 12139 -9756
rect 12195 -9800 12239 -9756
rect 12295 -9800 12339 -9756
rect 12395 -9800 12439 -9756
rect 12495 -9800 12539 -9756
rect 12595 -9800 12639 -9756
rect 12695 -9800 12739 -9756
rect 13195 -9800 13239 -9756
rect 13295 -9800 13339 -9756
rect 13395 -9800 13439 -9756
rect 13495 -9800 13539 -9756
rect 13595 -9800 13639 -9756
rect 13695 -9800 13739 -9756
rect 13795 -9800 13839 -9756
rect 13895 -9800 13939 -9756
rect 13995 -9800 14039 -9756
rect 14095 -9800 14139 -9756
rect 14195 -9800 14239 -9756
rect 14295 -9800 14339 -9756
rect 14395 -9800 14439 -9756
rect 14495 -9800 14539 -9756
rect 14595 -9800 14639 -9756
rect 14695 -9800 14739 -9756
rect 15195 -9800 15239 -9756
rect 15295 -9800 15339 -9756
rect 15395 -9800 15439 -9756
rect 15495 -9800 15539 -9756
rect 15595 -9800 15639 -9756
rect 15695 -9800 15739 -9756
rect 15795 -9800 15839 -9756
rect 15895 -9800 15939 -9756
rect 15995 -9800 16039 -9756
rect 16095 -9800 16139 -9756
rect 16195 -9800 16239 -9756
rect 16295 -9800 16339 -9756
rect 16395 -9800 16439 -9756
rect 16495 -9800 16539 -9756
rect 16595 -9800 16639 -9756
rect 16695 -9800 16739 -9756
rect 9195 -9900 9239 -9856
rect 9295 -9900 9339 -9856
rect 9395 -9900 9439 -9856
rect 9495 -9900 9539 -9856
rect 9595 -9900 9639 -9856
rect 9695 -9900 9739 -9856
rect 9795 -9900 9839 -9856
rect 9895 -9900 9939 -9856
rect 9995 -9900 10039 -9856
rect 10095 -9900 10139 -9856
rect 10195 -9900 10239 -9856
rect 10295 -9900 10339 -9856
rect 10395 -9900 10439 -9856
rect 10495 -9900 10539 -9856
rect 10595 -9900 10639 -9856
rect 10695 -9900 10739 -9856
rect 11195 -9900 11239 -9856
rect 11295 -9900 11339 -9856
rect 11395 -9900 11439 -9856
rect 11495 -9900 11539 -9856
rect 11595 -9900 11639 -9856
rect 11695 -9900 11739 -9856
rect 11795 -9900 11839 -9856
rect 11895 -9900 11939 -9856
rect 11995 -9900 12039 -9856
rect 12095 -9900 12139 -9856
rect 12195 -9900 12239 -9856
rect 12295 -9900 12339 -9856
rect 12395 -9900 12439 -9856
rect 12495 -9900 12539 -9856
rect 12595 -9900 12639 -9856
rect 12695 -9900 12739 -9856
rect 13195 -9900 13239 -9856
rect 13295 -9900 13339 -9856
rect 13395 -9900 13439 -9856
rect 13495 -9900 13539 -9856
rect 13595 -9900 13639 -9856
rect 13695 -9900 13739 -9856
rect 13795 -9900 13839 -9856
rect 13895 -9900 13939 -9856
rect 13995 -9900 14039 -9856
rect 14095 -9900 14139 -9856
rect 14195 -9900 14239 -9856
rect 14295 -9900 14339 -9856
rect 14395 -9900 14439 -9856
rect 14495 -9900 14539 -9856
rect 14595 -9900 14639 -9856
rect 14695 -9900 14739 -9856
rect 15195 -9900 15239 -9856
rect 15295 -9900 15339 -9856
rect 15395 -9900 15439 -9856
rect 15495 -9900 15539 -9856
rect 15595 -9900 15639 -9856
rect 15695 -9900 15739 -9856
rect 15795 -9900 15839 -9856
rect 15895 -9900 15939 -9856
rect 15995 -9900 16039 -9856
rect 16095 -9900 16139 -9856
rect 16195 -9900 16239 -9856
rect 16295 -9900 16339 -9856
rect 16395 -9900 16439 -9856
rect 16495 -9900 16539 -9856
rect 16595 -9900 16639 -9856
rect 16695 -9900 16739 -9856
rect 9195 -10000 9239 -9956
rect 9295 -10000 9339 -9956
rect 9395 -10000 9439 -9956
rect 9495 -10000 9539 -9956
rect 9595 -10000 9639 -9956
rect 9695 -10000 9739 -9956
rect 9795 -10000 9839 -9956
rect 9895 -10000 9939 -9956
rect 9995 -10000 10039 -9956
rect 10095 -10000 10139 -9956
rect 10195 -10000 10239 -9956
rect 10295 -10000 10339 -9956
rect 10395 -10000 10439 -9956
rect 10495 -10000 10539 -9956
rect 10595 -10000 10639 -9956
rect 10695 -10000 10739 -9956
rect 11195 -10000 11239 -9956
rect 11295 -10000 11339 -9956
rect 11395 -10000 11439 -9956
rect 11495 -10000 11539 -9956
rect 11595 -10000 11639 -9956
rect 11695 -10000 11739 -9956
rect 11795 -10000 11839 -9956
rect 11895 -10000 11939 -9956
rect 11995 -10000 12039 -9956
rect 12095 -10000 12139 -9956
rect 12195 -10000 12239 -9956
rect 12295 -10000 12339 -9956
rect 12395 -10000 12439 -9956
rect 12495 -10000 12539 -9956
rect 12595 -10000 12639 -9956
rect 12695 -10000 12739 -9956
rect 13195 -10000 13239 -9956
rect 13295 -10000 13339 -9956
rect 13395 -10000 13439 -9956
rect 13495 -10000 13539 -9956
rect 13595 -10000 13639 -9956
rect 13695 -10000 13739 -9956
rect 13795 -10000 13839 -9956
rect 13895 -10000 13939 -9956
rect 13995 -10000 14039 -9956
rect 14095 -10000 14139 -9956
rect 14195 -10000 14239 -9956
rect 14295 -10000 14339 -9956
rect 14395 -10000 14439 -9956
rect 14495 -10000 14539 -9956
rect 14595 -10000 14639 -9956
rect 14695 -10000 14739 -9956
rect 15195 -10000 15239 -9956
rect 15295 -10000 15339 -9956
rect 15395 -10000 15439 -9956
rect 15495 -10000 15539 -9956
rect 15595 -10000 15639 -9956
rect 15695 -10000 15739 -9956
rect 15795 -10000 15839 -9956
rect 15895 -10000 15939 -9956
rect 15995 -10000 16039 -9956
rect 16095 -10000 16139 -9956
rect 16195 -10000 16239 -9956
rect 16295 -10000 16339 -9956
rect 16395 -10000 16439 -9956
rect 16495 -10000 16539 -9956
rect 16595 -10000 16639 -9956
rect 16695 -10000 16739 -9956
rect 9195 -10100 9239 -10056
rect 9295 -10100 9339 -10056
rect 9395 -10100 9439 -10056
rect 9495 -10100 9539 -10056
rect 9595 -10100 9639 -10056
rect 9695 -10100 9739 -10056
rect 9795 -10100 9839 -10056
rect 9895 -10100 9939 -10056
rect 9995 -10100 10039 -10056
rect 10095 -10100 10139 -10056
rect 10195 -10100 10239 -10056
rect 10295 -10100 10339 -10056
rect 10395 -10100 10439 -10056
rect 10495 -10100 10539 -10056
rect 10595 -10100 10639 -10056
rect 10695 -10100 10739 -10056
rect 11195 -10100 11239 -10056
rect 11295 -10100 11339 -10056
rect 11395 -10100 11439 -10056
rect 11495 -10100 11539 -10056
rect 11595 -10100 11639 -10056
rect 11695 -10100 11739 -10056
rect 11795 -10100 11839 -10056
rect 11895 -10100 11939 -10056
rect 11995 -10100 12039 -10056
rect 12095 -10100 12139 -10056
rect 12195 -10100 12239 -10056
rect 12295 -10100 12339 -10056
rect 12395 -10100 12439 -10056
rect 12495 -10100 12539 -10056
rect 12595 -10100 12639 -10056
rect 12695 -10100 12739 -10056
rect 13195 -10100 13239 -10056
rect 13295 -10100 13339 -10056
rect 13395 -10100 13439 -10056
rect 13495 -10100 13539 -10056
rect 13595 -10100 13639 -10056
rect 13695 -10100 13739 -10056
rect 13795 -10100 13839 -10056
rect 13895 -10100 13939 -10056
rect 13995 -10100 14039 -10056
rect 14095 -10100 14139 -10056
rect 14195 -10100 14239 -10056
rect 14295 -10100 14339 -10056
rect 14395 -10100 14439 -10056
rect 14495 -10100 14539 -10056
rect 14595 -10100 14639 -10056
rect 14695 -10100 14739 -10056
rect 15195 -10100 15239 -10056
rect 15295 -10100 15339 -10056
rect 15395 -10100 15439 -10056
rect 15495 -10100 15539 -10056
rect 15595 -10100 15639 -10056
rect 15695 -10100 15739 -10056
rect 15795 -10100 15839 -10056
rect 15895 -10100 15939 -10056
rect 15995 -10100 16039 -10056
rect 16095 -10100 16139 -10056
rect 16195 -10100 16239 -10056
rect 16295 -10100 16339 -10056
rect 16395 -10100 16439 -10056
rect 16495 -10100 16539 -10056
rect 16595 -10100 16639 -10056
rect 16695 -10100 16739 -10056
rect 9195 -10200 9239 -10156
rect 9295 -10200 9339 -10156
rect 9395 -10200 9439 -10156
rect 9495 -10200 9539 -10156
rect 9595 -10200 9639 -10156
rect 9695 -10200 9739 -10156
rect 9795 -10200 9839 -10156
rect 9895 -10200 9939 -10156
rect 9995 -10200 10039 -10156
rect 10095 -10200 10139 -10156
rect 10195 -10200 10239 -10156
rect 10295 -10200 10339 -10156
rect 10395 -10200 10439 -10156
rect 10495 -10200 10539 -10156
rect 10595 -10200 10639 -10156
rect 10695 -10200 10739 -10156
rect 11195 -10200 11239 -10156
rect 11295 -10200 11339 -10156
rect 11395 -10200 11439 -10156
rect 11495 -10200 11539 -10156
rect 11595 -10200 11639 -10156
rect 11695 -10200 11739 -10156
rect 11795 -10200 11839 -10156
rect 11895 -10200 11939 -10156
rect 11995 -10200 12039 -10156
rect 12095 -10200 12139 -10156
rect 12195 -10200 12239 -10156
rect 12295 -10200 12339 -10156
rect 12395 -10200 12439 -10156
rect 12495 -10200 12539 -10156
rect 12595 -10200 12639 -10156
rect 12695 -10200 12739 -10156
rect 13195 -10200 13239 -10156
rect 13295 -10200 13339 -10156
rect 13395 -10200 13439 -10156
rect 13495 -10200 13539 -10156
rect 13595 -10200 13639 -10156
rect 13695 -10200 13739 -10156
rect 13795 -10200 13839 -10156
rect 13895 -10200 13939 -10156
rect 13995 -10200 14039 -10156
rect 14095 -10200 14139 -10156
rect 14195 -10200 14239 -10156
rect 14295 -10200 14339 -10156
rect 14395 -10200 14439 -10156
rect 14495 -10200 14539 -10156
rect 14595 -10200 14639 -10156
rect 14695 -10200 14739 -10156
rect 15195 -10200 15239 -10156
rect 15295 -10200 15339 -10156
rect 15395 -10200 15439 -10156
rect 15495 -10200 15539 -10156
rect 15595 -10200 15639 -10156
rect 15695 -10200 15739 -10156
rect 15795 -10200 15839 -10156
rect 15895 -10200 15939 -10156
rect 15995 -10200 16039 -10156
rect 16095 -10200 16139 -10156
rect 16195 -10200 16239 -10156
rect 16295 -10200 16339 -10156
rect 16395 -10200 16439 -10156
rect 16495 -10200 16539 -10156
rect 16595 -10200 16639 -10156
rect 16695 -10200 16739 -10156
rect 9195 -10300 9239 -10256
rect 9295 -10300 9339 -10256
rect 9395 -10300 9439 -10256
rect 9495 -10300 9539 -10256
rect 9595 -10300 9639 -10256
rect 9695 -10300 9739 -10256
rect 9795 -10300 9839 -10256
rect 9895 -10300 9939 -10256
rect 9995 -10300 10039 -10256
rect 10095 -10300 10139 -10256
rect 10195 -10300 10239 -10256
rect 10295 -10300 10339 -10256
rect 10395 -10300 10439 -10256
rect 10495 -10300 10539 -10256
rect 10595 -10300 10639 -10256
rect 10695 -10300 10739 -10256
rect 11195 -10300 11239 -10256
rect 11295 -10300 11339 -10256
rect 11395 -10300 11439 -10256
rect 11495 -10300 11539 -10256
rect 11595 -10300 11639 -10256
rect 11695 -10300 11739 -10256
rect 11795 -10300 11839 -10256
rect 11895 -10300 11939 -10256
rect 11995 -10300 12039 -10256
rect 12095 -10300 12139 -10256
rect 12195 -10300 12239 -10256
rect 12295 -10300 12339 -10256
rect 12395 -10300 12439 -10256
rect 12495 -10300 12539 -10256
rect 12595 -10300 12639 -10256
rect 12695 -10300 12739 -10256
rect 13195 -10300 13239 -10256
rect 13295 -10300 13339 -10256
rect 13395 -10300 13439 -10256
rect 13495 -10300 13539 -10256
rect 13595 -10300 13639 -10256
rect 13695 -10300 13739 -10256
rect 13795 -10300 13839 -10256
rect 13895 -10300 13939 -10256
rect 13995 -10300 14039 -10256
rect 14095 -10300 14139 -10256
rect 14195 -10300 14239 -10256
rect 14295 -10300 14339 -10256
rect 14395 -10300 14439 -10256
rect 14495 -10300 14539 -10256
rect 14595 -10300 14639 -10256
rect 14695 -10300 14739 -10256
rect 15195 -10300 15239 -10256
rect 15295 -10300 15339 -10256
rect 15395 -10300 15439 -10256
rect 15495 -10300 15539 -10256
rect 15595 -10300 15639 -10256
rect 15695 -10300 15739 -10256
rect 15795 -10300 15839 -10256
rect 15895 -10300 15939 -10256
rect 15995 -10300 16039 -10256
rect 16095 -10300 16139 -10256
rect 16195 -10300 16239 -10256
rect 16295 -10300 16339 -10256
rect 16395 -10300 16439 -10256
rect 16495 -10300 16539 -10256
rect 16595 -10300 16639 -10256
rect 16695 -10300 16739 -10256
rect 9195 -10400 9239 -10356
rect 9295 -10400 9339 -10356
rect 9395 -10400 9439 -10356
rect 9495 -10400 9539 -10356
rect 9595 -10400 9639 -10356
rect 9695 -10400 9739 -10356
rect 9795 -10400 9839 -10356
rect 9895 -10400 9939 -10356
rect 9995 -10400 10039 -10356
rect 10095 -10400 10139 -10356
rect 10195 -10400 10239 -10356
rect 10295 -10400 10339 -10356
rect 10395 -10400 10439 -10356
rect 10495 -10400 10539 -10356
rect 10595 -10400 10639 -10356
rect 10695 -10400 10739 -10356
rect 11195 -10400 11239 -10356
rect 11295 -10400 11339 -10356
rect 11395 -10400 11439 -10356
rect 11495 -10400 11539 -10356
rect 11595 -10400 11639 -10356
rect 11695 -10400 11739 -10356
rect 11795 -10400 11839 -10356
rect 11895 -10400 11939 -10356
rect 11995 -10400 12039 -10356
rect 12095 -10400 12139 -10356
rect 12195 -10400 12239 -10356
rect 12295 -10400 12339 -10356
rect 12395 -10400 12439 -10356
rect 12495 -10400 12539 -10356
rect 12595 -10400 12639 -10356
rect 12695 -10400 12739 -10356
rect 13195 -10400 13239 -10356
rect 13295 -10400 13339 -10356
rect 13395 -10400 13439 -10356
rect 13495 -10400 13539 -10356
rect 13595 -10400 13639 -10356
rect 13695 -10400 13739 -10356
rect 13795 -10400 13839 -10356
rect 13895 -10400 13939 -10356
rect 13995 -10400 14039 -10356
rect 14095 -10400 14139 -10356
rect 14195 -10400 14239 -10356
rect 14295 -10400 14339 -10356
rect 14395 -10400 14439 -10356
rect 14495 -10400 14539 -10356
rect 14595 -10400 14639 -10356
rect 14695 -10400 14739 -10356
rect 15195 -10400 15239 -10356
rect 15295 -10400 15339 -10356
rect 15395 -10400 15439 -10356
rect 15495 -10400 15539 -10356
rect 15595 -10400 15639 -10356
rect 15695 -10400 15739 -10356
rect 15795 -10400 15839 -10356
rect 15895 -10400 15939 -10356
rect 15995 -10400 16039 -10356
rect 16095 -10400 16139 -10356
rect 16195 -10400 16239 -10356
rect 16295 -10400 16339 -10356
rect 16395 -10400 16439 -10356
rect 16495 -10400 16539 -10356
rect 16595 -10400 16639 -10356
rect 16695 -10400 16739 -10356
rect 9195 -10500 9239 -10456
rect 9295 -10500 9339 -10456
rect 9395 -10500 9439 -10456
rect 9495 -10500 9539 -10456
rect 9595 -10500 9639 -10456
rect 9695 -10500 9739 -10456
rect 9795 -10500 9839 -10456
rect 9895 -10500 9939 -10456
rect 9995 -10500 10039 -10456
rect 10095 -10500 10139 -10456
rect 10195 -10500 10239 -10456
rect 10295 -10500 10339 -10456
rect 10395 -10500 10439 -10456
rect 10495 -10500 10539 -10456
rect 10595 -10500 10639 -10456
rect 10695 -10500 10739 -10456
rect 11195 -10500 11239 -10456
rect 11295 -10500 11339 -10456
rect 11395 -10500 11439 -10456
rect 11495 -10500 11539 -10456
rect 11595 -10500 11639 -10456
rect 11695 -10500 11739 -10456
rect 11795 -10500 11839 -10456
rect 11895 -10500 11939 -10456
rect 11995 -10500 12039 -10456
rect 12095 -10500 12139 -10456
rect 12195 -10500 12239 -10456
rect 12295 -10500 12339 -10456
rect 12395 -10500 12439 -10456
rect 12495 -10500 12539 -10456
rect 12595 -10500 12639 -10456
rect 12695 -10500 12739 -10456
rect 13195 -10500 13239 -10456
rect 13295 -10500 13339 -10456
rect 13395 -10500 13439 -10456
rect 13495 -10500 13539 -10456
rect 13595 -10500 13639 -10456
rect 13695 -10500 13739 -10456
rect 13795 -10500 13839 -10456
rect 13895 -10500 13939 -10456
rect 13995 -10500 14039 -10456
rect 14095 -10500 14139 -10456
rect 14195 -10500 14239 -10456
rect 14295 -10500 14339 -10456
rect 14395 -10500 14439 -10456
rect 14495 -10500 14539 -10456
rect 14595 -10500 14639 -10456
rect 14695 -10500 14739 -10456
rect 15195 -10500 15239 -10456
rect 15295 -10500 15339 -10456
rect 15395 -10500 15439 -10456
rect 15495 -10500 15539 -10456
rect 15595 -10500 15639 -10456
rect 15695 -10500 15739 -10456
rect 15795 -10500 15839 -10456
rect 15895 -10500 15939 -10456
rect 15995 -10500 16039 -10456
rect 16095 -10500 16139 -10456
rect 16195 -10500 16239 -10456
rect 16295 -10500 16339 -10456
rect 16395 -10500 16439 -10456
rect 16495 -10500 16539 -10456
rect 16595 -10500 16639 -10456
rect 16695 -10500 16739 -10456
rect 9195 -10600 9239 -10556
rect 9295 -10600 9339 -10556
rect 9395 -10600 9439 -10556
rect 9495 -10600 9539 -10556
rect 9595 -10600 9639 -10556
rect 9695 -10600 9739 -10556
rect 9795 -10600 9839 -10556
rect 9895 -10600 9939 -10556
rect 9995 -10600 10039 -10556
rect 10095 -10600 10139 -10556
rect 10195 -10600 10239 -10556
rect 10295 -10600 10339 -10556
rect 10395 -10600 10439 -10556
rect 10495 -10600 10539 -10556
rect 10595 -10600 10639 -10556
rect 10695 -10600 10739 -10556
rect 11195 -10600 11239 -10556
rect 11295 -10600 11339 -10556
rect 11395 -10600 11439 -10556
rect 11495 -10600 11539 -10556
rect 11595 -10600 11639 -10556
rect 11695 -10600 11739 -10556
rect 11795 -10600 11839 -10556
rect 11895 -10600 11939 -10556
rect 11995 -10600 12039 -10556
rect 12095 -10600 12139 -10556
rect 12195 -10600 12239 -10556
rect 12295 -10600 12339 -10556
rect 12395 -10600 12439 -10556
rect 12495 -10600 12539 -10556
rect 12595 -10600 12639 -10556
rect 12695 -10600 12739 -10556
rect 13195 -10600 13239 -10556
rect 13295 -10600 13339 -10556
rect 13395 -10600 13439 -10556
rect 13495 -10600 13539 -10556
rect 13595 -10600 13639 -10556
rect 13695 -10600 13739 -10556
rect 13795 -10600 13839 -10556
rect 13895 -10600 13939 -10556
rect 13995 -10600 14039 -10556
rect 14095 -10600 14139 -10556
rect 14195 -10600 14239 -10556
rect 14295 -10600 14339 -10556
rect 14395 -10600 14439 -10556
rect 14495 -10600 14539 -10556
rect 14595 -10600 14639 -10556
rect 14695 -10600 14739 -10556
rect 15195 -10600 15239 -10556
rect 15295 -10600 15339 -10556
rect 15395 -10600 15439 -10556
rect 15495 -10600 15539 -10556
rect 15595 -10600 15639 -10556
rect 15695 -10600 15739 -10556
rect 15795 -10600 15839 -10556
rect 15895 -10600 15939 -10556
rect 15995 -10600 16039 -10556
rect 16095 -10600 16139 -10556
rect 16195 -10600 16239 -10556
rect 16295 -10600 16339 -10556
rect 16395 -10600 16439 -10556
rect 16495 -10600 16539 -10556
rect 16595 -10600 16639 -10556
rect 16695 -10600 16739 -10556
rect 9195 -10700 9239 -10656
rect 9295 -10700 9339 -10656
rect 9395 -10700 9439 -10656
rect 9495 -10700 9539 -10656
rect 9595 -10700 9639 -10656
rect 9695 -10700 9739 -10656
rect 9795 -10700 9839 -10656
rect 9895 -10700 9939 -10656
rect 9995 -10700 10039 -10656
rect 10095 -10700 10139 -10656
rect 10195 -10700 10239 -10656
rect 10295 -10700 10339 -10656
rect 10395 -10700 10439 -10656
rect 10495 -10700 10539 -10656
rect 10595 -10700 10639 -10656
rect 10695 -10700 10739 -10656
rect 11195 -10700 11239 -10656
rect 11295 -10700 11339 -10656
rect 11395 -10700 11439 -10656
rect 11495 -10700 11539 -10656
rect 11595 -10700 11639 -10656
rect 11695 -10700 11739 -10656
rect 11795 -10700 11839 -10656
rect 11895 -10700 11939 -10656
rect 11995 -10700 12039 -10656
rect 12095 -10700 12139 -10656
rect 12195 -10700 12239 -10656
rect 12295 -10700 12339 -10656
rect 12395 -10700 12439 -10656
rect 12495 -10700 12539 -10656
rect 12595 -10700 12639 -10656
rect 12695 -10700 12739 -10656
rect 13195 -10700 13239 -10656
rect 13295 -10700 13339 -10656
rect 13395 -10700 13439 -10656
rect 13495 -10700 13539 -10656
rect 13595 -10700 13639 -10656
rect 13695 -10700 13739 -10656
rect 13795 -10700 13839 -10656
rect 13895 -10700 13939 -10656
rect 13995 -10700 14039 -10656
rect 14095 -10700 14139 -10656
rect 14195 -10700 14239 -10656
rect 14295 -10700 14339 -10656
rect 14395 -10700 14439 -10656
rect 14495 -10700 14539 -10656
rect 14595 -10700 14639 -10656
rect 14695 -10700 14739 -10656
rect 15195 -10700 15239 -10656
rect 15295 -10700 15339 -10656
rect 15395 -10700 15439 -10656
rect 15495 -10700 15539 -10656
rect 15595 -10700 15639 -10656
rect 15695 -10700 15739 -10656
rect 15795 -10700 15839 -10656
rect 15895 -10700 15939 -10656
rect 15995 -10700 16039 -10656
rect 16095 -10700 16139 -10656
rect 16195 -10700 16239 -10656
rect 16295 -10700 16339 -10656
rect 16395 -10700 16439 -10656
rect 16495 -10700 16539 -10656
rect 16595 -10700 16639 -10656
rect 16695 -10700 16739 -10656
rect 9195 -10800 9239 -10756
rect 9295 -10800 9339 -10756
rect 9395 -10800 9439 -10756
rect 9495 -10800 9539 -10756
rect 9595 -10800 9639 -10756
rect 9695 -10800 9739 -10756
rect 9795 -10800 9839 -10756
rect 9895 -10800 9939 -10756
rect 9995 -10800 10039 -10756
rect 10095 -10800 10139 -10756
rect 10195 -10800 10239 -10756
rect 10295 -10800 10339 -10756
rect 10395 -10800 10439 -10756
rect 10495 -10800 10539 -10756
rect 10595 -10800 10639 -10756
rect 10695 -10800 10739 -10756
rect 11195 -10800 11239 -10756
rect 11295 -10800 11339 -10756
rect 11395 -10800 11439 -10756
rect 11495 -10800 11539 -10756
rect 11595 -10800 11639 -10756
rect 11695 -10800 11739 -10756
rect 11795 -10800 11839 -10756
rect 11895 -10800 11939 -10756
rect 11995 -10800 12039 -10756
rect 12095 -10800 12139 -10756
rect 12195 -10800 12239 -10756
rect 12295 -10800 12339 -10756
rect 12395 -10800 12439 -10756
rect 12495 -10800 12539 -10756
rect 12595 -10800 12639 -10756
rect 12695 -10800 12739 -10756
rect 13195 -10800 13239 -10756
rect 13295 -10800 13339 -10756
rect 13395 -10800 13439 -10756
rect 13495 -10800 13539 -10756
rect 13595 -10800 13639 -10756
rect 13695 -10800 13739 -10756
rect 13795 -10800 13839 -10756
rect 13895 -10800 13939 -10756
rect 13995 -10800 14039 -10756
rect 14095 -10800 14139 -10756
rect 14195 -10800 14239 -10756
rect 14295 -10800 14339 -10756
rect 14395 -10800 14439 -10756
rect 14495 -10800 14539 -10756
rect 14595 -10800 14639 -10756
rect 14695 -10800 14739 -10756
rect 15195 -10800 15239 -10756
rect 15295 -10800 15339 -10756
rect 15395 -10800 15439 -10756
rect 15495 -10800 15539 -10756
rect 15595 -10800 15639 -10756
rect 15695 -10800 15739 -10756
rect 15795 -10800 15839 -10756
rect 15895 -10800 15939 -10756
rect 15995 -10800 16039 -10756
rect 16095 -10800 16139 -10756
rect 16195 -10800 16239 -10756
rect 16295 -10800 16339 -10756
rect 16395 -10800 16439 -10756
rect 16495 -10800 16539 -10756
rect 16595 -10800 16639 -10756
rect 16695 -10800 16739 -10756
rect 9195 -10900 9239 -10856
rect 9295 -10900 9339 -10856
rect 9395 -10900 9439 -10856
rect 9495 -10900 9539 -10856
rect 9595 -10900 9639 -10856
rect 9695 -10900 9739 -10856
rect 9795 -10900 9839 -10856
rect 9895 -10900 9939 -10856
rect 9995 -10900 10039 -10856
rect 10095 -10900 10139 -10856
rect 10195 -10900 10239 -10856
rect 10295 -10900 10339 -10856
rect 10395 -10900 10439 -10856
rect 10495 -10900 10539 -10856
rect 10595 -10900 10639 -10856
rect 10695 -10900 10739 -10856
rect 11195 -10900 11239 -10856
rect 11295 -10900 11339 -10856
rect 11395 -10900 11439 -10856
rect 11495 -10900 11539 -10856
rect 11595 -10900 11639 -10856
rect 11695 -10900 11739 -10856
rect 11795 -10900 11839 -10856
rect 11895 -10900 11939 -10856
rect 11995 -10900 12039 -10856
rect 12095 -10900 12139 -10856
rect 12195 -10900 12239 -10856
rect 12295 -10900 12339 -10856
rect 12395 -10900 12439 -10856
rect 12495 -10900 12539 -10856
rect 12595 -10900 12639 -10856
rect 12695 -10900 12739 -10856
rect 13195 -10900 13239 -10856
rect 13295 -10900 13339 -10856
rect 13395 -10900 13439 -10856
rect 13495 -10900 13539 -10856
rect 13595 -10900 13639 -10856
rect 13695 -10900 13739 -10856
rect 13795 -10900 13839 -10856
rect 13895 -10900 13939 -10856
rect 13995 -10900 14039 -10856
rect 14095 -10900 14139 -10856
rect 14195 -10900 14239 -10856
rect 14295 -10900 14339 -10856
rect 14395 -10900 14439 -10856
rect 14495 -10900 14539 -10856
rect 14595 -10900 14639 -10856
rect 14695 -10900 14739 -10856
rect 15195 -10900 15239 -10856
rect 15295 -10900 15339 -10856
rect 15395 -10900 15439 -10856
rect 15495 -10900 15539 -10856
rect 15595 -10900 15639 -10856
rect 15695 -10900 15739 -10856
rect 15795 -10900 15839 -10856
rect 15895 -10900 15939 -10856
rect 15995 -10900 16039 -10856
rect 16095 -10900 16139 -10856
rect 16195 -10900 16239 -10856
rect 16295 -10900 16339 -10856
rect 16395 -10900 16439 -10856
rect 16495 -10900 16539 -10856
rect 16595 -10900 16639 -10856
rect 16695 -10900 16739 -10856
rect 9195 -11000 9239 -10956
rect 9295 -11000 9339 -10956
rect 9395 -11000 9439 -10956
rect 9495 -11000 9539 -10956
rect 9595 -11000 9639 -10956
rect 9695 -11000 9739 -10956
rect 9795 -11000 9839 -10956
rect 9895 -11000 9939 -10956
rect 9995 -11000 10039 -10956
rect 10095 -11000 10139 -10956
rect 10195 -11000 10239 -10956
rect 10295 -11000 10339 -10956
rect 10395 -11000 10439 -10956
rect 10495 -11000 10539 -10956
rect 10595 -11000 10639 -10956
rect 10695 -11000 10739 -10956
rect 11195 -11000 11239 -10956
rect 11295 -11000 11339 -10956
rect 11395 -11000 11439 -10956
rect 11495 -11000 11539 -10956
rect 11595 -11000 11639 -10956
rect 11695 -11000 11739 -10956
rect 11795 -11000 11839 -10956
rect 11895 -11000 11939 -10956
rect 11995 -11000 12039 -10956
rect 12095 -11000 12139 -10956
rect 12195 -11000 12239 -10956
rect 12295 -11000 12339 -10956
rect 12395 -11000 12439 -10956
rect 12495 -11000 12539 -10956
rect 12595 -11000 12639 -10956
rect 12695 -11000 12739 -10956
rect 13195 -11000 13239 -10956
rect 13295 -11000 13339 -10956
rect 13395 -11000 13439 -10956
rect 13495 -11000 13539 -10956
rect 13595 -11000 13639 -10956
rect 13695 -11000 13739 -10956
rect 13795 -11000 13839 -10956
rect 13895 -11000 13939 -10956
rect 13995 -11000 14039 -10956
rect 14095 -11000 14139 -10956
rect 14195 -11000 14239 -10956
rect 14295 -11000 14339 -10956
rect 14395 -11000 14439 -10956
rect 14495 -11000 14539 -10956
rect 14595 -11000 14639 -10956
rect 14695 -11000 14739 -10956
rect 15195 -11000 15239 -10956
rect 15295 -11000 15339 -10956
rect 15395 -11000 15439 -10956
rect 15495 -11000 15539 -10956
rect 15595 -11000 15639 -10956
rect 15695 -11000 15739 -10956
rect 15795 -11000 15839 -10956
rect 15895 -11000 15939 -10956
rect 15995 -11000 16039 -10956
rect 16095 -11000 16139 -10956
rect 16195 -11000 16239 -10956
rect 16295 -11000 16339 -10956
rect 16395 -11000 16439 -10956
rect 16495 -11000 16539 -10956
rect 16595 -11000 16639 -10956
rect 16695 -11000 16739 -10956
rect 9195 -11100 9239 -11056
rect 9295 -11100 9339 -11056
rect 9395 -11100 9439 -11056
rect 9495 -11100 9539 -11056
rect 9595 -11100 9639 -11056
rect 9695 -11100 9739 -11056
rect 9795 -11100 9839 -11056
rect 9895 -11100 9939 -11056
rect 9995 -11100 10039 -11056
rect 10095 -11100 10139 -11056
rect 10195 -11100 10239 -11056
rect 10295 -11100 10339 -11056
rect 10395 -11100 10439 -11056
rect 10495 -11100 10539 -11056
rect 10595 -11100 10639 -11056
rect 10695 -11100 10739 -11056
rect 11195 -11100 11239 -11056
rect 11295 -11100 11339 -11056
rect 11395 -11100 11439 -11056
rect 11495 -11100 11539 -11056
rect 11595 -11100 11639 -11056
rect 11695 -11100 11739 -11056
rect 11795 -11100 11839 -11056
rect 11895 -11100 11939 -11056
rect 11995 -11100 12039 -11056
rect 12095 -11100 12139 -11056
rect 12195 -11100 12239 -11056
rect 12295 -11100 12339 -11056
rect 12395 -11100 12439 -11056
rect 12495 -11100 12539 -11056
rect 12595 -11100 12639 -11056
rect 12695 -11100 12739 -11056
rect 13195 -11100 13239 -11056
rect 13295 -11100 13339 -11056
rect 13395 -11100 13439 -11056
rect 13495 -11100 13539 -11056
rect 13595 -11100 13639 -11056
rect 13695 -11100 13739 -11056
rect 13795 -11100 13839 -11056
rect 13895 -11100 13939 -11056
rect 13995 -11100 14039 -11056
rect 14095 -11100 14139 -11056
rect 14195 -11100 14239 -11056
rect 14295 -11100 14339 -11056
rect 14395 -11100 14439 -11056
rect 14495 -11100 14539 -11056
rect 14595 -11100 14639 -11056
rect 14695 -11100 14739 -11056
rect 15195 -11100 15239 -11056
rect 15295 -11100 15339 -11056
rect 15395 -11100 15439 -11056
rect 15495 -11100 15539 -11056
rect 15595 -11100 15639 -11056
rect 15695 -11100 15739 -11056
rect 15795 -11100 15839 -11056
rect 15895 -11100 15939 -11056
rect 15995 -11100 16039 -11056
rect 16095 -11100 16139 -11056
rect 16195 -11100 16239 -11056
rect 16295 -11100 16339 -11056
rect 16395 -11100 16439 -11056
rect 16495 -11100 16539 -11056
rect 16595 -11100 16639 -11056
rect 16695 -11100 16739 -11056
rect 9195 -11200 9239 -11156
rect 9295 -11200 9339 -11156
rect 9395 -11200 9439 -11156
rect 9495 -11200 9539 -11156
rect 9595 -11200 9639 -11156
rect 9695 -11200 9739 -11156
rect 9795 -11200 9839 -11156
rect 9895 -11200 9939 -11156
rect 9995 -11200 10039 -11156
rect 10095 -11200 10139 -11156
rect 10195 -11200 10239 -11156
rect 10295 -11200 10339 -11156
rect 10395 -11200 10439 -11156
rect 10495 -11200 10539 -11156
rect 10595 -11200 10639 -11156
rect 10695 -11200 10739 -11156
rect 11195 -11200 11239 -11156
rect 11295 -11200 11339 -11156
rect 11395 -11200 11439 -11156
rect 11495 -11200 11539 -11156
rect 11595 -11200 11639 -11156
rect 11695 -11200 11739 -11156
rect 11795 -11200 11839 -11156
rect 11895 -11200 11939 -11156
rect 11995 -11200 12039 -11156
rect 12095 -11200 12139 -11156
rect 12195 -11200 12239 -11156
rect 12295 -11200 12339 -11156
rect 12395 -11200 12439 -11156
rect 12495 -11200 12539 -11156
rect 12595 -11200 12639 -11156
rect 12695 -11200 12739 -11156
rect 13195 -11200 13239 -11156
rect 13295 -11200 13339 -11156
rect 13395 -11200 13439 -11156
rect 13495 -11200 13539 -11156
rect 13595 -11200 13639 -11156
rect 13695 -11200 13739 -11156
rect 13795 -11200 13839 -11156
rect 13895 -11200 13939 -11156
rect 13995 -11200 14039 -11156
rect 14095 -11200 14139 -11156
rect 14195 -11200 14239 -11156
rect 14295 -11200 14339 -11156
rect 14395 -11200 14439 -11156
rect 14495 -11200 14539 -11156
rect 14595 -11200 14639 -11156
rect 14695 -11200 14739 -11156
rect 15195 -11200 15239 -11156
rect 15295 -11200 15339 -11156
rect 15395 -11200 15439 -11156
rect 15495 -11200 15539 -11156
rect 15595 -11200 15639 -11156
rect 15695 -11200 15739 -11156
rect 15795 -11200 15839 -11156
rect 15895 -11200 15939 -11156
rect 15995 -11200 16039 -11156
rect 16095 -11200 16139 -11156
rect 16195 -11200 16239 -11156
rect 16295 -11200 16339 -11156
rect 16395 -11200 16439 -11156
rect 16495 -11200 16539 -11156
rect 16595 -11200 16639 -11156
rect 16695 -11200 16739 -11156
rect 9195 -11300 9239 -11256
rect 9295 -11300 9339 -11256
rect 9395 -11300 9439 -11256
rect 9495 -11300 9539 -11256
rect 9595 -11300 9639 -11256
rect 9695 -11300 9739 -11256
rect 9795 -11300 9839 -11256
rect 9895 -11300 9939 -11256
rect 9995 -11300 10039 -11256
rect 10095 -11300 10139 -11256
rect 10195 -11300 10239 -11256
rect 10295 -11300 10339 -11256
rect 10395 -11300 10439 -11256
rect 10495 -11300 10539 -11256
rect 10595 -11300 10639 -11256
rect 10695 -11300 10739 -11256
rect 11195 -11300 11239 -11256
rect 11295 -11300 11339 -11256
rect 11395 -11300 11439 -11256
rect 11495 -11300 11539 -11256
rect 11595 -11300 11639 -11256
rect 11695 -11300 11739 -11256
rect 11795 -11300 11839 -11256
rect 11895 -11300 11939 -11256
rect 11995 -11300 12039 -11256
rect 12095 -11300 12139 -11256
rect 12195 -11300 12239 -11256
rect 12295 -11300 12339 -11256
rect 12395 -11300 12439 -11256
rect 12495 -11300 12539 -11256
rect 12595 -11300 12639 -11256
rect 12695 -11300 12739 -11256
rect 13195 -11300 13239 -11256
rect 13295 -11300 13339 -11256
rect 13395 -11300 13439 -11256
rect 13495 -11300 13539 -11256
rect 13595 -11300 13639 -11256
rect 13695 -11300 13739 -11256
rect 13795 -11300 13839 -11256
rect 13895 -11300 13939 -11256
rect 13995 -11300 14039 -11256
rect 14095 -11300 14139 -11256
rect 14195 -11300 14239 -11256
rect 14295 -11300 14339 -11256
rect 14395 -11300 14439 -11256
rect 14495 -11300 14539 -11256
rect 14595 -11300 14639 -11256
rect 14695 -11300 14739 -11256
rect 15195 -11300 15239 -11256
rect 15295 -11300 15339 -11256
rect 15395 -11300 15439 -11256
rect 15495 -11300 15539 -11256
rect 15595 -11300 15639 -11256
rect 15695 -11300 15739 -11256
rect 15795 -11300 15839 -11256
rect 15895 -11300 15939 -11256
rect 15995 -11300 16039 -11256
rect 16095 -11300 16139 -11256
rect 16195 -11300 16239 -11256
rect 16295 -11300 16339 -11256
rect 16395 -11300 16439 -11256
rect 16495 -11300 16539 -11256
rect 16595 -11300 16639 -11256
rect 16695 -11300 16739 -11256
rect 37223 -9682 37267 -9638
rect 37323 -9682 37367 -9638
rect 37423 -9682 37467 -9638
rect 37523 -9682 37567 -9638
rect 37623 -9682 37667 -9638
rect 37723 -9682 37767 -9638
rect 37823 -9682 37867 -9638
rect 37923 -9682 37967 -9638
rect 38023 -9682 38067 -9638
rect 38123 -9682 38167 -9638
rect 38223 -9682 38267 -9638
rect 38323 -9682 38367 -9638
rect 38423 -9682 38467 -9638
rect 38523 -9682 38567 -9638
rect 38623 -9682 38667 -9638
rect 38723 -9682 38767 -9638
rect 39223 -9682 39267 -9638
rect 39323 -9682 39367 -9638
rect 39423 -9682 39467 -9638
rect 39523 -9682 39567 -9638
rect 39623 -9682 39667 -9638
rect 39723 -9682 39767 -9638
rect 39823 -9682 39867 -9638
rect 39923 -9682 39967 -9638
rect 40023 -9682 40067 -9638
rect 40123 -9682 40167 -9638
rect 40223 -9682 40267 -9638
rect 40323 -9682 40367 -9638
rect 40423 -9682 40467 -9638
rect 40523 -9682 40567 -9638
rect 40623 -9682 40667 -9638
rect 40723 -9682 40767 -9638
rect 41223 -9682 41267 -9638
rect 41323 -9682 41367 -9638
rect 41423 -9682 41467 -9638
rect 41523 -9682 41567 -9638
rect 41623 -9682 41667 -9638
rect 41723 -9682 41767 -9638
rect 41823 -9682 41867 -9638
rect 41923 -9682 41967 -9638
rect 42023 -9682 42067 -9638
rect 42123 -9682 42167 -9638
rect 42223 -9682 42267 -9638
rect 42323 -9682 42367 -9638
rect 42423 -9682 42467 -9638
rect 42523 -9682 42567 -9638
rect 42623 -9682 42667 -9638
rect 42723 -9682 42767 -9638
rect 43223 -9682 43267 -9638
rect 43323 -9682 43367 -9638
rect 43423 -9682 43467 -9638
rect 43523 -9682 43567 -9638
rect 43623 -9682 43667 -9638
rect 43723 -9682 43767 -9638
rect 43823 -9682 43867 -9638
rect 43923 -9682 43967 -9638
rect 44023 -9682 44067 -9638
rect 44123 -9682 44167 -9638
rect 44223 -9682 44267 -9638
rect 44323 -9682 44367 -9638
rect 44423 -9682 44467 -9638
rect 44523 -9682 44567 -9638
rect 44623 -9682 44667 -9638
rect 44723 -9682 44767 -9638
rect 37223 -9782 37267 -9738
rect 37323 -9782 37367 -9738
rect 37423 -9782 37467 -9738
rect 37523 -9782 37567 -9738
rect 37623 -9782 37667 -9738
rect 37723 -9782 37767 -9738
rect 37823 -9782 37867 -9738
rect 37923 -9782 37967 -9738
rect 38023 -9782 38067 -9738
rect 38123 -9782 38167 -9738
rect 38223 -9782 38267 -9738
rect 38323 -9782 38367 -9738
rect 38423 -9782 38467 -9738
rect 38523 -9782 38567 -9738
rect 38623 -9782 38667 -9738
rect 38723 -9782 38767 -9738
rect 39223 -9782 39267 -9738
rect 39323 -9782 39367 -9738
rect 39423 -9782 39467 -9738
rect 39523 -9782 39567 -9738
rect 39623 -9782 39667 -9738
rect 39723 -9782 39767 -9738
rect 39823 -9782 39867 -9738
rect 39923 -9782 39967 -9738
rect 40023 -9782 40067 -9738
rect 40123 -9782 40167 -9738
rect 40223 -9782 40267 -9738
rect 40323 -9782 40367 -9738
rect 40423 -9782 40467 -9738
rect 40523 -9782 40567 -9738
rect 40623 -9782 40667 -9738
rect 40723 -9782 40767 -9738
rect 41223 -9782 41267 -9738
rect 41323 -9782 41367 -9738
rect 41423 -9782 41467 -9738
rect 41523 -9782 41567 -9738
rect 41623 -9782 41667 -9738
rect 41723 -9782 41767 -9738
rect 41823 -9782 41867 -9738
rect 41923 -9782 41967 -9738
rect 42023 -9782 42067 -9738
rect 42123 -9782 42167 -9738
rect 42223 -9782 42267 -9738
rect 42323 -9782 42367 -9738
rect 42423 -9782 42467 -9738
rect 42523 -9782 42567 -9738
rect 42623 -9782 42667 -9738
rect 42723 -9782 42767 -9738
rect 43223 -9782 43267 -9738
rect 43323 -9782 43367 -9738
rect 43423 -9782 43467 -9738
rect 43523 -9782 43567 -9738
rect 43623 -9782 43667 -9738
rect 43723 -9782 43767 -9738
rect 43823 -9782 43867 -9738
rect 43923 -9782 43967 -9738
rect 44023 -9782 44067 -9738
rect 44123 -9782 44167 -9738
rect 44223 -9782 44267 -9738
rect 44323 -9782 44367 -9738
rect 44423 -9782 44467 -9738
rect 44523 -9782 44567 -9738
rect 44623 -9782 44667 -9738
rect 44723 -9782 44767 -9738
rect 37223 -9882 37267 -9838
rect 37323 -9882 37367 -9838
rect 37423 -9882 37467 -9838
rect 37523 -9882 37567 -9838
rect 37623 -9882 37667 -9838
rect 37723 -9882 37767 -9838
rect 37823 -9882 37867 -9838
rect 37923 -9882 37967 -9838
rect 38023 -9882 38067 -9838
rect 38123 -9882 38167 -9838
rect 38223 -9882 38267 -9838
rect 38323 -9882 38367 -9838
rect 38423 -9882 38467 -9838
rect 38523 -9882 38567 -9838
rect 38623 -9882 38667 -9838
rect 38723 -9882 38767 -9838
rect 39223 -9882 39267 -9838
rect 39323 -9882 39367 -9838
rect 39423 -9882 39467 -9838
rect 39523 -9882 39567 -9838
rect 39623 -9882 39667 -9838
rect 39723 -9882 39767 -9838
rect 39823 -9882 39867 -9838
rect 39923 -9882 39967 -9838
rect 40023 -9882 40067 -9838
rect 40123 -9882 40167 -9838
rect 40223 -9882 40267 -9838
rect 40323 -9882 40367 -9838
rect 40423 -9882 40467 -9838
rect 40523 -9882 40567 -9838
rect 40623 -9882 40667 -9838
rect 40723 -9882 40767 -9838
rect 41223 -9882 41267 -9838
rect 41323 -9882 41367 -9838
rect 41423 -9882 41467 -9838
rect 41523 -9882 41567 -9838
rect 41623 -9882 41667 -9838
rect 41723 -9882 41767 -9838
rect 41823 -9882 41867 -9838
rect 41923 -9882 41967 -9838
rect 42023 -9882 42067 -9838
rect 42123 -9882 42167 -9838
rect 42223 -9882 42267 -9838
rect 42323 -9882 42367 -9838
rect 42423 -9882 42467 -9838
rect 42523 -9882 42567 -9838
rect 42623 -9882 42667 -9838
rect 42723 -9882 42767 -9838
rect 43223 -9882 43267 -9838
rect 43323 -9882 43367 -9838
rect 43423 -9882 43467 -9838
rect 43523 -9882 43567 -9838
rect 43623 -9882 43667 -9838
rect 43723 -9882 43767 -9838
rect 43823 -9882 43867 -9838
rect 43923 -9882 43967 -9838
rect 44023 -9882 44067 -9838
rect 44123 -9882 44167 -9838
rect 44223 -9882 44267 -9838
rect 44323 -9882 44367 -9838
rect 44423 -9882 44467 -9838
rect 44523 -9882 44567 -9838
rect 44623 -9882 44667 -9838
rect 44723 -9882 44767 -9838
rect 37223 -9982 37267 -9938
rect 37323 -9982 37367 -9938
rect 37423 -9982 37467 -9938
rect 37523 -9982 37567 -9938
rect 37623 -9982 37667 -9938
rect 37723 -9982 37767 -9938
rect 37823 -9982 37867 -9938
rect 37923 -9982 37967 -9938
rect 38023 -9982 38067 -9938
rect 38123 -9982 38167 -9938
rect 38223 -9982 38267 -9938
rect 38323 -9982 38367 -9938
rect 38423 -9982 38467 -9938
rect 38523 -9982 38567 -9938
rect 38623 -9982 38667 -9938
rect 38723 -9982 38767 -9938
rect 39223 -9982 39267 -9938
rect 39323 -9982 39367 -9938
rect 39423 -9982 39467 -9938
rect 39523 -9982 39567 -9938
rect 39623 -9982 39667 -9938
rect 39723 -9982 39767 -9938
rect 39823 -9982 39867 -9938
rect 39923 -9982 39967 -9938
rect 40023 -9982 40067 -9938
rect 40123 -9982 40167 -9938
rect 40223 -9982 40267 -9938
rect 40323 -9982 40367 -9938
rect 40423 -9982 40467 -9938
rect 40523 -9982 40567 -9938
rect 40623 -9982 40667 -9938
rect 40723 -9982 40767 -9938
rect 41223 -9982 41267 -9938
rect 41323 -9982 41367 -9938
rect 41423 -9982 41467 -9938
rect 41523 -9982 41567 -9938
rect 41623 -9982 41667 -9938
rect 41723 -9982 41767 -9938
rect 41823 -9982 41867 -9938
rect 41923 -9982 41967 -9938
rect 42023 -9982 42067 -9938
rect 42123 -9982 42167 -9938
rect 42223 -9982 42267 -9938
rect 42323 -9982 42367 -9938
rect 42423 -9982 42467 -9938
rect 42523 -9982 42567 -9938
rect 42623 -9982 42667 -9938
rect 42723 -9982 42767 -9938
rect 43223 -9982 43267 -9938
rect 43323 -9982 43367 -9938
rect 43423 -9982 43467 -9938
rect 43523 -9982 43567 -9938
rect 43623 -9982 43667 -9938
rect 43723 -9982 43767 -9938
rect 43823 -9982 43867 -9938
rect 43923 -9982 43967 -9938
rect 44023 -9982 44067 -9938
rect 44123 -9982 44167 -9938
rect 44223 -9982 44267 -9938
rect 44323 -9982 44367 -9938
rect 44423 -9982 44467 -9938
rect 44523 -9982 44567 -9938
rect 44623 -9982 44667 -9938
rect 44723 -9982 44767 -9938
rect 37223 -10082 37267 -10038
rect 37323 -10082 37367 -10038
rect 37423 -10082 37467 -10038
rect 37523 -10082 37567 -10038
rect 37623 -10082 37667 -10038
rect 37723 -10082 37767 -10038
rect 37823 -10082 37867 -10038
rect 37923 -10082 37967 -10038
rect 38023 -10082 38067 -10038
rect 38123 -10082 38167 -10038
rect 38223 -10082 38267 -10038
rect 38323 -10082 38367 -10038
rect 38423 -10082 38467 -10038
rect 38523 -10082 38567 -10038
rect 38623 -10082 38667 -10038
rect 38723 -10082 38767 -10038
rect 39223 -10082 39267 -10038
rect 39323 -10082 39367 -10038
rect 39423 -10082 39467 -10038
rect 39523 -10082 39567 -10038
rect 39623 -10082 39667 -10038
rect 39723 -10082 39767 -10038
rect 39823 -10082 39867 -10038
rect 39923 -10082 39967 -10038
rect 40023 -10082 40067 -10038
rect 40123 -10082 40167 -10038
rect 40223 -10082 40267 -10038
rect 40323 -10082 40367 -10038
rect 40423 -10082 40467 -10038
rect 40523 -10082 40567 -10038
rect 40623 -10082 40667 -10038
rect 40723 -10082 40767 -10038
rect 41223 -10082 41267 -10038
rect 41323 -10082 41367 -10038
rect 41423 -10082 41467 -10038
rect 41523 -10082 41567 -10038
rect 41623 -10082 41667 -10038
rect 41723 -10082 41767 -10038
rect 41823 -10082 41867 -10038
rect 41923 -10082 41967 -10038
rect 42023 -10082 42067 -10038
rect 42123 -10082 42167 -10038
rect 42223 -10082 42267 -10038
rect 42323 -10082 42367 -10038
rect 42423 -10082 42467 -10038
rect 42523 -10082 42567 -10038
rect 42623 -10082 42667 -10038
rect 42723 -10082 42767 -10038
rect 43223 -10082 43267 -10038
rect 43323 -10082 43367 -10038
rect 43423 -10082 43467 -10038
rect 43523 -10082 43567 -10038
rect 43623 -10082 43667 -10038
rect 43723 -10082 43767 -10038
rect 43823 -10082 43867 -10038
rect 43923 -10082 43967 -10038
rect 44023 -10082 44067 -10038
rect 44123 -10082 44167 -10038
rect 44223 -10082 44267 -10038
rect 44323 -10082 44367 -10038
rect 44423 -10082 44467 -10038
rect 44523 -10082 44567 -10038
rect 44623 -10082 44667 -10038
rect 44723 -10082 44767 -10038
rect 37223 -10182 37267 -10138
rect 37323 -10182 37367 -10138
rect 37423 -10182 37467 -10138
rect 37523 -10182 37567 -10138
rect 37623 -10182 37667 -10138
rect 37723 -10182 37767 -10138
rect 37823 -10182 37867 -10138
rect 37923 -10182 37967 -10138
rect 38023 -10182 38067 -10138
rect 38123 -10182 38167 -10138
rect 38223 -10182 38267 -10138
rect 38323 -10182 38367 -10138
rect 38423 -10182 38467 -10138
rect 38523 -10182 38567 -10138
rect 38623 -10182 38667 -10138
rect 38723 -10182 38767 -10138
rect 39223 -10182 39267 -10138
rect 39323 -10182 39367 -10138
rect 39423 -10182 39467 -10138
rect 39523 -10182 39567 -10138
rect 39623 -10182 39667 -10138
rect 39723 -10182 39767 -10138
rect 39823 -10182 39867 -10138
rect 39923 -10182 39967 -10138
rect 40023 -10182 40067 -10138
rect 40123 -10182 40167 -10138
rect 40223 -10182 40267 -10138
rect 40323 -10182 40367 -10138
rect 40423 -10182 40467 -10138
rect 40523 -10182 40567 -10138
rect 40623 -10182 40667 -10138
rect 40723 -10182 40767 -10138
rect 41223 -10182 41267 -10138
rect 41323 -10182 41367 -10138
rect 41423 -10182 41467 -10138
rect 41523 -10182 41567 -10138
rect 41623 -10182 41667 -10138
rect 41723 -10182 41767 -10138
rect 41823 -10182 41867 -10138
rect 41923 -10182 41967 -10138
rect 42023 -10182 42067 -10138
rect 42123 -10182 42167 -10138
rect 42223 -10182 42267 -10138
rect 42323 -10182 42367 -10138
rect 42423 -10182 42467 -10138
rect 42523 -10182 42567 -10138
rect 42623 -10182 42667 -10138
rect 42723 -10182 42767 -10138
rect 43223 -10182 43267 -10138
rect 43323 -10182 43367 -10138
rect 43423 -10182 43467 -10138
rect 43523 -10182 43567 -10138
rect 43623 -10182 43667 -10138
rect 43723 -10182 43767 -10138
rect 43823 -10182 43867 -10138
rect 43923 -10182 43967 -10138
rect 44023 -10182 44067 -10138
rect 44123 -10182 44167 -10138
rect 44223 -10182 44267 -10138
rect 44323 -10182 44367 -10138
rect 44423 -10182 44467 -10138
rect 44523 -10182 44567 -10138
rect 44623 -10182 44667 -10138
rect 44723 -10182 44767 -10138
rect 37223 -10282 37267 -10238
rect 37323 -10282 37367 -10238
rect 37423 -10282 37467 -10238
rect 37523 -10282 37567 -10238
rect 37623 -10282 37667 -10238
rect 37723 -10282 37767 -10238
rect 37823 -10282 37867 -10238
rect 37923 -10282 37967 -10238
rect 38023 -10282 38067 -10238
rect 38123 -10282 38167 -10238
rect 38223 -10282 38267 -10238
rect 38323 -10282 38367 -10238
rect 38423 -10282 38467 -10238
rect 38523 -10282 38567 -10238
rect 38623 -10282 38667 -10238
rect 38723 -10282 38767 -10238
rect 39223 -10282 39267 -10238
rect 39323 -10282 39367 -10238
rect 39423 -10282 39467 -10238
rect 39523 -10282 39567 -10238
rect 39623 -10282 39667 -10238
rect 39723 -10282 39767 -10238
rect 39823 -10282 39867 -10238
rect 39923 -10282 39967 -10238
rect 40023 -10282 40067 -10238
rect 40123 -10282 40167 -10238
rect 40223 -10282 40267 -10238
rect 40323 -10282 40367 -10238
rect 40423 -10282 40467 -10238
rect 40523 -10282 40567 -10238
rect 40623 -10282 40667 -10238
rect 40723 -10282 40767 -10238
rect 41223 -10282 41267 -10238
rect 41323 -10282 41367 -10238
rect 41423 -10282 41467 -10238
rect 41523 -10282 41567 -10238
rect 41623 -10282 41667 -10238
rect 41723 -10282 41767 -10238
rect 41823 -10282 41867 -10238
rect 41923 -10282 41967 -10238
rect 42023 -10282 42067 -10238
rect 42123 -10282 42167 -10238
rect 42223 -10282 42267 -10238
rect 42323 -10282 42367 -10238
rect 42423 -10282 42467 -10238
rect 42523 -10282 42567 -10238
rect 42623 -10282 42667 -10238
rect 42723 -10282 42767 -10238
rect 43223 -10282 43267 -10238
rect 43323 -10282 43367 -10238
rect 43423 -10282 43467 -10238
rect 43523 -10282 43567 -10238
rect 43623 -10282 43667 -10238
rect 43723 -10282 43767 -10238
rect 43823 -10282 43867 -10238
rect 43923 -10282 43967 -10238
rect 44023 -10282 44067 -10238
rect 44123 -10282 44167 -10238
rect 44223 -10282 44267 -10238
rect 44323 -10282 44367 -10238
rect 44423 -10282 44467 -10238
rect 44523 -10282 44567 -10238
rect 44623 -10282 44667 -10238
rect 44723 -10282 44767 -10238
rect 37223 -10382 37267 -10338
rect 37323 -10382 37367 -10338
rect 37423 -10382 37467 -10338
rect 37523 -10382 37567 -10338
rect 37623 -10382 37667 -10338
rect 37723 -10382 37767 -10338
rect 37823 -10382 37867 -10338
rect 37923 -10382 37967 -10338
rect 38023 -10382 38067 -10338
rect 38123 -10382 38167 -10338
rect 38223 -10382 38267 -10338
rect 38323 -10382 38367 -10338
rect 38423 -10382 38467 -10338
rect 38523 -10382 38567 -10338
rect 38623 -10382 38667 -10338
rect 38723 -10382 38767 -10338
rect 39223 -10382 39267 -10338
rect 39323 -10382 39367 -10338
rect 39423 -10382 39467 -10338
rect 39523 -10382 39567 -10338
rect 39623 -10382 39667 -10338
rect 39723 -10382 39767 -10338
rect 39823 -10382 39867 -10338
rect 39923 -10382 39967 -10338
rect 40023 -10382 40067 -10338
rect 40123 -10382 40167 -10338
rect 40223 -10382 40267 -10338
rect 40323 -10382 40367 -10338
rect 40423 -10382 40467 -10338
rect 40523 -10382 40567 -10338
rect 40623 -10382 40667 -10338
rect 40723 -10382 40767 -10338
rect 41223 -10382 41267 -10338
rect 41323 -10382 41367 -10338
rect 41423 -10382 41467 -10338
rect 41523 -10382 41567 -10338
rect 41623 -10382 41667 -10338
rect 41723 -10382 41767 -10338
rect 41823 -10382 41867 -10338
rect 41923 -10382 41967 -10338
rect 42023 -10382 42067 -10338
rect 42123 -10382 42167 -10338
rect 42223 -10382 42267 -10338
rect 42323 -10382 42367 -10338
rect 42423 -10382 42467 -10338
rect 42523 -10382 42567 -10338
rect 42623 -10382 42667 -10338
rect 42723 -10382 42767 -10338
rect 43223 -10382 43267 -10338
rect 43323 -10382 43367 -10338
rect 43423 -10382 43467 -10338
rect 43523 -10382 43567 -10338
rect 43623 -10382 43667 -10338
rect 43723 -10382 43767 -10338
rect 43823 -10382 43867 -10338
rect 43923 -10382 43967 -10338
rect 44023 -10382 44067 -10338
rect 44123 -10382 44167 -10338
rect 44223 -10382 44267 -10338
rect 44323 -10382 44367 -10338
rect 44423 -10382 44467 -10338
rect 44523 -10382 44567 -10338
rect 44623 -10382 44667 -10338
rect 44723 -10382 44767 -10338
rect 37223 -10482 37267 -10438
rect 37323 -10482 37367 -10438
rect 37423 -10482 37467 -10438
rect 37523 -10482 37567 -10438
rect 37623 -10482 37667 -10438
rect 37723 -10482 37767 -10438
rect 37823 -10482 37867 -10438
rect 37923 -10482 37967 -10438
rect 38023 -10482 38067 -10438
rect 38123 -10482 38167 -10438
rect 38223 -10482 38267 -10438
rect 38323 -10482 38367 -10438
rect 38423 -10482 38467 -10438
rect 38523 -10482 38567 -10438
rect 38623 -10482 38667 -10438
rect 38723 -10482 38767 -10438
rect 39223 -10482 39267 -10438
rect 39323 -10482 39367 -10438
rect 39423 -10482 39467 -10438
rect 39523 -10482 39567 -10438
rect 39623 -10482 39667 -10438
rect 39723 -10482 39767 -10438
rect 39823 -10482 39867 -10438
rect 39923 -10482 39967 -10438
rect 40023 -10482 40067 -10438
rect 40123 -10482 40167 -10438
rect 40223 -10482 40267 -10438
rect 40323 -10482 40367 -10438
rect 40423 -10482 40467 -10438
rect 40523 -10482 40567 -10438
rect 40623 -10482 40667 -10438
rect 40723 -10482 40767 -10438
rect 41223 -10482 41267 -10438
rect 41323 -10482 41367 -10438
rect 41423 -10482 41467 -10438
rect 41523 -10482 41567 -10438
rect 41623 -10482 41667 -10438
rect 41723 -10482 41767 -10438
rect 41823 -10482 41867 -10438
rect 41923 -10482 41967 -10438
rect 42023 -10482 42067 -10438
rect 42123 -10482 42167 -10438
rect 42223 -10482 42267 -10438
rect 42323 -10482 42367 -10438
rect 42423 -10482 42467 -10438
rect 42523 -10482 42567 -10438
rect 42623 -10482 42667 -10438
rect 42723 -10482 42767 -10438
rect 43223 -10482 43267 -10438
rect 43323 -10482 43367 -10438
rect 43423 -10482 43467 -10438
rect 43523 -10482 43567 -10438
rect 43623 -10482 43667 -10438
rect 43723 -10482 43767 -10438
rect 43823 -10482 43867 -10438
rect 43923 -10482 43967 -10438
rect 44023 -10482 44067 -10438
rect 44123 -10482 44167 -10438
rect 44223 -10482 44267 -10438
rect 44323 -10482 44367 -10438
rect 44423 -10482 44467 -10438
rect 44523 -10482 44567 -10438
rect 44623 -10482 44667 -10438
rect 44723 -10482 44767 -10438
rect 37223 -10582 37267 -10538
rect 37323 -10582 37367 -10538
rect 37423 -10582 37467 -10538
rect 37523 -10582 37567 -10538
rect 37623 -10582 37667 -10538
rect 37723 -10582 37767 -10538
rect 37823 -10582 37867 -10538
rect 37923 -10582 37967 -10538
rect 38023 -10582 38067 -10538
rect 38123 -10582 38167 -10538
rect 38223 -10582 38267 -10538
rect 38323 -10582 38367 -10538
rect 38423 -10582 38467 -10538
rect 38523 -10582 38567 -10538
rect 38623 -10582 38667 -10538
rect 38723 -10582 38767 -10538
rect 39223 -10582 39267 -10538
rect 39323 -10582 39367 -10538
rect 39423 -10582 39467 -10538
rect 39523 -10582 39567 -10538
rect 39623 -10582 39667 -10538
rect 39723 -10582 39767 -10538
rect 39823 -10582 39867 -10538
rect 39923 -10582 39967 -10538
rect 40023 -10582 40067 -10538
rect 40123 -10582 40167 -10538
rect 40223 -10582 40267 -10538
rect 40323 -10582 40367 -10538
rect 40423 -10582 40467 -10538
rect 40523 -10582 40567 -10538
rect 40623 -10582 40667 -10538
rect 40723 -10582 40767 -10538
rect 41223 -10582 41267 -10538
rect 41323 -10582 41367 -10538
rect 41423 -10582 41467 -10538
rect 41523 -10582 41567 -10538
rect 41623 -10582 41667 -10538
rect 41723 -10582 41767 -10538
rect 41823 -10582 41867 -10538
rect 41923 -10582 41967 -10538
rect 42023 -10582 42067 -10538
rect 42123 -10582 42167 -10538
rect 42223 -10582 42267 -10538
rect 42323 -10582 42367 -10538
rect 42423 -10582 42467 -10538
rect 42523 -10582 42567 -10538
rect 42623 -10582 42667 -10538
rect 42723 -10582 42767 -10538
rect 43223 -10582 43267 -10538
rect 43323 -10582 43367 -10538
rect 43423 -10582 43467 -10538
rect 43523 -10582 43567 -10538
rect 43623 -10582 43667 -10538
rect 43723 -10582 43767 -10538
rect 43823 -10582 43867 -10538
rect 43923 -10582 43967 -10538
rect 44023 -10582 44067 -10538
rect 44123 -10582 44167 -10538
rect 44223 -10582 44267 -10538
rect 44323 -10582 44367 -10538
rect 44423 -10582 44467 -10538
rect 44523 -10582 44567 -10538
rect 44623 -10582 44667 -10538
rect 44723 -10582 44767 -10538
rect 37223 -10682 37267 -10638
rect 37323 -10682 37367 -10638
rect 37423 -10682 37467 -10638
rect 37523 -10682 37567 -10638
rect 37623 -10682 37667 -10638
rect 37723 -10682 37767 -10638
rect 37823 -10682 37867 -10638
rect 37923 -10682 37967 -10638
rect 38023 -10682 38067 -10638
rect 38123 -10682 38167 -10638
rect 38223 -10682 38267 -10638
rect 38323 -10682 38367 -10638
rect 38423 -10682 38467 -10638
rect 38523 -10682 38567 -10638
rect 38623 -10682 38667 -10638
rect 38723 -10682 38767 -10638
rect 39223 -10682 39267 -10638
rect 39323 -10682 39367 -10638
rect 39423 -10682 39467 -10638
rect 39523 -10682 39567 -10638
rect 39623 -10682 39667 -10638
rect 39723 -10682 39767 -10638
rect 39823 -10682 39867 -10638
rect 39923 -10682 39967 -10638
rect 40023 -10682 40067 -10638
rect 40123 -10682 40167 -10638
rect 40223 -10682 40267 -10638
rect 40323 -10682 40367 -10638
rect 40423 -10682 40467 -10638
rect 40523 -10682 40567 -10638
rect 40623 -10682 40667 -10638
rect 40723 -10682 40767 -10638
rect 41223 -10682 41267 -10638
rect 41323 -10682 41367 -10638
rect 41423 -10682 41467 -10638
rect 41523 -10682 41567 -10638
rect 41623 -10682 41667 -10638
rect 41723 -10682 41767 -10638
rect 41823 -10682 41867 -10638
rect 41923 -10682 41967 -10638
rect 42023 -10682 42067 -10638
rect 42123 -10682 42167 -10638
rect 42223 -10682 42267 -10638
rect 42323 -10682 42367 -10638
rect 42423 -10682 42467 -10638
rect 42523 -10682 42567 -10638
rect 42623 -10682 42667 -10638
rect 42723 -10682 42767 -10638
rect 43223 -10682 43267 -10638
rect 43323 -10682 43367 -10638
rect 43423 -10682 43467 -10638
rect 43523 -10682 43567 -10638
rect 43623 -10682 43667 -10638
rect 43723 -10682 43767 -10638
rect 43823 -10682 43867 -10638
rect 43923 -10682 43967 -10638
rect 44023 -10682 44067 -10638
rect 44123 -10682 44167 -10638
rect 44223 -10682 44267 -10638
rect 44323 -10682 44367 -10638
rect 44423 -10682 44467 -10638
rect 44523 -10682 44567 -10638
rect 44623 -10682 44667 -10638
rect 44723 -10682 44767 -10638
rect 37223 -10782 37267 -10738
rect 37323 -10782 37367 -10738
rect 37423 -10782 37467 -10738
rect 37523 -10782 37567 -10738
rect 37623 -10782 37667 -10738
rect 37723 -10782 37767 -10738
rect 37823 -10782 37867 -10738
rect 37923 -10782 37967 -10738
rect 38023 -10782 38067 -10738
rect 38123 -10782 38167 -10738
rect 38223 -10782 38267 -10738
rect 38323 -10782 38367 -10738
rect 38423 -10782 38467 -10738
rect 38523 -10782 38567 -10738
rect 38623 -10782 38667 -10738
rect 38723 -10782 38767 -10738
rect 39223 -10782 39267 -10738
rect 39323 -10782 39367 -10738
rect 39423 -10782 39467 -10738
rect 39523 -10782 39567 -10738
rect 39623 -10782 39667 -10738
rect 39723 -10782 39767 -10738
rect 39823 -10782 39867 -10738
rect 39923 -10782 39967 -10738
rect 40023 -10782 40067 -10738
rect 40123 -10782 40167 -10738
rect 40223 -10782 40267 -10738
rect 40323 -10782 40367 -10738
rect 40423 -10782 40467 -10738
rect 40523 -10782 40567 -10738
rect 40623 -10782 40667 -10738
rect 40723 -10782 40767 -10738
rect 41223 -10782 41267 -10738
rect 41323 -10782 41367 -10738
rect 41423 -10782 41467 -10738
rect 41523 -10782 41567 -10738
rect 41623 -10782 41667 -10738
rect 41723 -10782 41767 -10738
rect 41823 -10782 41867 -10738
rect 41923 -10782 41967 -10738
rect 42023 -10782 42067 -10738
rect 42123 -10782 42167 -10738
rect 42223 -10782 42267 -10738
rect 42323 -10782 42367 -10738
rect 42423 -10782 42467 -10738
rect 42523 -10782 42567 -10738
rect 42623 -10782 42667 -10738
rect 42723 -10782 42767 -10738
rect 43223 -10782 43267 -10738
rect 43323 -10782 43367 -10738
rect 43423 -10782 43467 -10738
rect 43523 -10782 43567 -10738
rect 43623 -10782 43667 -10738
rect 43723 -10782 43767 -10738
rect 43823 -10782 43867 -10738
rect 43923 -10782 43967 -10738
rect 44023 -10782 44067 -10738
rect 44123 -10782 44167 -10738
rect 44223 -10782 44267 -10738
rect 44323 -10782 44367 -10738
rect 44423 -10782 44467 -10738
rect 44523 -10782 44567 -10738
rect 44623 -10782 44667 -10738
rect 44723 -10782 44767 -10738
rect 37223 -10882 37267 -10838
rect 37323 -10882 37367 -10838
rect 37423 -10882 37467 -10838
rect 37523 -10882 37567 -10838
rect 37623 -10882 37667 -10838
rect 37723 -10882 37767 -10838
rect 37823 -10882 37867 -10838
rect 37923 -10882 37967 -10838
rect 38023 -10882 38067 -10838
rect 38123 -10882 38167 -10838
rect 38223 -10882 38267 -10838
rect 38323 -10882 38367 -10838
rect 38423 -10882 38467 -10838
rect 38523 -10882 38567 -10838
rect 38623 -10882 38667 -10838
rect 38723 -10882 38767 -10838
rect 39223 -10882 39267 -10838
rect 39323 -10882 39367 -10838
rect 39423 -10882 39467 -10838
rect 39523 -10882 39567 -10838
rect 39623 -10882 39667 -10838
rect 39723 -10882 39767 -10838
rect 39823 -10882 39867 -10838
rect 39923 -10882 39967 -10838
rect 40023 -10882 40067 -10838
rect 40123 -10882 40167 -10838
rect 40223 -10882 40267 -10838
rect 40323 -10882 40367 -10838
rect 40423 -10882 40467 -10838
rect 40523 -10882 40567 -10838
rect 40623 -10882 40667 -10838
rect 40723 -10882 40767 -10838
rect 41223 -10882 41267 -10838
rect 41323 -10882 41367 -10838
rect 41423 -10882 41467 -10838
rect 41523 -10882 41567 -10838
rect 41623 -10882 41667 -10838
rect 41723 -10882 41767 -10838
rect 41823 -10882 41867 -10838
rect 41923 -10882 41967 -10838
rect 42023 -10882 42067 -10838
rect 42123 -10882 42167 -10838
rect 42223 -10882 42267 -10838
rect 42323 -10882 42367 -10838
rect 42423 -10882 42467 -10838
rect 42523 -10882 42567 -10838
rect 42623 -10882 42667 -10838
rect 42723 -10882 42767 -10838
rect 43223 -10882 43267 -10838
rect 43323 -10882 43367 -10838
rect 43423 -10882 43467 -10838
rect 43523 -10882 43567 -10838
rect 43623 -10882 43667 -10838
rect 43723 -10882 43767 -10838
rect 43823 -10882 43867 -10838
rect 43923 -10882 43967 -10838
rect 44023 -10882 44067 -10838
rect 44123 -10882 44167 -10838
rect 44223 -10882 44267 -10838
rect 44323 -10882 44367 -10838
rect 44423 -10882 44467 -10838
rect 44523 -10882 44567 -10838
rect 44623 -10882 44667 -10838
rect 44723 -10882 44767 -10838
rect 37223 -10982 37267 -10938
rect 37323 -10982 37367 -10938
rect 37423 -10982 37467 -10938
rect 37523 -10982 37567 -10938
rect 37623 -10982 37667 -10938
rect 37723 -10982 37767 -10938
rect 37823 -10982 37867 -10938
rect 37923 -10982 37967 -10938
rect 38023 -10982 38067 -10938
rect 38123 -10982 38167 -10938
rect 38223 -10982 38267 -10938
rect 38323 -10982 38367 -10938
rect 38423 -10982 38467 -10938
rect 38523 -10982 38567 -10938
rect 38623 -10982 38667 -10938
rect 38723 -10982 38767 -10938
rect 39223 -10982 39267 -10938
rect 39323 -10982 39367 -10938
rect 39423 -10982 39467 -10938
rect 39523 -10982 39567 -10938
rect 39623 -10982 39667 -10938
rect 39723 -10982 39767 -10938
rect 39823 -10982 39867 -10938
rect 39923 -10982 39967 -10938
rect 40023 -10982 40067 -10938
rect 40123 -10982 40167 -10938
rect 40223 -10982 40267 -10938
rect 40323 -10982 40367 -10938
rect 40423 -10982 40467 -10938
rect 40523 -10982 40567 -10938
rect 40623 -10982 40667 -10938
rect 40723 -10982 40767 -10938
rect 41223 -10982 41267 -10938
rect 41323 -10982 41367 -10938
rect 41423 -10982 41467 -10938
rect 41523 -10982 41567 -10938
rect 41623 -10982 41667 -10938
rect 41723 -10982 41767 -10938
rect 41823 -10982 41867 -10938
rect 41923 -10982 41967 -10938
rect 42023 -10982 42067 -10938
rect 42123 -10982 42167 -10938
rect 42223 -10982 42267 -10938
rect 42323 -10982 42367 -10938
rect 42423 -10982 42467 -10938
rect 42523 -10982 42567 -10938
rect 42623 -10982 42667 -10938
rect 42723 -10982 42767 -10938
rect 43223 -10982 43267 -10938
rect 43323 -10982 43367 -10938
rect 43423 -10982 43467 -10938
rect 43523 -10982 43567 -10938
rect 43623 -10982 43667 -10938
rect 43723 -10982 43767 -10938
rect 43823 -10982 43867 -10938
rect 43923 -10982 43967 -10938
rect 44023 -10982 44067 -10938
rect 44123 -10982 44167 -10938
rect 44223 -10982 44267 -10938
rect 44323 -10982 44367 -10938
rect 44423 -10982 44467 -10938
rect 44523 -10982 44567 -10938
rect 44623 -10982 44667 -10938
rect 44723 -10982 44767 -10938
rect 37223 -11082 37267 -11038
rect 37323 -11082 37367 -11038
rect 37423 -11082 37467 -11038
rect 37523 -11082 37567 -11038
rect 37623 -11082 37667 -11038
rect 37723 -11082 37767 -11038
rect 37823 -11082 37867 -11038
rect 37923 -11082 37967 -11038
rect 38023 -11082 38067 -11038
rect 38123 -11082 38167 -11038
rect 38223 -11082 38267 -11038
rect 38323 -11082 38367 -11038
rect 38423 -11082 38467 -11038
rect 38523 -11082 38567 -11038
rect 38623 -11082 38667 -11038
rect 38723 -11082 38767 -11038
rect 39223 -11082 39267 -11038
rect 39323 -11082 39367 -11038
rect 39423 -11082 39467 -11038
rect 39523 -11082 39567 -11038
rect 39623 -11082 39667 -11038
rect 39723 -11082 39767 -11038
rect 39823 -11082 39867 -11038
rect 39923 -11082 39967 -11038
rect 40023 -11082 40067 -11038
rect 40123 -11082 40167 -11038
rect 40223 -11082 40267 -11038
rect 40323 -11082 40367 -11038
rect 40423 -11082 40467 -11038
rect 40523 -11082 40567 -11038
rect 40623 -11082 40667 -11038
rect 40723 -11082 40767 -11038
rect 41223 -11082 41267 -11038
rect 41323 -11082 41367 -11038
rect 41423 -11082 41467 -11038
rect 41523 -11082 41567 -11038
rect 41623 -11082 41667 -11038
rect 41723 -11082 41767 -11038
rect 41823 -11082 41867 -11038
rect 41923 -11082 41967 -11038
rect 42023 -11082 42067 -11038
rect 42123 -11082 42167 -11038
rect 42223 -11082 42267 -11038
rect 42323 -11082 42367 -11038
rect 42423 -11082 42467 -11038
rect 42523 -11082 42567 -11038
rect 42623 -11082 42667 -11038
rect 42723 -11082 42767 -11038
rect 43223 -11082 43267 -11038
rect 43323 -11082 43367 -11038
rect 43423 -11082 43467 -11038
rect 43523 -11082 43567 -11038
rect 43623 -11082 43667 -11038
rect 43723 -11082 43767 -11038
rect 43823 -11082 43867 -11038
rect 43923 -11082 43967 -11038
rect 44023 -11082 44067 -11038
rect 44123 -11082 44167 -11038
rect 44223 -11082 44267 -11038
rect 44323 -11082 44367 -11038
rect 44423 -11082 44467 -11038
rect 44523 -11082 44567 -11038
rect 44623 -11082 44667 -11038
rect 44723 -11082 44767 -11038
rect 37223 -11182 37267 -11138
rect 37323 -11182 37367 -11138
rect 37423 -11182 37467 -11138
rect 37523 -11182 37567 -11138
rect 37623 -11182 37667 -11138
rect 37723 -11182 37767 -11138
rect 37823 -11182 37867 -11138
rect 37923 -11182 37967 -11138
rect 38023 -11182 38067 -11138
rect 38123 -11182 38167 -11138
rect 38223 -11182 38267 -11138
rect 38323 -11182 38367 -11138
rect 38423 -11182 38467 -11138
rect 38523 -11182 38567 -11138
rect 38623 -11182 38667 -11138
rect 38723 -11182 38767 -11138
rect 39223 -11182 39267 -11138
rect 39323 -11182 39367 -11138
rect 39423 -11182 39467 -11138
rect 39523 -11182 39567 -11138
rect 39623 -11182 39667 -11138
rect 39723 -11182 39767 -11138
rect 39823 -11182 39867 -11138
rect 39923 -11182 39967 -11138
rect 40023 -11182 40067 -11138
rect 40123 -11182 40167 -11138
rect 40223 -11182 40267 -11138
rect 40323 -11182 40367 -11138
rect 40423 -11182 40467 -11138
rect 40523 -11182 40567 -11138
rect 40623 -11182 40667 -11138
rect 40723 -11182 40767 -11138
rect 41223 -11182 41267 -11138
rect 41323 -11182 41367 -11138
rect 41423 -11182 41467 -11138
rect 41523 -11182 41567 -11138
rect 41623 -11182 41667 -11138
rect 41723 -11182 41767 -11138
rect 41823 -11182 41867 -11138
rect 41923 -11182 41967 -11138
rect 42023 -11182 42067 -11138
rect 42123 -11182 42167 -11138
rect 42223 -11182 42267 -11138
rect 42323 -11182 42367 -11138
rect 42423 -11182 42467 -11138
rect 42523 -11182 42567 -11138
rect 42623 -11182 42667 -11138
rect 42723 -11182 42767 -11138
rect 43223 -11182 43267 -11138
rect 43323 -11182 43367 -11138
rect 43423 -11182 43467 -11138
rect 43523 -11182 43567 -11138
rect 43623 -11182 43667 -11138
rect 43723 -11182 43767 -11138
rect 43823 -11182 43867 -11138
rect 43923 -11182 43967 -11138
rect 44023 -11182 44067 -11138
rect 44123 -11182 44167 -11138
rect 44223 -11182 44267 -11138
rect 44323 -11182 44367 -11138
rect 44423 -11182 44467 -11138
rect 44523 -11182 44567 -11138
rect 44623 -11182 44667 -11138
rect 44723 -11182 44767 -11138
rect 144904 -17489 144948 -17445
rect 145004 -17489 145048 -17445
rect 145104 -17489 145148 -17445
rect 145204 -17489 145248 -17445
rect 145304 -17489 145348 -17445
rect 145404 -17489 145448 -17445
rect 145504 -17489 145548 -17445
rect 145604 -17489 145648 -17445
rect 145704 -17489 145748 -17445
rect 145804 -17489 145848 -17445
rect 145904 -17489 145948 -17445
rect 146004 -17489 146048 -17445
rect 146104 -17489 146148 -17445
rect 146204 -17489 146248 -17445
rect 146304 -17489 146348 -17445
rect 146404 -17489 146448 -17445
rect 146904 -17489 146948 -17445
rect 147004 -17489 147048 -17445
rect 147104 -17489 147148 -17445
rect 147204 -17489 147248 -17445
rect 147304 -17489 147348 -17445
rect 147404 -17489 147448 -17445
rect 147504 -17489 147548 -17445
rect 147604 -17489 147648 -17445
rect 147704 -17489 147748 -17445
rect 147804 -17489 147848 -17445
rect 147904 -17489 147948 -17445
rect 148004 -17489 148048 -17445
rect 148104 -17489 148148 -17445
rect 148204 -17489 148248 -17445
rect 148304 -17489 148348 -17445
rect 148404 -17489 148448 -17445
rect 148904 -17489 148948 -17445
rect 149004 -17489 149048 -17445
rect 149104 -17489 149148 -17445
rect 149204 -17489 149248 -17445
rect 149304 -17489 149348 -17445
rect 149404 -17489 149448 -17445
rect 149504 -17489 149548 -17445
rect 149604 -17489 149648 -17445
rect 149704 -17489 149748 -17445
rect 149804 -17489 149848 -17445
rect 149904 -17489 149948 -17445
rect 150004 -17489 150048 -17445
rect 150104 -17489 150148 -17445
rect 150204 -17489 150248 -17445
rect 150304 -17489 150348 -17445
rect 150404 -17489 150448 -17445
rect 150904 -17489 150948 -17445
rect 151004 -17489 151048 -17445
rect 151104 -17489 151148 -17445
rect 151204 -17489 151248 -17445
rect 151304 -17489 151348 -17445
rect 151404 -17489 151448 -17445
rect 151504 -17489 151548 -17445
rect 151604 -17489 151648 -17445
rect 151704 -17489 151748 -17445
rect 151804 -17489 151848 -17445
rect 151904 -17489 151948 -17445
rect 152004 -17489 152048 -17445
rect 152104 -17489 152148 -17445
rect 152204 -17489 152248 -17445
rect 152304 -17489 152348 -17445
rect 152404 -17489 152448 -17445
rect 144904 -17589 144948 -17545
rect 145004 -17589 145048 -17545
rect 145104 -17589 145148 -17545
rect 145204 -17589 145248 -17545
rect 145304 -17589 145348 -17545
rect 145404 -17589 145448 -17545
rect 145504 -17589 145548 -17545
rect 145604 -17589 145648 -17545
rect 145704 -17589 145748 -17545
rect 145804 -17589 145848 -17545
rect 145904 -17589 145948 -17545
rect 146004 -17589 146048 -17545
rect 146104 -17589 146148 -17545
rect 146204 -17589 146248 -17545
rect 146304 -17589 146348 -17545
rect 146404 -17589 146448 -17545
rect 146904 -17589 146948 -17545
rect 147004 -17589 147048 -17545
rect 147104 -17589 147148 -17545
rect 147204 -17589 147248 -17545
rect 147304 -17589 147348 -17545
rect 147404 -17589 147448 -17545
rect 147504 -17589 147548 -17545
rect 147604 -17589 147648 -17545
rect 147704 -17589 147748 -17545
rect 147804 -17589 147848 -17545
rect 147904 -17589 147948 -17545
rect 148004 -17589 148048 -17545
rect 148104 -17589 148148 -17545
rect 148204 -17589 148248 -17545
rect 148304 -17589 148348 -17545
rect 148404 -17589 148448 -17545
rect 148904 -17589 148948 -17545
rect 149004 -17589 149048 -17545
rect 149104 -17589 149148 -17545
rect 149204 -17589 149248 -17545
rect 149304 -17589 149348 -17545
rect 149404 -17589 149448 -17545
rect 149504 -17589 149548 -17545
rect 149604 -17589 149648 -17545
rect 149704 -17589 149748 -17545
rect 149804 -17589 149848 -17545
rect 149904 -17589 149948 -17545
rect 150004 -17589 150048 -17545
rect 150104 -17589 150148 -17545
rect 150204 -17589 150248 -17545
rect 150304 -17589 150348 -17545
rect 150404 -17589 150448 -17545
rect 150904 -17589 150948 -17545
rect 151004 -17589 151048 -17545
rect 151104 -17589 151148 -17545
rect 151204 -17589 151248 -17545
rect 151304 -17589 151348 -17545
rect 151404 -17589 151448 -17545
rect 151504 -17589 151548 -17545
rect 151604 -17589 151648 -17545
rect 151704 -17589 151748 -17545
rect 151804 -17589 151848 -17545
rect 151904 -17589 151948 -17545
rect 152004 -17589 152048 -17545
rect 152104 -17589 152148 -17545
rect 152204 -17589 152248 -17545
rect 152304 -17589 152348 -17545
rect 152404 -17589 152448 -17545
rect 144904 -17689 144948 -17645
rect 145004 -17689 145048 -17645
rect 145104 -17689 145148 -17645
rect 145204 -17689 145248 -17645
rect 145304 -17689 145348 -17645
rect 145404 -17689 145448 -17645
rect 145504 -17689 145548 -17645
rect 145604 -17689 145648 -17645
rect 145704 -17689 145748 -17645
rect 145804 -17689 145848 -17645
rect 145904 -17689 145948 -17645
rect 146004 -17689 146048 -17645
rect 146104 -17689 146148 -17645
rect 146204 -17689 146248 -17645
rect 146304 -17689 146348 -17645
rect 146404 -17689 146448 -17645
rect 146904 -17689 146948 -17645
rect 147004 -17689 147048 -17645
rect 147104 -17689 147148 -17645
rect 147204 -17689 147248 -17645
rect 147304 -17689 147348 -17645
rect 147404 -17689 147448 -17645
rect 147504 -17689 147548 -17645
rect 147604 -17689 147648 -17645
rect 147704 -17689 147748 -17645
rect 147804 -17689 147848 -17645
rect 147904 -17689 147948 -17645
rect 148004 -17689 148048 -17645
rect 148104 -17689 148148 -17645
rect 148204 -17689 148248 -17645
rect 148304 -17689 148348 -17645
rect 148404 -17689 148448 -17645
rect 148904 -17689 148948 -17645
rect 149004 -17689 149048 -17645
rect 149104 -17689 149148 -17645
rect 149204 -17689 149248 -17645
rect 149304 -17689 149348 -17645
rect 149404 -17689 149448 -17645
rect 149504 -17689 149548 -17645
rect 149604 -17689 149648 -17645
rect 149704 -17689 149748 -17645
rect 149804 -17689 149848 -17645
rect 149904 -17689 149948 -17645
rect 150004 -17689 150048 -17645
rect 150104 -17689 150148 -17645
rect 150204 -17689 150248 -17645
rect 150304 -17689 150348 -17645
rect 150404 -17689 150448 -17645
rect 150904 -17689 150948 -17645
rect 151004 -17689 151048 -17645
rect 151104 -17689 151148 -17645
rect 151204 -17689 151248 -17645
rect 151304 -17689 151348 -17645
rect 151404 -17689 151448 -17645
rect 151504 -17689 151548 -17645
rect 151604 -17689 151648 -17645
rect 151704 -17689 151748 -17645
rect 151804 -17689 151848 -17645
rect 151904 -17689 151948 -17645
rect 152004 -17689 152048 -17645
rect 152104 -17689 152148 -17645
rect 152204 -17689 152248 -17645
rect 152304 -17689 152348 -17645
rect 152404 -17689 152448 -17645
rect 144904 -17789 144948 -17745
rect 145004 -17789 145048 -17745
rect 145104 -17789 145148 -17745
rect 145204 -17789 145248 -17745
rect 145304 -17789 145348 -17745
rect 145404 -17789 145448 -17745
rect 145504 -17789 145548 -17745
rect 145604 -17789 145648 -17745
rect 145704 -17789 145748 -17745
rect 145804 -17789 145848 -17745
rect 145904 -17789 145948 -17745
rect 146004 -17789 146048 -17745
rect 146104 -17789 146148 -17745
rect 146204 -17789 146248 -17745
rect 146304 -17789 146348 -17745
rect 146404 -17789 146448 -17745
rect 146904 -17789 146948 -17745
rect 147004 -17789 147048 -17745
rect 147104 -17789 147148 -17745
rect 147204 -17789 147248 -17745
rect 147304 -17789 147348 -17745
rect 147404 -17789 147448 -17745
rect 147504 -17789 147548 -17745
rect 147604 -17789 147648 -17745
rect 147704 -17789 147748 -17745
rect 147804 -17789 147848 -17745
rect 147904 -17789 147948 -17745
rect 148004 -17789 148048 -17745
rect 148104 -17789 148148 -17745
rect 148204 -17789 148248 -17745
rect 148304 -17789 148348 -17745
rect 148404 -17789 148448 -17745
rect 148904 -17789 148948 -17745
rect 149004 -17789 149048 -17745
rect 149104 -17789 149148 -17745
rect 149204 -17789 149248 -17745
rect 149304 -17789 149348 -17745
rect 149404 -17789 149448 -17745
rect 149504 -17789 149548 -17745
rect 149604 -17789 149648 -17745
rect 149704 -17789 149748 -17745
rect 149804 -17789 149848 -17745
rect 149904 -17789 149948 -17745
rect 150004 -17789 150048 -17745
rect 150104 -17789 150148 -17745
rect 150204 -17789 150248 -17745
rect 150304 -17789 150348 -17745
rect 150404 -17789 150448 -17745
rect 150904 -17789 150948 -17745
rect 151004 -17789 151048 -17745
rect 151104 -17789 151148 -17745
rect 151204 -17789 151248 -17745
rect 151304 -17789 151348 -17745
rect 151404 -17789 151448 -17745
rect 151504 -17789 151548 -17745
rect 151604 -17789 151648 -17745
rect 151704 -17789 151748 -17745
rect 151804 -17789 151848 -17745
rect 151904 -17789 151948 -17745
rect 152004 -17789 152048 -17745
rect 152104 -17789 152148 -17745
rect 152204 -17789 152248 -17745
rect 152304 -17789 152348 -17745
rect 152404 -17789 152448 -17745
rect 173611 -17830 174124 -17214
rect 144904 -17889 144948 -17845
rect 145004 -17889 145048 -17845
rect 145104 -17889 145148 -17845
rect 145204 -17889 145248 -17845
rect 145304 -17889 145348 -17845
rect 145404 -17889 145448 -17845
rect 145504 -17889 145548 -17845
rect 145604 -17889 145648 -17845
rect 145704 -17889 145748 -17845
rect 145804 -17889 145848 -17845
rect 145904 -17889 145948 -17845
rect 146004 -17889 146048 -17845
rect 146104 -17889 146148 -17845
rect 146204 -17889 146248 -17845
rect 146304 -17889 146348 -17845
rect 146404 -17889 146448 -17845
rect 146904 -17889 146948 -17845
rect 147004 -17889 147048 -17845
rect 147104 -17889 147148 -17845
rect 147204 -17889 147248 -17845
rect 147304 -17889 147348 -17845
rect 147404 -17889 147448 -17845
rect 147504 -17889 147548 -17845
rect 147604 -17889 147648 -17845
rect 147704 -17889 147748 -17845
rect 147804 -17889 147848 -17845
rect 147904 -17889 147948 -17845
rect 148004 -17889 148048 -17845
rect 148104 -17889 148148 -17845
rect 148204 -17889 148248 -17845
rect 148304 -17889 148348 -17845
rect 148404 -17889 148448 -17845
rect 148904 -17889 148948 -17845
rect 149004 -17889 149048 -17845
rect 149104 -17889 149148 -17845
rect 149204 -17889 149248 -17845
rect 149304 -17889 149348 -17845
rect 149404 -17889 149448 -17845
rect 149504 -17889 149548 -17845
rect 149604 -17889 149648 -17845
rect 149704 -17889 149748 -17845
rect 149804 -17889 149848 -17845
rect 149904 -17889 149948 -17845
rect 150004 -17889 150048 -17845
rect 150104 -17889 150148 -17845
rect 150204 -17889 150248 -17845
rect 150304 -17889 150348 -17845
rect 150404 -17889 150448 -17845
rect 150904 -17889 150948 -17845
rect 151004 -17889 151048 -17845
rect 151104 -17889 151148 -17845
rect 151204 -17889 151248 -17845
rect 151304 -17889 151348 -17845
rect 151404 -17889 151448 -17845
rect 151504 -17889 151548 -17845
rect 151604 -17889 151648 -17845
rect 151704 -17889 151748 -17845
rect 151804 -17889 151848 -17845
rect 151904 -17889 151948 -17845
rect 152004 -17889 152048 -17845
rect 152104 -17889 152148 -17845
rect 152204 -17889 152248 -17845
rect 152304 -17889 152348 -17845
rect 152404 -17889 152448 -17845
rect 144904 -17989 144948 -17945
rect 145004 -17989 145048 -17945
rect 145104 -17989 145148 -17945
rect 145204 -17989 145248 -17945
rect 145304 -17989 145348 -17945
rect 145404 -17989 145448 -17945
rect 145504 -17989 145548 -17945
rect 145604 -17989 145648 -17945
rect 145704 -17989 145748 -17945
rect 145804 -17989 145848 -17945
rect 145904 -17989 145948 -17945
rect 146004 -17989 146048 -17945
rect 146104 -17989 146148 -17945
rect 146204 -17989 146248 -17945
rect 146304 -17989 146348 -17945
rect 146404 -17989 146448 -17945
rect 146904 -17989 146948 -17945
rect 147004 -17989 147048 -17945
rect 147104 -17989 147148 -17945
rect 147204 -17989 147248 -17945
rect 147304 -17989 147348 -17945
rect 147404 -17989 147448 -17945
rect 147504 -17989 147548 -17945
rect 147604 -17989 147648 -17945
rect 147704 -17989 147748 -17945
rect 147804 -17989 147848 -17945
rect 147904 -17989 147948 -17945
rect 148004 -17989 148048 -17945
rect 148104 -17989 148148 -17945
rect 148204 -17989 148248 -17945
rect 148304 -17989 148348 -17945
rect 148404 -17989 148448 -17945
rect 148904 -17989 148948 -17945
rect 149004 -17989 149048 -17945
rect 149104 -17989 149148 -17945
rect 149204 -17989 149248 -17945
rect 149304 -17989 149348 -17945
rect 149404 -17989 149448 -17945
rect 149504 -17989 149548 -17945
rect 149604 -17989 149648 -17945
rect 149704 -17989 149748 -17945
rect 149804 -17989 149848 -17945
rect 149904 -17989 149948 -17945
rect 150004 -17989 150048 -17945
rect 150104 -17989 150148 -17945
rect 150204 -17989 150248 -17945
rect 150304 -17989 150348 -17945
rect 150404 -17989 150448 -17945
rect 150904 -17989 150948 -17945
rect 151004 -17989 151048 -17945
rect 151104 -17989 151148 -17945
rect 151204 -17989 151248 -17945
rect 151304 -17989 151348 -17945
rect 151404 -17989 151448 -17945
rect 151504 -17989 151548 -17945
rect 151604 -17989 151648 -17945
rect 151704 -17989 151748 -17945
rect 151804 -17989 151848 -17945
rect 151904 -17989 151948 -17945
rect 152004 -17989 152048 -17945
rect 152104 -17989 152148 -17945
rect 152204 -17989 152248 -17945
rect 152304 -17989 152348 -17945
rect 152404 -17989 152448 -17945
rect 144904 -18089 144948 -18045
rect 145004 -18089 145048 -18045
rect 145104 -18089 145148 -18045
rect 145204 -18089 145248 -18045
rect 145304 -18089 145348 -18045
rect 145404 -18089 145448 -18045
rect 145504 -18089 145548 -18045
rect 145604 -18089 145648 -18045
rect 145704 -18089 145748 -18045
rect 145804 -18089 145848 -18045
rect 145904 -18089 145948 -18045
rect 146004 -18089 146048 -18045
rect 146104 -18089 146148 -18045
rect 146204 -18089 146248 -18045
rect 146304 -18089 146348 -18045
rect 146404 -18089 146448 -18045
rect 146904 -18089 146948 -18045
rect 147004 -18089 147048 -18045
rect 147104 -18089 147148 -18045
rect 147204 -18089 147248 -18045
rect 147304 -18089 147348 -18045
rect 147404 -18089 147448 -18045
rect 147504 -18089 147548 -18045
rect 147604 -18089 147648 -18045
rect 147704 -18089 147748 -18045
rect 147804 -18089 147848 -18045
rect 147904 -18089 147948 -18045
rect 148004 -18089 148048 -18045
rect 148104 -18089 148148 -18045
rect 148204 -18089 148248 -18045
rect 148304 -18089 148348 -18045
rect 148404 -18089 148448 -18045
rect 148904 -18089 148948 -18045
rect 149004 -18089 149048 -18045
rect 149104 -18089 149148 -18045
rect 149204 -18089 149248 -18045
rect 149304 -18089 149348 -18045
rect 149404 -18089 149448 -18045
rect 149504 -18089 149548 -18045
rect 149604 -18089 149648 -18045
rect 149704 -18089 149748 -18045
rect 149804 -18089 149848 -18045
rect 149904 -18089 149948 -18045
rect 150004 -18089 150048 -18045
rect 150104 -18089 150148 -18045
rect 150204 -18089 150248 -18045
rect 150304 -18089 150348 -18045
rect 150404 -18089 150448 -18045
rect 150904 -18089 150948 -18045
rect 151004 -18089 151048 -18045
rect 151104 -18089 151148 -18045
rect 151204 -18089 151248 -18045
rect 151304 -18089 151348 -18045
rect 151404 -18089 151448 -18045
rect 151504 -18089 151548 -18045
rect 151604 -18089 151648 -18045
rect 151704 -18089 151748 -18045
rect 151804 -18089 151848 -18045
rect 151904 -18089 151948 -18045
rect 152004 -18089 152048 -18045
rect 152104 -18089 152148 -18045
rect 152204 -18089 152248 -18045
rect 152304 -18089 152348 -18045
rect 152404 -18089 152448 -18045
rect 144904 -18189 144948 -18145
rect 145004 -18189 145048 -18145
rect 145104 -18189 145148 -18145
rect 145204 -18189 145248 -18145
rect 145304 -18189 145348 -18145
rect 145404 -18189 145448 -18145
rect 145504 -18189 145548 -18145
rect 145604 -18189 145648 -18145
rect 145704 -18189 145748 -18145
rect 145804 -18189 145848 -18145
rect 145904 -18189 145948 -18145
rect 146004 -18189 146048 -18145
rect 146104 -18189 146148 -18145
rect 146204 -18189 146248 -18145
rect 146304 -18189 146348 -18145
rect 146404 -18189 146448 -18145
rect 146904 -18189 146948 -18145
rect 147004 -18189 147048 -18145
rect 147104 -18189 147148 -18145
rect 147204 -18189 147248 -18145
rect 147304 -18189 147348 -18145
rect 147404 -18189 147448 -18145
rect 147504 -18189 147548 -18145
rect 147604 -18189 147648 -18145
rect 147704 -18189 147748 -18145
rect 147804 -18189 147848 -18145
rect 147904 -18189 147948 -18145
rect 148004 -18189 148048 -18145
rect 148104 -18189 148148 -18145
rect 148204 -18189 148248 -18145
rect 148304 -18189 148348 -18145
rect 148404 -18189 148448 -18145
rect 148904 -18189 148948 -18145
rect 149004 -18189 149048 -18145
rect 149104 -18189 149148 -18145
rect 149204 -18189 149248 -18145
rect 149304 -18189 149348 -18145
rect 149404 -18189 149448 -18145
rect 149504 -18189 149548 -18145
rect 149604 -18189 149648 -18145
rect 149704 -18189 149748 -18145
rect 149804 -18189 149848 -18145
rect 149904 -18189 149948 -18145
rect 150004 -18189 150048 -18145
rect 150104 -18189 150148 -18145
rect 150204 -18189 150248 -18145
rect 150304 -18189 150348 -18145
rect 150404 -18189 150448 -18145
rect 150904 -18189 150948 -18145
rect 151004 -18189 151048 -18145
rect 151104 -18189 151148 -18145
rect 151204 -18189 151248 -18145
rect 151304 -18189 151348 -18145
rect 151404 -18189 151448 -18145
rect 151504 -18189 151548 -18145
rect 151604 -18189 151648 -18145
rect 151704 -18189 151748 -18145
rect 151804 -18189 151848 -18145
rect 151904 -18189 151948 -18145
rect 152004 -18189 152048 -18145
rect 152104 -18189 152148 -18145
rect 152204 -18189 152248 -18145
rect 152304 -18189 152348 -18145
rect 152404 -18189 152448 -18145
rect 144904 -18289 144948 -18245
rect 145004 -18289 145048 -18245
rect 145104 -18289 145148 -18245
rect 145204 -18289 145248 -18245
rect 145304 -18289 145348 -18245
rect 145404 -18289 145448 -18245
rect 145504 -18289 145548 -18245
rect 145604 -18289 145648 -18245
rect 145704 -18289 145748 -18245
rect 145804 -18289 145848 -18245
rect 145904 -18289 145948 -18245
rect 146004 -18289 146048 -18245
rect 146104 -18289 146148 -18245
rect 146204 -18289 146248 -18245
rect 146304 -18289 146348 -18245
rect 146404 -18289 146448 -18245
rect 146904 -18289 146948 -18245
rect 147004 -18289 147048 -18245
rect 147104 -18289 147148 -18245
rect 147204 -18289 147248 -18245
rect 147304 -18289 147348 -18245
rect 147404 -18289 147448 -18245
rect 147504 -18289 147548 -18245
rect 147604 -18289 147648 -18245
rect 147704 -18289 147748 -18245
rect 147804 -18289 147848 -18245
rect 147904 -18289 147948 -18245
rect 148004 -18289 148048 -18245
rect 148104 -18289 148148 -18245
rect 148204 -18289 148248 -18245
rect 148304 -18289 148348 -18245
rect 148404 -18289 148448 -18245
rect 148904 -18289 148948 -18245
rect 149004 -18289 149048 -18245
rect 149104 -18289 149148 -18245
rect 149204 -18289 149248 -18245
rect 149304 -18289 149348 -18245
rect 149404 -18289 149448 -18245
rect 149504 -18289 149548 -18245
rect 149604 -18289 149648 -18245
rect 149704 -18289 149748 -18245
rect 149804 -18289 149848 -18245
rect 149904 -18289 149948 -18245
rect 150004 -18289 150048 -18245
rect 150104 -18289 150148 -18245
rect 150204 -18289 150248 -18245
rect 150304 -18289 150348 -18245
rect 150404 -18289 150448 -18245
rect 150904 -18289 150948 -18245
rect 151004 -18289 151048 -18245
rect 151104 -18289 151148 -18245
rect 151204 -18289 151248 -18245
rect 151304 -18289 151348 -18245
rect 151404 -18289 151448 -18245
rect 151504 -18289 151548 -18245
rect 151604 -18289 151648 -18245
rect 151704 -18289 151748 -18245
rect 151804 -18289 151848 -18245
rect 151904 -18289 151948 -18245
rect 152004 -18289 152048 -18245
rect 152104 -18289 152148 -18245
rect 152204 -18289 152248 -18245
rect 152304 -18289 152348 -18245
rect 152404 -18289 152448 -18245
rect 144904 -18389 144948 -18345
rect 145004 -18389 145048 -18345
rect 145104 -18389 145148 -18345
rect 145204 -18389 145248 -18345
rect 145304 -18389 145348 -18345
rect 145404 -18389 145448 -18345
rect 145504 -18389 145548 -18345
rect 145604 -18389 145648 -18345
rect 145704 -18389 145748 -18345
rect 145804 -18389 145848 -18345
rect 145904 -18389 145948 -18345
rect 146004 -18389 146048 -18345
rect 146104 -18389 146148 -18345
rect 146204 -18389 146248 -18345
rect 146304 -18389 146348 -18345
rect 146404 -18389 146448 -18345
rect 146904 -18389 146948 -18345
rect 147004 -18389 147048 -18345
rect 147104 -18389 147148 -18345
rect 147204 -18389 147248 -18345
rect 147304 -18389 147348 -18345
rect 147404 -18389 147448 -18345
rect 147504 -18389 147548 -18345
rect 147604 -18389 147648 -18345
rect 147704 -18389 147748 -18345
rect 147804 -18389 147848 -18345
rect 147904 -18389 147948 -18345
rect 148004 -18389 148048 -18345
rect 148104 -18389 148148 -18345
rect 148204 -18389 148248 -18345
rect 148304 -18389 148348 -18345
rect 148404 -18389 148448 -18345
rect 148904 -18389 148948 -18345
rect 149004 -18389 149048 -18345
rect 149104 -18389 149148 -18345
rect 149204 -18389 149248 -18345
rect 149304 -18389 149348 -18345
rect 149404 -18389 149448 -18345
rect 149504 -18389 149548 -18345
rect 149604 -18389 149648 -18345
rect 149704 -18389 149748 -18345
rect 149804 -18389 149848 -18345
rect 149904 -18389 149948 -18345
rect 150004 -18389 150048 -18345
rect 150104 -18389 150148 -18345
rect 150204 -18389 150248 -18345
rect 150304 -18389 150348 -18345
rect 150404 -18389 150448 -18345
rect 150904 -18389 150948 -18345
rect 151004 -18389 151048 -18345
rect 151104 -18389 151148 -18345
rect 151204 -18389 151248 -18345
rect 151304 -18389 151348 -18345
rect 151404 -18389 151448 -18345
rect 151504 -18389 151548 -18345
rect 151604 -18389 151648 -18345
rect 151704 -18389 151748 -18345
rect 151804 -18389 151848 -18345
rect 151904 -18389 151948 -18345
rect 152004 -18389 152048 -18345
rect 152104 -18389 152148 -18345
rect 152204 -18389 152248 -18345
rect 152304 -18389 152348 -18345
rect 152404 -18389 152448 -18345
rect 144904 -18489 144948 -18445
rect 145004 -18489 145048 -18445
rect 145104 -18489 145148 -18445
rect 145204 -18489 145248 -18445
rect 145304 -18489 145348 -18445
rect 145404 -18489 145448 -18445
rect 145504 -18489 145548 -18445
rect 145604 -18489 145648 -18445
rect 145704 -18489 145748 -18445
rect 145804 -18489 145848 -18445
rect 145904 -18489 145948 -18445
rect 146004 -18489 146048 -18445
rect 146104 -18489 146148 -18445
rect 146204 -18489 146248 -18445
rect 146304 -18489 146348 -18445
rect 146404 -18489 146448 -18445
rect 146904 -18489 146948 -18445
rect 147004 -18489 147048 -18445
rect 147104 -18489 147148 -18445
rect 147204 -18489 147248 -18445
rect 147304 -18489 147348 -18445
rect 147404 -18489 147448 -18445
rect 147504 -18489 147548 -18445
rect 147604 -18489 147648 -18445
rect 147704 -18489 147748 -18445
rect 147804 -18489 147848 -18445
rect 147904 -18489 147948 -18445
rect 148004 -18489 148048 -18445
rect 148104 -18489 148148 -18445
rect 148204 -18489 148248 -18445
rect 148304 -18489 148348 -18445
rect 148404 -18489 148448 -18445
rect 148904 -18489 148948 -18445
rect 149004 -18489 149048 -18445
rect 149104 -18489 149148 -18445
rect 149204 -18489 149248 -18445
rect 149304 -18489 149348 -18445
rect 149404 -18489 149448 -18445
rect 149504 -18489 149548 -18445
rect 149604 -18489 149648 -18445
rect 149704 -18489 149748 -18445
rect 149804 -18489 149848 -18445
rect 149904 -18489 149948 -18445
rect 150004 -18489 150048 -18445
rect 150104 -18489 150148 -18445
rect 150204 -18489 150248 -18445
rect 150304 -18489 150348 -18445
rect 150404 -18489 150448 -18445
rect 150904 -18489 150948 -18445
rect 151004 -18489 151048 -18445
rect 151104 -18489 151148 -18445
rect 151204 -18489 151248 -18445
rect 151304 -18489 151348 -18445
rect 151404 -18489 151448 -18445
rect 151504 -18489 151548 -18445
rect 151604 -18489 151648 -18445
rect 151704 -18489 151748 -18445
rect 151804 -18489 151848 -18445
rect 151904 -18489 151948 -18445
rect 152004 -18489 152048 -18445
rect 152104 -18489 152148 -18445
rect 152204 -18489 152248 -18445
rect 152304 -18489 152348 -18445
rect 152404 -18489 152448 -18445
rect 144904 -18589 144948 -18545
rect 145004 -18589 145048 -18545
rect 145104 -18589 145148 -18545
rect 145204 -18589 145248 -18545
rect 145304 -18589 145348 -18545
rect 145404 -18589 145448 -18545
rect 145504 -18589 145548 -18545
rect 145604 -18589 145648 -18545
rect 145704 -18589 145748 -18545
rect 145804 -18589 145848 -18545
rect 145904 -18589 145948 -18545
rect 146004 -18589 146048 -18545
rect 146104 -18589 146148 -18545
rect 146204 -18589 146248 -18545
rect 146304 -18589 146348 -18545
rect 146404 -18589 146448 -18545
rect 146904 -18589 146948 -18545
rect 147004 -18589 147048 -18545
rect 147104 -18589 147148 -18545
rect 147204 -18589 147248 -18545
rect 147304 -18589 147348 -18545
rect 147404 -18589 147448 -18545
rect 147504 -18589 147548 -18545
rect 147604 -18589 147648 -18545
rect 147704 -18589 147748 -18545
rect 147804 -18589 147848 -18545
rect 147904 -18589 147948 -18545
rect 148004 -18589 148048 -18545
rect 148104 -18589 148148 -18545
rect 148204 -18589 148248 -18545
rect 148304 -18589 148348 -18545
rect 148404 -18589 148448 -18545
rect 148904 -18589 148948 -18545
rect 149004 -18589 149048 -18545
rect 149104 -18589 149148 -18545
rect 149204 -18589 149248 -18545
rect 149304 -18589 149348 -18545
rect 149404 -18589 149448 -18545
rect 149504 -18589 149548 -18545
rect 149604 -18589 149648 -18545
rect 149704 -18589 149748 -18545
rect 149804 -18589 149848 -18545
rect 149904 -18589 149948 -18545
rect 150004 -18589 150048 -18545
rect 150104 -18589 150148 -18545
rect 150204 -18589 150248 -18545
rect 150304 -18589 150348 -18545
rect 150404 -18589 150448 -18545
rect 150904 -18589 150948 -18545
rect 151004 -18589 151048 -18545
rect 151104 -18589 151148 -18545
rect 151204 -18589 151248 -18545
rect 151304 -18589 151348 -18545
rect 151404 -18589 151448 -18545
rect 151504 -18589 151548 -18545
rect 151604 -18589 151648 -18545
rect 151704 -18589 151748 -18545
rect 151804 -18589 151848 -18545
rect 151904 -18589 151948 -18545
rect 152004 -18589 152048 -18545
rect 152104 -18589 152148 -18545
rect 152204 -18589 152248 -18545
rect 152304 -18589 152348 -18545
rect 152404 -18589 152448 -18545
rect 144904 -18689 144948 -18645
rect 145004 -18689 145048 -18645
rect 145104 -18689 145148 -18645
rect 145204 -18689 145248 -18645
rect 145304 -18689 145348 -18645
rect 145404 -18689 145448 -18645
rect 145504 -18689 145548 -18645
rect 145604 -18689 145648 -18645
rect 145704 -18689 145748 -18645
rect 145804 -18689 145848 -18645
rect 145904 -18689 145948 -18645
rect 146004 -18689 146048 -18645
rect 146104 -18689 146148 -18645
rect 146204 -18689 146248 -18645
rect 146304 -18689 146348 -18645
rect 146404 -18689 146448 -18645
rect 146904 -18689 146948 -18645
rect 147004 -18689 147048 -18645
rect 147104 -18689 147148 -18645
rect 147204 -18689 147248 -18645
rect 147304 -18689 147348 -18645
rect 147404 -18689 147448 -18645
rect 147504 -18689 147548 -18645
rect 147604 -18689 147648 -18645
rect 147704 -18689 147748 -18645
rect 147804 -18689 147848 -18645
rect 147904 -18689 147948 -18645
rect 148004 -18689 148048 -18645
rect 148104 -18689 148148 -18645
rect 148204 -18689 148248 -18645
rect 148304 -18689 148348 -18645
rect 148404 -18689 148448 -18645
rect 148904 -18689 148948 -18645
rect 149004 -18689 149048 -18645
rect 149104 -18689 149148 -18645
rect 149204 -18689 149248 -18645
rect 149304 -18689 149348 -18645
rect 149404 -18689 149448 -18645
rect 149504 -18689 149548 -18645
rect 149604 -18689 149648 -18645
rect 149704 -18689 149748 -18645
rect 149804 -18689 149848 -18645
rect 149904 -18689 149948 -18645
rect 150004 -18689 150048 -18645
rect 150104 -18689 150148 -18645
rect 150204 -18689 150248 -18645
rect 150304 -18689 150348 -18645
rect 150404 -18689 150448 -18645
rect 150904 -18689 150948 -18645
rect 151004 -18689 151048 -18645
rect 151104 -18689 151148 -18645
rect 151204 -18689 151248 -18645
rect 151304 -18689 151348 -18645
rect 151404 -18689 151448 -18645
rect 151504 -18689 151548 -18645
rect 151604 -18689 151648 -18645
rect 151704 -18689 151748 -18645
rect 151804 -18689 151848 -18645
rect 151904 -18689 151948 -18645
rect 152004 -18689 152048 -18645
rect 152104 -18689 152148 -18645
rect 152204 -18689 152248 -18645
rect 152304 -18689 152348 -18645
rect 152404 -18689 152448 -18645
rect 144904 -18789 144948 -18745
rect 145004 -18789 145048 -18745
rect 145104 -18789 145148 -18745
rect 145204 -18789 145248 -18745
rect 145304 -18789 145348 -18745
rect 145404 -18789 145448 -18745
rect 145504 -18789 145548 -18745
rect 145604 -18789 145648 -18745
rect 145704 -18789 145748 -18745
rect 145804 -18789 145848 -18745
rect 145904 -18789 145948 -18745
rect 146004 -18789 146048 -18745
rect 146104 -18789 146148 -18745
rect 146204 -18789 146248 -18745
rect 146304 -18789 146348 -18745
rect 146404 -18789 146448 -18745
rect 146904 -18789 146948 -18745
rect 147004 -18789 147048 -18745
rect 147104 -18789 147148 -18745
rect 147204 -18789 147248 -18745
rect 147304 -18789 147348 -18745
rect 147404 -18789 147448 -18745
rect 147504 -18789 147548 -18745
rect 147604 -18789 147648 -18745
rect 147704 -18789 147748 -18745
rect 147804 -18789 147848 -18745
rect 147904 -18789 147948 -18745
rect 148004 -18789 148048 -18745
rect 148104 -18789 148148 -18745
rect 148204 -18789 148248 -18745
rect 148304 -18789 148348 -18745
rect 148404 -18789 148448 -18745
rect 148904 -18789 148948 -18745
rect 149004 -18789 149048 -18745
rect 149104 -18789 149148 -18745
rect 149204 -18789 149248 -18745
rect 149304 -18789 149348 -18745
rect 149404 -18789 149448 -18745
rect 149504 -18789 149548 -18745
rect 149604 -18789 149648 -18745
rect 149704 -18789 149748 -18745
rect 149804 -18789 149848 -18745
rect 149904 -18789 149948 -18745
rect 150004 -18789 150048 -18745
rect 150104 -18789 150148 -18745
rect 150204 -18789 150248 -18745
rect 150304 -18789 150348 -18745
rect 150404 -18789 150448 -18745
rect 150904 -18789 150948 -18745
rect 151004 -18789 151048 -18745
rect 151104 -18789 151148 -18745
rect 151204 -18789 151248 -18745
rect 151304 -18789 151348 -18745
rect 151404 -18789 151448 -18745
rect 151504 -18789 151548 -18745
rect 151604 -18789 151648 -18745
rect 151704 -18789 151748 -18745
rect 151804 -18789 151848 -18745
rect 151904 -18789 151948 -18745
rect 152004 -18789 152048 -18745
rect 152104 -18789 152148 -18745
rect 152204 -18789 152248 -18745
rect 152304 -18789 152348 -18745
rect 152404 -18789 152448 -18745
rect 144904 -18889 144948 -18845
rect 145004 -18889 145048 -18845
rect 145104 -18889 145148 -18845
rect 145204 -18889 145248 -18845
rect 145304 -18889 145348 -18845
rect 145404 -18889 145448 -18845
rect 145504 -18889 145548 -18845
rect 145604 -18889 145648 -18845
rect 145704 -18889 145748 -18845
rect 145804 -18889 145848 -18845
rect 145904 -18889 145948 -18845
rect 146004 -18889 146048 -18845
rect 146104 -18889 146148 -18845
rect 146204 -18889 146248 -18845
rect 146304 -18889 146348 -18845
rect 146404 -18889 146448 -18845
rect 146904 -18889 146948 -18845
rect 147004 -18889 147048 -18845
rect 147104 -18889 147148 -18845
rect 147204 -18889 147248 -18845
rect 147304 -18889 147348 -18845
rect 147404 -18889 147448 -18845
rect 147504 -18889 147548 -18845
rect 147604 -18889 147648 -18845
rect 147704 -18889 147748 -18845
rect 147804 -18889 147848 -18845
rect 147904 -18889 147948 -18845
rect 148004 -18889 148048 -18845
rect 148104 -18889 148148 -18845
rect 148204 -18889 148248 -18845
rect 148304 -18889 148348 -18845
rect 148404 -18889 148448 -18845
rect 148904 -18889 148948 -18845
rect 149004 -18889 149048 -18845
rect 149104 -18889 149148 -18845
rect 149204 -18889 149248 -18845
rect 149304 -18889 149348 -18845
rect 149404 -18889 149448 -18845
rect 149504 -18889 149548 -18845
rect 149604 -18889 149648 -18845
rect 149704 -18889 149748 -18845
rect 149804 -18889 149848 -18845
rect 149904 -18889 149948 -18845
rect 150004 -18889 150048 -18845
rect 150104 -18889 150148 -18845
rect 150204 -18889 150248 -18845
rect 150304 -18889 150348 -18845
rect 150404 -18889 150448 -18845
rect 150904 -18889 150948 -18845
rect 151004 -18889 151048 -18845
rect 151104 -18889 151148 -18845
rect 151204 -18889 151248 -18845
rect 151304 -18889 151348 -18845
rect 151404 -18889 151448 -18845
rect 151504 -18889 151548 -18845
rect 151604 -18889 151648 -18845
rect 151704 -18889 151748 -18845
rect 151804 -18889 151848 -18845
rect 151904 -18889 151948 -18845
rect 152004 -18889 152048 -18845
rect 152104 -18889 152148 -18845
rect 152204 -18889 152248 -18845
rect 152304 -18889 152348 -18845
rect 152404 -18889 152448 -18845
rect 144904 -18989 144948 -18945
rect 145004 -18989 145048 -18945
rect 145104 -18989 145148 -18945
rect 145204 -18989 145248 -18945
rect 145304 -18989 145348 -18945
rect 145404 -18989 145448 -18945
rect 145504 -18989 145548 -18945
rect 145604 -18989 145648 -18945
rect 145704 -18989 145748 -18945
rect 145804 -18989 145848 -18945
rect 145904 -18989 145948 -18945
rect 146004 -18989 146048 -18945
rect 146104 -18989 146148 -18945
rect 146204 -18989 146248 -18945
rect 146304 -18989 146348 -18945
rect 146404 -18989 146448 -18945
rect 146904 -18989 146948 -18945
rect 147004 -18989 147048 -18945
rect 147104 -18989 147148 -18945
rect 147204 -18989 147248 -18945
rect 147304 -18989 147348 -18945
rect 147404 -18989 147448 -18945
rect 147504 -18989 147548 -18945
rect 147604 -18989 147648 -18945
rect 147704 -18989 147748 -18945
rect 147804 -18989 147848 -18945
rect 147904 -18989 147948 -18945
rect 148004 -18989 148048 -18945
rect 148104 -18989 148148 -18945
rect 148204 -18989 148248 -18945
rect 148304 -18989 148348 -18945
rect 148404 -18989 148448 -18945
rect 148904 -18989 148948 -18945
rect 149004 -18989 149048 -18945
rect 149104 -18989 149148 -18945
rect 149204 -18989 149248 -18945
rect 149304 -18989 149348 -18945
rect 149404 -18989 149448 -18945
rect 149504 -18989 149548 -18945
rect 149604 -18989 149648 -18945
rect 149704 -18989 149748 -18945
rect 149804 -18989 149848 -18945
rect 149904 -18989 149948 -18945
rect 150004 -18989 150048 -18945
rect 150104 -18989 150148 -18945
rect 150204 -18989 150248 -18945
rect 150304 -18989 150348 -18945
rect 150404 -18989 150448 -18945
rect 150904 -18989 150948 -18945
rect 151004 -18989 151048 -18945
rect 151104 -18989 151148 -18945
rect 151204 -18989 151248 -18945
rect 151304 -18989 151348 -18945
rect 151404 -18989 151448 -18945
rect 151504 -18989 151548 -18945
rect 151604 -18989 151648 -18945
rect 151704 -18989 151748 -18945
rect 151804 -18989 151848 -18945
rect 151904 -18989 151948 -18945
rect 152004 -18989 152048 -18945
rect 152104 -18989 152148 -18945
rect 152204 -18989 152248 -18945
rect 152304 -18989 152348 -18945
rect 152404 -18989 152448 -18945
rect 80849 -24070 80893 -24026
rect 80949 -24070 80993 -24026
rect 81049 -24070 81093 -24026
rect 81149 -24070 81193 -24026
rect 81249 -24070 81293 -24026
rect 81349 -24070 81393 -24026
rect 81449 -24070 81493 -24026
rect 81549 -24070 81593 -24026
rect 81649 -24070 81693 -24026
rect 81749 -24070 81793 -24026
rect 81849 -24070 81893 -24026
rect 81949 -24070 81993 -24026
rect 82049 -24070 82093 -24026
rect 82149 -24070 82193 -24026
rect 82249 -24070 82293 -24026
rect 82349 -24070 82393 -24026
rect 82849 -24070 82893 -24026
rect 82949 -24070 82993 -24026
rect 83049 -24070 83093 -24026
rect 83149 -24070 83193 -24026
rect 83249 -24070 83293 -24026
rect 83349 -24070 83393 -24026
rect 83449 -24070 83493 -24026
rect 83549 -24070 83593 -24026
rect 83649 -24070 83693 -24026
rect 83749 -24070 83793 -24026
rect 83849 -24070 83893 -24026
rect 83949 -24070 83993 -24026
rect 84049 -24070 84093 -24026
rect 84149 -24070 84193 -24026
rect 84249 -24070 84293 -24026
rect 84349 -24070 84393 -24026
rect 84849 -24070 84893 -24026
rect 84949 -24070 84993 -24026
rect 85049 -24070 85093 -24026
rect 85149 -24070 85193 -24026
rect 85249 -24070 85293 -24026
rect 85349 -24070 85393 -24026
rect 85449 -24070 85493 -24026
rect 85549 -24070 85593 -24026
rect 85649 -24070 85693 -24026
rect 85749 -24070 85793 -24026
rect 85849 -24070 85893 -24026
rect 85949 -24070 85993 -24026
rect 86049 -24070 86093 -24026
rect 86149 -24070 86193 -24026
rect 86249 -24070 86293 -24026
rect 86349 -24070 86393 -24026
rect 86849 -24070 86893 -24026
rect 86949 -24070 86993 -24026
rect 87049 -24070 87093 -24026
rect 87149 -24070 87193 -24026
rect 87249 -24070 87293 -24026
rect 87349 -24070 87393 -24026
rect 87449 -24070 87493 -24026
rect 87549 -24070 87593 -24026
rect 87649 -24070 87693 -24026
rect 87749 -24070 87793 -24026
rect 87849 -24070 87893 -24026
rect 87949 -24070 87993 -24026
rect 88049 -24070 88093 -24026
rect 88149 -24070 88193 -24026
rect 88249 -24070 88293 -24026
rect 88349 -24070 88393 -24026
rect 80849 -24170 80893 -24126
rect 80949 -24170 80993 -24126
rect 81049 -24170 81093 -24126
rect 81149 -24170 81193 -24126
rect 81249 -24170 81293 -24126
rect 81349 -24170 81393 -24126
rect 81449 -24170 81493 -24126
rect 81549 -24170 81593 -24126
rect 81649 -24170 81693 -24126
rect 81749 -24170 81793 -24126
rect 81849 -24170 81893 -24126
rect 81949 -24170 81993 -24126
rect 82049 -24170 82093 -24126
rect 82149 -24170 82193 -24126
rect 82249 -24170 82293 -24126
rect 82349 -24170 82393 -24126
rect 82849 -24170 82893 -24126
rect 82949 -24170 82993 -24126
rect 83049 -24170 83093 -24126
rect 83149 -24170 83193 -24126
rect 83249 -24170 83293 -24126
rect 83349 -24170 83393 -24126
rect 83449 -24170 83493 -24126
rect 83549 -24170 83593 -24126
rect 83649 -24170 83693 -24126
rect 83749 -24170 83793 -24126
rect 83849 -24170 83893 -24126
rect 83949 -24170 83993 -24126
rect 84049 -24170 84093 -24126
rect 84149 -24170 84193 -24126
rect 84249 -24170 84293 -24126
rect 84349 -24170 84393 -24126
rect 84849 -24170 84893 -24126
rect 84949 -24170 84993 -24126
rect 85049 -24170 85093 -24126
rect 85149 -24170 85193 -24126
rect 85249 -24170 85293 -24126
rect 85349 -24170 85393 -24126
rect 85449 -24170 85493 -24126
rect 85549 -24170 85593 -24126
rect 85649 -24170 85693 -24126
rect 85749 -24170 85793 -24126
rect 85849 -24170 85893 -24126
rect 85949 -24170 85993 -24126
rect 86049 -24170 86093 -24126
rect 86149 -24170 86193 -24126
rect 86249 -24170 86293 -24126
rect 86349 -24170 86393 -24126
rect 86849 -24170 86893 -24126
rect 86949 -24170 86993 -24126
rect 87049 -24170 87093 -24126
rect 87149 -24170 87193 -24126
rect 87249 -24170 87293 -24126
rect 87349 -24170 87393 -24126
rect 87449 -24170 87493 -24126
rect 87549 -24170 87593 -24126
rect 87649 -24170 87693 -24126
rect 87749 -24170 87793 -24126
rect 87849 -24170 87893 -24126
rect 87949 -24170 87993 -24126
rect 88049 -24170 88093 -24126
rect 88149 -24170 88193 -24126
rect 88249 -24170 88293 -24126
rect 88349 -24170 88393 -24126
rect 80849 -24270 80893 -24226
rect 80949 -24270 80993 -24226
rect 81049 -24270 81093 -24226
rect 81149 -24270 81193 -24226
rect 81249 -24270 81293 -24226
rect 81349 -24270 81393 -24226
rect 81449 -24270 81493 -24226
rect 81549 -24270 81593 -24226
rect 81649 -24270 81693 -24226
rect 81749 -24270 81793 -24226
rect 81849 -24270 81893 -24226
rect 81949 -24270 81993 -24226
rect 82049 -24270 82093 -24226
rect 82149 -24270 82193 -24226
rect 82249 -24270 82293 -24226
rect 82349 -24270 82393 -24226
rect 82849 -24270 82893 -24226
rect 82949 -24270 82993 -24226
rect 83049 -24270 83093 -24226
rect 83149 -24270 83193 -24226
rect 83249 -24270 83293 -24226
rect 83349 -24270 83393 -24226
rect 83449 -24270 83493 -24226
rect 83549 -24270 83593 -24226
rect 83649 -24270 83693 -24226
rect 83749 -24270 83793 -24226
rect 83849 -24270 83893 -24226
rect 83949 -24270 83993 -24226
rect 84049 -24270 84093 -24226
rect 84149 -24270 84193 -24226
rect 84249 -24270 84293 -24226
rect 84349 -24270 84393 -24226
rect 84849 -24270 84893 -24226
rect 84949 -24270 84993 -24226
rect 85049 -24270 85093 -24226
rect 85149 -24270 85193 -24226
rect 85249 -24270 85293 -24226
rect 85349 -24270 85393 -24226
rect 85449 -24270 85493 -24226
rect 85549 -24270 85593 -24226
rect 85649 -24270 85693 -24226
rect 85749 -24270 85793 -24226
rect 85849 -24270 85893 -24226
rect 85949 -24270 85993 -24226
rect 86049 -24270 86093 -24226
rect 86149 -24270 86193 -24226
rect 86249 -24270 86293 -24226
rect 86349 -24270 86393 -24226
rect 86849 -24270 86893 -24226
rect 86949 -24270 86993 -24226
rect 87049 -24270 87093 -24226
rect 87149 -24270 87193 -24226
rect 87249 -24270 87293 -24226
rect 87349 -24270 87393 -24226
rect 87449 -24270 87493 -24226
rect 87549 -24270 87593 -24226
rect 87649 -24270 87693 -24226
rect 87749 -24270 87793 -24226
rect 87849 -24270 87893 -24226
rect 87949 -24270 87993 -24226
rect 88049 -24270 88093 -24226
rect 88149 -24270 88193 -24226
rect 88249 -24270 88293 -24226
rect 88349 -24270 88393 -24226
rect 109104 -24239 109148 -24195
rect 109204 -24239 109248 -24195
rect 109304 -24239 109348 -24195
rect 109404 -24239 109448 -24195
rect 109504 -24239 109548 -24195
rect 109604 -24239 109648 -24195
rect 109704 -24239 109748 -24195
rect 109804 -24239 109848 -24195
rect 109904 -24239 109948 -24195
rect 110004 -24239 110048 -24195
rect 110104 -24239 110148 -24195
rect 110204 -24239 110248 -24195
rect 110304 -24239 110348 -24195
rect 110404 -24239 110448 -24195
rect 110504 -24239 110548 -24195
rect 110604 -24239 110648 -24195
rect 111104 -24239 111148 -24195
rect 111204 -24239 111248 -24195
rect 111304 -24239 111348 -24195
rect 111404 -24239 111448 -24195
rect 111504 -24239 111548 -24195
rect 111604 -24239 111648 -24195
rect 111704 -24239 111748 -24195
rect 111804 -24239 111848 -24195
rect 111904 -24239 111948 -24195
rect 112004 -24239 112048 -24195
rect 112104 -24239 112148 -24195
rect 112204 -24239 112248 -24195
rect 112304 -24239 112348 -24195
rect 112404 -24239 112448 -24195
rect 112504 -24239 112548 -24195
rect 112604 -24239 112648 -24195
rect 113104 -24239 113148 -24195
rect 113204 -24239 113248 -24195
rect 113304 -24239 113348 -24195
rect 113404 -24239 113448 -24195
rect 113504 -24239 113548 -24195
rect 113604 -24239 113648 -24195
rect 113704 -24239 113748 -24195
rect 113804 -24239 113848 -24195
rect 113904 -24239 113948 -24195
rect 114004 -24239 114048 -24195
rect 114104 -24239 114148 -24195
rect 114204 -24239 114248 -24195
rect 114304 -24239 114348 -24195
rect 114404 -24239 114448 -24195
rect 114504 -24239 114548 -24195
rect 114604 -24239 114648 -24195
rect 115104 -24239 115148 -24195
rect 115204 -24239 115248 -24195
rect 115304 -24239 115348 -24195
rect 115404 -24239 115448 -24195
rect 115504 -24239 115548 -24195
rect 115604 -24239 115648 -24195
rect 115704 -24239 115748 -24195
rect 115804 -24239 115848 -24195
rect 115904 -24239 115948 -24195
rect 116004 -24239 116048 -24195
rect 116104 -24239 116148 -24195
rect 116204 -24239 116248 -24195
rect 116304 -24239 116348 -24195
rect 116404 -24239 116448 -24195
rect 116504 -24239 116548 -24195
rect 116604 -24239 116648 -24195
rect -82799 -24410 -82755 -24366
rect -82699 -24410 -82655 -24366
rect -82599 -24410 -82555 -24366
rect -82499 -24410 -82455 -24366
rect -82399 -24410 -82355 -24366
rect -82299 -24410 -82255 -24366
rect -82199 -24410 -82155 -24366
rect -82099 -24410 -82055 -24366
rect -81999 -24410 -81955 -24366
rect -81899 -24410 -81855 -24366
rect -81799 -24410 -81755 -24366
rect -81699 -24410 -81655 -24366
rect -81599 -24410 -81555 -24366
rect -81499 -24410 -81455 -24366
rect -81399 -24410 -81355 -24366
rect -81299 -24410 -81255 -24366
rect -80799 -24410 -80755 -24366
rect -80699 -24410 -80655 -24366
rect -80599 -24410 -80555 -24366
rect -80499 -24410 -80455 -24366
rect -80399 -24410 -80355 -24366
rect -80299 -24410 -80255 -24366
rect -80199 -24410 -80155 -24366
rect -80099 -24410 -80055 -24366
rect -79999 -24410 -79955 -24366
rect -79899 -24410 -79855 -24366
rect -79799 -24410 -79755 -24366
rect -79699 -24410 -79655 -24366
rect -79599 -24410 -79555 -24366
rect -79499 -24410 -79455 -24366
rect -79399 -24410 -79355 -24366
rect -79299 -24410 -79255 -24366
rect -78799 -24410 -78755 -24366
rect -78699 -24410 -78655 -24366
rect -78599 -24410 -78555 -24366
rect -78499 -24410 -78455 -24366
rect -78399 -24410 -78355 -24366
rect -78299 -24410 -78255 -24366
rect -78199 -24410 -78155 -24366
rect -78099 -24410 -78055 -24366
rect -77999 -24410 -77955 -24366
rect -77899 -24410 -77855 -24366
rect -77799 -24410 -77755 -24366
rect -77699 -24410 -77655 -24366
rect -77599 -24410 -77555 -24366
rect -77499 -24410 -77455 -24366
rect -77399 -24410 -77355 -24366
rect -77299 -24410 -77255 -24366
rect -76799 -24410 -76755 -24366
rect -76699 -24410 -76655 -24366
rect -76599 -24410 -76555 -24366
rect -76499 -24410 -76455 -24366
rect -76399 -24410 -76355 -24366
rect -76299 -24410 -76255 -24366
rect -76199 -24410 -76155 -24366
rect -76099 -24410 -76055 -24366
rect -75999 -24410 -75955 -24366
rect -75899 -24410 -75855 -24366
rect -75799 -24410 -75755 -24366
rect -75699 -24410 -75655 -24366
rect -75599 -24410 -75555 -24366
rect -75499 -24410 -75455 -24366
rect -75399 -24410 -75355 -24366
rect -75299 -24410 -75255 -24366
rect 80849 -24370 80893 -24326
rect 80949 -24370 80993 -24326
rect 81049 -24370 81093 -24326
rect 81149 -24370 81193 -24326
rect 81249 -24370 81293 -24326
rect 81349 -24370 81393 -24326
rect 81449 -24370 81493 -24326
rect 81549 -24370 81593 -24326
rect 81649 -24370 81693 -24326
rect 81749 -24370 81793 -24326
rect 81849 -24370 81893 -24326
rect 81949 -24370 81993 -24326
rect 82049 -24370 82093 -24326
rect 82149 -24370 82193 -24326
rect 82249 -24370 82293 -24326
rect 82349 -24370 82393 -24326
rect 82849 -24370 82893 -24326
rect 82949 -24370 82993 -24326
rect 83049 -24370 83093 -24326
rect 83149 -24370 83193 -24326
rect 83249 -24370 83293 -24326
rect 83349 -24370 83393 -24326
rect 83449 -24370 83493 -24326
rect 83549 -24370 83593 -24326
rect 83649 -24370 83693 -24326
rect 83749 -24370 83793 -24326
rect 83849 -24370 83893 -24326
rect 83949 -24370 83993 -24326
rect 84049 -24370 84093 -24326
rect 84149 -24370 84193 -24326
rect 84249 -24370 84293 -24326
rect 84349 -24370 84393 -24326
rect 84849 -24370 84893 -24326
rect 84949 -24370 84993 -24326
rect 85049 -24370 85093 -24326
rect 85149 -24370 85193 -24326
rect 85249 -24370 85293 -24326
rect 85349 -24370 85393 -24326
rect 85449 -24370 85493 -24326
rect 85549 -24370 85593 -24326
rect 85649 -24370 85693 -24326
rect 85749 -24370 85793 -24326
rect 85849 -24370 85893 -24326
rect 85949 -24370 85993 -24326
rect 86049 -24370 86093 -24326
rect 86149 -24370 86193 -24326
rect 86249 -24370 86293 -24326
rect 86349 -24370 86393 -24326
rect 86849 -24370 86893 -24326
rect 86949 -24370 86993 -24326
rect 87049 -24370 87093 -24326
rect 87149 -24370 87193 -24326
rect 87249 -24370 87293 -24326
rect 87349 -24370 87393 -24326
rect 87449 -24370 87493 -24326
rect 87549 -24370 87593 -24326
rect 87649 -24370 87693 -24326
rect 87749 -24370 87793 -24326
rect 87849 -24370 87893 -24326
rect 87949 -24370 87993 -24326
rect 88049 -24370 88093 -24326
rect 88149 -24370 88193 -24326
rect 88249 -24370 88293 -24326
rect 88349 -24370 88393 -24326
rect 109104 -24339 109148 -24295
rect 109204 -24339 109248 -24295
rect 109304 -24339 109348 -24295
rect 109404 -24339 109448 -24295
rect 109504 -24339 109548 -24295
rect 109604 -24339 109648 -24295
rect 109704 -24339 109748 -24295
rect 109804 -24339 109848 -24295
rect 109904 -24339 109948 -24295
rect 110004 -24339 110048 -24295
rect 110104 -24339 110148 -24295
rect 110204 -24339 110248 -24295
rect 110304 -24339 110348 -24295
rect 110404 -24339 110448 -24295
rect 110504 -24339 110548 -24295
rect 110604 -24339 110648 -24295
rect 111104 -24339 111148 -24295
rect 111204 -24339 111248 -24295
rect 111304 -24339 111348 -24295
rect 111404 -24339 111448 -24295
rect 111504 -24339 111548 -24295
rect 111604 -24339 111648 -24295
rect 111704 -24339 111748 -24295
rect 111804 -24339 111848 -24295
rect 111904 -24339 111948 -24295
rect 112004 -24339 112048 -24295
rect 112104 -24339 112148 -24295
rect 112204 -24339 112248 -24295
rect 112304 -24339 112348 -24295
rect 112404 -24339 112448 -24295
rect 112504 -24339 112548 -24295
rect 112604 -24339 112648 -24295
rect 113104 -24339 113148 -24295
rect 113204 -24339 113248 -24295
rect 113304 -24339 113348 -24295
rect 113404 -24339 113448 -24295
rect 113504 -24339 113548 -24295
rect 113604 -24339 113648 -24295
rect 113704 -24339 113748 -24295
rect 113804 -24339 113848 -24295
rect 113904 -24339 113948 -24295
rect 114004 -24339 114048 -24295
rect 114104 -24339 114148 -24295
rect 114204 -24339 114248 -24295
rect 114304 -24339 114348 -24295
rect 114404 -24339 114448 -24295
rect 114504 -24339 114548 -24295
rect 114604 -24339 114648 -24295
rect 115104 -24339 115148 -24295
rect 115204 -24339 115248 -24295
rect 115304 -24339 115348 -24295
rect 115404 -24339 115448 -24295
rect 115504 -24339 115548 -24295
rect 115604 -24339 115648 -24295
rect 115704 -24339 115748 -24295
rect 115804 -24339 115848 -24295
rect 115904 -24339 115948 -24295
rect 116004 -24339 116048 -24295
rect 116104 -24339 116148 -24295
rect 116204 -24339 116248 -24295
rect 116304 -24339 116348 -24295
rect 116404 -24339 116448 -24295
rect 116504 -24339 116548 -24295
rect 116604 -24339 116648 -24295
rect -82799 -24510 -82755 -24466
rect -82699 -24510 -82655 -24466
rect -82599 -24510 -82555 -24466
rect -82499 -24510 -82455 -24466
rect -82399 -24510 -82355 -24466
rect -82299 -24510 -82255 -24466
rect -82199 -24510 -82155 -24466
rect -82099 -24510 -82055 -24466
rect -81999 -24510 -81955 -24466
rect -81899 -24510 -81855 -24466
rect -81799 -24510 -81755 -24466
rect -81699 -24510 -81655 -24466
rect -81599 -24510 -81555 -24466
rect -81499 -24510 -81455 -24466
rect -81399 -24510 -81355 -24466
rect -81299 -24510 -81255 -24466
rect -80799 -24510 -80755 -24466
rect -80699 -24510 -80655 -24466
rect -80599 -24510 -80555 -24466
rect -80499 -24510 -80455 -24466
rect -80399 -24510 -80355 -24466
rect -80299 -24510 -80255 -24466
rect -80199 -24510 -80155 -24466
rect -80099 -24510 -80055 -24466
rect -79999 -24510 -79955 -24466
rect -79899 -24510 -79855 -24466
rect -79799 -24510 -79755 -24466
rect -79699 -24510 -79655 -24466
rect -79599 -24510 -79555 -24466
rect -79499 -24510 -79455 -24466
rect -79399 -24510 -79355 -24466
rect -79299 -24510 -79255 -24466
rect -78799 -24510 -78755 -24466
rect -78699 -24510 -78655 -24466
rect -78599 -24510 -78555 -24466
rect -78499 -24510 -78455 -24466
rect -78399 -24510 -78355 -24466
rect -78299 -24510 -78255 -24466
rect -78199 -24510 -78155 -24466
rect -78099 -24510 -78055 -24466
rect -77999 -24510 -77955 -24466
rect -77899 -24510 -77855 -24466
rect -77799 -24510 -77755 -24466
rect -77699 -24510 -77655 -24466
rect -77599 -24510 -77555 -24466
rect -77499 -24510 -77455 -24466
rect -77399 -24510 -77355 -24466
rect -77299 -24510 -77255 -24466
rect -76799 -24510 -76755 -24466
rect -76699 -24510 -76655 -24466
rect -76599 -24510 -76555 -24466
rect -76499 -24510 -76455 -24466
rect -76399 -24510 -76355 -24466
rect -76299 -24510 -76255 -24466
rect -76199 -24510 -76155 -24466
rect -76099 -24510 -76055 -24466
rect -75999 -24510 -75955 -24466
rect -75899 -24510 -75855 -24466
rect -75799 -24510 -75755 -24466
rect -75699 -24510 -75655 -24466
rect -75599 -24510 -75555 -24466
rect -75499 -24510 -75455 -24466
rect -75399 -24510 -75355 -24466
rect -75299 -24510 -75255 -24466
rect 80849 -24470 80893 -24426
rect 80949 -24470 80993 -24426
rect 81049 -24470 81093 -24426
rect 81149 -24470 81193 -24426
rect 81249 -24470 81293 -24426
rect 81349 -24470 81393 -24426
rect 81449 -24470 81493 -24426
rect 81549 -24470 81593 -24426
rect 81649 -24470 81693 -24426
rect 81749 -24470 81793 -24426
rect 81849 -24470 81893 -24426
rect 81949 -24470 81993 -24426
rect 82049 -24470 82093 -24426
rect 82149 -24470 82193 -24426
rect 82249 -24470 82293 -24426
rect 82349 -24470 82393 -24426
rect 82849 -24470 82893 -24426
rect 82949 -24470 82993 -24426
rect 83049 -24470 83093 -24426
rect 83149 -24470 83193 -24426
rect 83249 -24470 83293 -24426
rect 83349 -24470 83393 -24426
rect 83449 -24470 83493 -24426
rect 83549 -24470 83593 -24426
rect 83649 -24470 83693 -24426
rect 83749 -24470 83793 -24426
rect 83849 -24470 83893 -24426
rect 83949 -24470 83993 -24426
rect 84049 -24470 84093 -24426
rect 84149 -24470 84193 -24426
rect 84249 -24470 84293 -24426
rect 84349 -24470 84393 -24426
rect 84849 -24470 84893 -24426
rect 84949 -24470 84993 -24426
rect 85049 -24470 85093 -24426
rect 85149 -24470 85193 -24426
rect 85249 -24470 85293 -24426
rect 85349 -24470 85393 -24426
rect 85449 -24470 85493 -24426
rect 85549 -24470 85593 -24426
rect 85649 -24470 85693 -24426
rect 85749 -24470 85793 -24426
rect 85849 -24470 85893 -24426
rect 85949 -24470 85993 -24426
rect 86049 -24470 86093 -24426
rect 86149 -24470 86193 -24426
rect 86249 -24470 86293 -24426
rect 86349 -24470 86393 -24426
rect 86849 -24470 86893 -24426
rect 86949 -24470 86993 -24426
rect 87049 -24470 87093 -24426
rect 87149 -24470 87193 -24426
rect 87249 -24470 87293 -24426
rect 87349 -24470 87393 -24426
rect 87449 -24470 87493 -24426
rect 87549 -24470 87593 -24426
rect 87649 -24470 87693 -24426
rect 87749 -24470 87793 -24426
rect 87849 -24470 87893 -24426
rect 87949 -24470 87993 -24426
rect 88049 -24470 88093 -24426
rect 88149 -24470 88193 -24426
rect 88249 -24470 88293 -24426
rect 88349 -24470 88393 -24426
rect 109104 -24439 109148 -24395
rect 109204 -24439 109248 -24395
rect 109304 -24439 109348 -24395
rect 109404 -24439 109448 -24395
rect 109504 -24439 109548 -24395
rect 109604 -24439 109648 -24395
rect 109704 -24439 109748 -24395
rect 109804 -24439 109848 -24395
rect 109904 -24439 109948 -24395
rect 110004 -24439 110048 -24395
rect 110104 -24439 110148 -24395
rect 110204 -24439 110248 -24395
rect 110304 -24439 110348 -24395
rect 110404 -24439 110448 -24395
rect 110504 -24439 110548 -24395
rect 110604 -24439 110648 -24395
rect 111104 -24439 111148 -24395
rect 111204 -24439 111248 -24395
rect 111304 -24439 111348 -24395
rect 111404 -24439 111448 -24395
rect 111504 -24439 111548 -24395
rect 111604 -24439 111648 -24395
rect 111704 -24439 111748 -24395
rect 111804 -24439 111848 -24395
rect 111904 -24439 111948 -24395
rect 112004 -24439 112048 -24395
rect 112104 -24439 112148 -24395
rect 112204 -24439 112248 -24395
rect 112304 -24439 112348 -24395
rect 112404 -24439 112448 -24395
rect 112504 -24439 112548 -24395
rect 112604 -24439 112648 -24395
rect 113104 -24439 113148 -24395
rect 113204 -24439 113248 -24395
rect 113304 -24439 113348 -24395
rect 113404 -24439 113448 -24395
rect 113504 -24439 113548 -24395
rect 113604 -24439 113648 -24395
rect 113704 -24439 113748 -24395
rect 113804 -24439 113848 -24395
rect 113904 -24439 113948 -24395
rect 114004 -24439 114048 -24395
rect 114104 -24439 114148 -24395
rect 114204 -24439 114248 -24395
rect 114304 -24439 114348 -24395
rect 114404 -24439 114448 -24395
rect 114504 -24439 114548 -24395
rect 114604 -24439 114648 -24395
rect 115104 -24439 115148 -24395
rect 115204 -24439 115248 -24395
rect 115304 -24439 115348 -24395
rect 115404 -24439 115448 -24395
rect 115504 -24439 115548 -24395
rect 115604 -24439 115648 -24395
rect 115704 -24439 115748 -24395
rect 115804 -24439 115848 -24395
rect 115904 -24439 115948 -24395
rect 116004 -24439 116048 -24395
rect 116104 -24439 116148 -24395
rect 116204 -24439 116248 -24395
rect 116304 -24439 116348 -24395
rect 116404 -24439 116448 -24395
rect 116504 -24439 116548 -24395
rect 116604 -24439 116648 -24395
rect -82799 -24610 -82755 -24566
rect -82699 -24610 -82655 -24566
rect -82599 -24610 -82555 -24566
rect -82499 -24610 -82455 -24566
rect -82399 -24610 -82355 -24566
rect -82299 -24610 -82255 -24566
rect -82199 -24610 -82155 -24566
rect -82099 -24610 -82055 -24566
rect -81999 -24610 -81955 -24566
rect -81899 -24610 -81855 -24566
rect -81799 -24610 -81755 -24566
rect -81699 -24610 -81655 -24566
rect -81599 -24610 -81555 -24566
rect -81499 -24610 -81455 -24566
rect -81399 -24610 -81355 -24566
rect -81299 -24610 -81255 -24566
rect -80799 -24610 -80755 -24566
rect -80699 -24610 -80655 -24566
rect -80599 -24610 -80555 -24566
rect -80499 -24610 -80455 -24566
rect -80399 -24610 -80355 -24566
rect -80299 -24610 -80255 -24566
rect -80199 -24610 -80155 -24566
rect -80099 -24610 -80055 -24566
rect -79999 -24610 -79955 -24566
rect -79899 -24610 -79855 -24566
rect -79799 -24610 -79755 -24566
rect -79699 -24610 -79655 -24566
rect -79599 -24610 -79555 -24566
rect -79499 -24610 -79455 -24566
rect -79399 -24610 -79355 -24566
rect -79299 -24610 -79255 -24566
rect -78799 -24610 -78755 -24566
rect -78699 -24610 -78655 -24566
rect -78599 -24610 -78555 -24566
rect -78499 -24610 -78455 -24566
rect -78399 -24610 -78355 -24566
rect -78299 -24610 -78255 -24566
rect -78199 -24610 -78155 -24566
rect -78099 -24610 -78055 -24566
rect -77999 -24610 -77955 -24566
rect -77899 -24610 -77855 -24566
rect -77799 -24610 -77755 -24566
rect -77699 -24610 -77655 -24566
rect -77599 -24610 -77555 -24566
rect -77499 -24610 -77455 -24566
rect -77399 -24610 -77355 -24566
rect -77299 -24610 -77255 -24566
rect -76799 -24610 -76755 -24566
rect -76699 -24610 -76655 -24566
rect -76599 -24610 -76555 -24566
rect -76499 -24610 -76455 -24566
rect -76399 -24610 -76355 -24566
rect -76299 -24610 -76255 -24566
rect -76199 -24610 -76155 -24566
rect -76099 -24610 -76055 -24566
rect -75999 -24610 -75955 -24566
rect -75899 -24610 -75855 -24566
rect -75799 -24610 -75755 -24566
rect -75699 -24610 -75655 -24566
rect -75599 -24610 -75555 -24566
rect -75499 -24610 -75455 -24566
rect -75399 -24610 -75355 -24566
rect -75299 -24610 -75255 -24566
rect 80849 -24570 80893 -24526
rect 80949 -24570 80993 -24526
rect 81049 -24570 81093 -24526
rect 81149 -24570 81193 -24526
rect 81249 -24570 81293 -24526
rect 81349 -24570 81393 -24526
rect 81449 -24570 81493 -24526
rect 81549 -24570 81593 -24526
rect 81649 -24570 81693 -24526
rect 81749 -24570 81793 -24526
rect 81849 -24570 81893 -24526
rect 81949 -24570 81993 -24526
rect 82049 -24570 82093 -24526
rect 82149 -24570 82193 -24526
rect 82249 -24570 82293 -24526
rect 82349 -24570 82393 -24526
rect 82849 -24570 82893 -24526
rect 82949 -24570 82993 -24526
rect 83049 -24570 83093 -24526
rect 83149 -24570 83193 -24526
rect 83249 -24570 83293 -24526
rect 83349 -24570 83393 -24526
rect 83449 -24570 83493 -24526
rect 83549 -24570 83593 -24526
rect 83649 -24570 83693 -24526
rect 83749 -24570 83793 -24526
rect 83849 -24570 83893 -24526
rect 83949 -24570 83993 -24526
rect 84049 -24570 84093 -24526
rect 84149 -24570 84193 -24526
rect 84249 -24570 84293 -24526
rect 84349 -24570 84393 -24526
rect 84849 -24570 84893 -24526
rect 84949 -24570 84993 -24526
rect 85049 -24570 85093 -24526
rect 85149 -24570 85193 -24526
rect 85249 -24570 85293 -24526
rect 85349 -24570 85393 -24526
rect 85449 -24570 85493 -24526
rect 85549 -24570 85593 -24526
rect 85649 -24570 85693 -24526
rect 85749 -24570 85793 -24526
rect 85849 -24570 85893 -24526
rect 85949 -24570 85993 -24526
rect 86049 -24570 86093 -24526
rect 86149 -24570 86193 -24526
rect 86249 -24570 86293 -24526
rect 86349 -24570 86393 -24526
rect 86849 -24570 86893 -24526
rect 86949 -24570 86993 -24526
rect 87049 -24570 87093 -24526
rect 87149 -24570 87193 -24526
rect 87249 -24570 87293 -24526
rect 87349 -24570 87393 -24526
rect 87449 -24570 87493 -24526
rect 87549 -24570 87593 -24526
rect 87649 -24570 87693 -24526
rect 87749 -24570 87793 -24526
rect 87849 -24570 87893 -24526
rect 87949 -24570 87993 -24526
rect 88049 -24570 88093 -24526
rect 88149 -24570 88193 -24526
rect 88249 -24570 88293 -24526
rect 88349 -24570 88393 -24526
rect 109104 -24539 109148 -24495
rect 109204 -24539 109248 -24495
rect 109304 -24539 109348 -24495
rect 109404 -24539 109448 -24495
rect 109504 -24539 109548 -24495
rect 109604 -24539 109648 -24495
rect 109704 -24539 109748 -24495
rect 109804 -24539 109848 -24495
rect 109904 -24539 109948 -24495
rect 110004 -24539 110048 -24495
rect 110104 -24539 110148 -24495
rect 110204 -24539 110248 -24495
rect 110304 -24539 110348 -24495
rect 110404 -24539 110448 -24495
rect 110504 -24539 110548 -24495
rect 110604 -24539 110648 -24495
rect 111104 -24539 111148 -24495
rect 111204 -24539 111248 -24495
rect 111304 -24539 111348 -24495
rect 111404 -24539 111448 -24495
rect 111504 -24539 111548 -24495
rect 111604 -24539 111648 -24495
rect 111704 -24539 111748 -24495
rect 111804 -24539 111848 -24495
rect 111904 -24539 111948 -24495
rect 112004 -24539 112048 -24495
rect 112104 -24539 112148 -24495
rect 112204 -24539 112248 -24495
rect 112304 -24539 112348 -24495
rect 112404 -24539 112448 -24495
rect 112504 -24539 112548 -24495
rect 112604 -24539 112648 -24495
rect 113104 -24539 113148 -24495
rect 113204 -24539 113248 -24495
rect 113304 -24539 113348 -24495
rect 113404 -24539 113448 -24495
rect 113504 -24539 113548 -24495
rect 113604 -24539 113648 -24495
rect 113704 -24539 113748 -24495
rect 113804 -24539 113848 -24495
rect 113904 -24539 113948 -24495
rect 114004 -24539 114048 -24495
rect 114104 -24539 114148 -24495
rect 114204 -24539 114248 -24495
rect 114304 -24539 114348 -24495
rect 114404 -24539 114448 -24495
rect 114504 -24539 114548 -24495
rect 114604 -24539 114648 -24495
rect 115104 -24539 115148 -24495
rect 115204 -24539 115248 -24495
rect 115304 -24539 115348 -24495
rect 115404 -24539 115448 -24495
rect 115504 -24539 115548 -24495
rect 115604 -24539 115648 -24495
rect 115704 -24539 115748 -24495
rect 115804 -24539 115848 -24495
rect 115904 -24539 115948 -24495
rect 116004 -24539 116048 -24495
rect 116104 -24539 116148 -24495
rect 116204 -24539 116248 -24495
rect 116304 -24539 116348 -24495
rect 116404 -24539 116448 -24495
rect 116504 -24539 116548 -24495
rect 116604 -24539 116648 -24495
rect -82799 -24710 -82755 -24666
rect -82699 -24710 -82655 -24666
rect -82599 -24710 -82555 -24666
rect -82499 -24710 -82455 -24666
rect -82399 -24710 -82355 -24666
rect -82299 -24710 -82255 -24666
rect -82199 -24710 -82155 -24666
rect -82099 -24710 -82055 -24666
rect -81999 -24710 -81955 -24666
rect -81899 -24710 -81855 -24666
rect -81799 -24710 -81755 -24666
rect -81699 -24710 -81655 -24666
rect -81599 -24710 -81555 -24666
rect -81499 -24710 -81455 -24666
rect -81399 -24710 -81355 -24666
rect -81299 -24710 -81255 -24666
rect -80799 -24710 -80755 -24666
rect -80699 -24710 -80655 -24666
rect -80599 -24710 -80555 -24666
rect -80499 -24710 -80455 -24666
rect -80399 -24710 -80355 -24666
rect -80299 -24710 -80255 -24666
rect -80199 -24710 -80155 -24666
rect -80099 -24710 -80055 -24666
rect -79999 -24710 -79955 -24666
rect -79899 -24710 -79855 -24666
rect -79799 -24710 -79755 -24666
rect -79699 -24710 -79655 -24666
rect -79599 -24710 -79555 -24666
rect -79499 -24710 -79455 -24666
rect -79399 -24710 -79355 -24666
rect -79299 -24710 -79255 -24666
rect -78799 -24710 -78755 -24666
rect -78699 -24710 -78655 -24666
rect -78599 -24710 -78555 -24666
rect -78499 -24710 -78455 -24666
rect -78399 -24710 -78355 -24666
rect -78299 -24710 -78255 -24666
rect -78199 -24710 -78155 -24666
rect -78099 -24710 -78055 -24666
rect -77999 -24710 -77955 -24666
rect -77899 -24710 -77855 -24666
rect -77799 -24710 -77755 -24666
rect -77699 -24710 -77655 -24666
rect -77599 -24710 -77555 -24666
rect -77499 -24710 -77455 -24666
rect -77399 -24710 -77355 -24666
rect -77299 -24710 -77255 -24666
rect -76799 -24710 -76755 -24666
rect -76699 -24710 -76655 -24666
rect -76599 -24710 -76555 -24666
rect -76499 -24710 -76455 -24666
rect -76399 -24710 -76355 -24666
rect -76299 -24710 -76255 -24666
rect -76199 -24710 -76155 -24666
rect -76099 -24710 -76055 -24666
rect -75999 -24710 -75955 -24666
rect -75899 -24710 -75855 -24666
rect -75799 -24710 -75755 -24666
rect -75699 -24710 -75655 -24666
rect -75599 -24710 -75555 -24666
rect -75499 -24710 -75455 -24666
rect -75399 -24710 -75355 -24666
rect -75299 -24710 -75255 -24666
rect 80849 -24670 80893 -24626
rect 80949 -24670 80993 -24626
rect 81049 -24670 81093 -24626
rect 81149 -24670 81193 -24626
rect 81249 -24670 81293 -24626
rect 81349 -24670 81393 -24626
rect 81449 -24670 81493 -24626
rect 81549 -24670 81593 -24626
rect 81649 -24670 81693 -24626
rect 81749 -24670 81793 -24626
rect 81849 -24670 81893 -24626
rect 81949 -24670 81993 -24626
rect 82049 -24670 82093 -24626
rect 82149 -24670 82193 -24626
rect 82249 -24670 82293 -24626
rect 82349 -24670 82393 -24626
rect 82849 -24670 82893 -24626
rect 82949 -24670 82993 -24626
rect 83049 -24670 83093 -24626
rect 83149 -24670 83193 -24626
rect 83249 -24670 83293 -24626
rect 83349 -24670 83393 -24626
rect 83449 -24670 83493 -24626
rect 83549 -24670 83593 -24626
rect 83649 -24670 83693 -24626
rect 83749 -24670 83793 -24626
rect 83849 -24670 83893 -24626
rect 83949 -24670 83993 -24626
rect 84049 -24670 84093 -24626
rect 84149 -24670 84193 -24626
rect 84249 -24670 84293 -24626
rect 84349 -24670 84393 -24626
rect 84849 -24670 84893 -24626
rect 84949 -24670 84993 -24626
rect 85049 -24670 85093 -24626
rect 85149 -24670 85193 -24626
rect 85249 -24670 85293 -24626
rect 85349 -24670 85393 -24626
rect 85449 -24670 85493 -24626
rect 85549 -24670 85593 -24626
rect 85649 -24670 85693 -24626
rect 85749 -24670 85793 -24626
rect 85849 -24670 85893 -24626
rect 85949 -24670 85993 -24626
rect 86049 -24670 86093 -24626
rect 86149 -24670 86193 -24626
rect 86249 -24670 86293 -24626
rect 86349 -24670 86393 -24626
rect 86849 -24670 86893 -24626
rect 86949 -24670 86993 -24626
rect 87049 -24670 87093 -24626
rect 87149 -24670 87193 -24626
rect 87249 -24670 87293 -24626
rect 87349 -24670 87393 -24626
rect 87449 -24670 87493 -24626
rect 87549 -24670 87593 -24626
rect 87649 -24670 87693 -24626
rect 87749 -24670 87793 -24626
rect 87849 -24670 87893 -24626
rect 87949 -24670 87993 -24626
rect 88049 -24670 88093 -24626
rect 88149 -24670 88193 -24626
rect 88249 -24670 88293 -24626
rect 88349 -24670 88393 -24626
rect 109104 -24639 109148 -24595
rect 109204 -24639 109248 -24595
rect 109304 -24639 109348 -24595
rect 109404 -24639 109448 -24595
rect 109504 -24639 109548 -24595
rect 109604 -24639 109648 -24595
rect 109704 -24639 109748 -24595
rect 109804 -24639 109848 -24595
rect 109904 -24639 109948 -24595
rect 110004 -24639 110048 -24595
rect 110104 -24639 110148 -24595
rect 110204 -24639 110248 -24595
rect 110304 -24639 110348 -24595
rect 110404 -24639 110448 -24595
rect 110504 -24639 110548 -24595
rect 110604 -24639 110648 -24595
rect 111104 -24639 111148 -24595
rect 111204 -24639 111248 -24595
rect 111304 -24639 111348 -24595
rect 111404 -24639 111448 -24595
rect 111504 -24639 111548 -24595
rect 111604 -24639 111648 -24595
rect 111704 -24639 111748 -24595
rect 111804 -24639 111848 -24595
rect 111904 -24639 111948 -24595
rect 112004 -24639 112048 -24595
rect 112104 -24639 112148 -24595
rect 112204 -24639 112248 -24595
rect 112304 -24639 112348 -24595
rect 112404 -24639 112448 -24595
rect 112504 -24639 112548 -24595
rect 112604 -24639 112648 -24595
rect 113104 -24639 113148 -24595
rect 113204 -24639 113248 -24595
rect 113304 -24639 113348 -24595
rect 113404 -24639 113448 -24595
rect 113504 -24639 113548 -24595
rect 113604 -24639 113648 -24595
rect 113704 -24639 113748 -24595
rect 113804 -24639 113848 -24595
rect 113904 -24639 113948 -24595
rect 114004 -24639 114048 -24595
rect 114104 -24639 114148 -24595
rect 114204 -24639 114248 -24595
rect 114304 -24639 114348 -24595
rect 114404 -24639 114448 -24595
rect 114504 -24639 114548 -24595
rect 114604 -24639 114648 -24595
rect 115104 -24639 115148 -24595
rect 115204 -24639 115248 -24595
rect 115304 -24639 115348 -24595
rect 115404 -24639 115448 -24595
rect 115504 -24639 115548 -24595
rect 115604 -24639 115648 -24595
rect 115704 -24639 115748 -24595
rect 115804 -24639 115848 -24595
rect 115904 -24639 115948 -24595
rect 116004 -24639 116048 -24595
rect 116104 -24639 116148 -24595
rect 116204 -24639 116248 -24595
rect 116304 -24639 116348 -24595
rect 116404 -24639 116448 -24595
rect 116504 -24639 116548 -24595
rect 116604 -24639 116648 -24595
rect -82799 -24810 -82755 -24766
rect -82699 -24810 -82655 -24766
rect -82599 -24810 -82555 -24766
rect -82499 -24810 -82455 -24766
rect -82399 -24810 -82355 -24766
rect -82299 -24810 -82255 -24766
rect -82199 -24810 -82155 -24766
rect -82099 -24810 -82055 -24766
rect -81999 -24810 -81955 -24766
rect -81899 -24810 -81855 -24766
rect -81799 -24810 -81755 -24766
rect -81699 -24810 -81655 -24766
rect -81599 -24810 -81555 -24766
rect -81499 -24810 -81455 -24766
rect -81399 -24810 -81355 -24766
rect -81299 -24810 -81255 -24766
rect -80799 -24810 -80755 -24766
rect -80699 -24810 -80655 -24766
rect -80599 -24810 -80555 -24766
rect -80499 -24810 -80455 -24766
rect -80399 -24810 -80355 -24766
rect -80299 -24810 -80255 -24766
rect -80199 -24810 -80155 -24766
rect -80099 -24810 -80055 -24766
rect -79999 -24810 -79955 -24766
rect -79899 -24810 -79855 -24766
rect -79799 -24810 -79755 -24766
rect -79699 -24810 -79655 -24766
rect -79599 -24810 -79555 -24766
rect -79499 -24810 -79455 -24766
rect -79399 -24810 -79355 -24766
rect -79299 -24810 -79255 -24766
rect -78799 -24810 -78755 -24766
rect -78699 -24810 -78655 -24766
rect -78599 -24810 -78555 -24766
rect -78499 -24810 -78455 -24766
rect -78399 -24810 -78355 -24766
rect -78299 -24810 -78255 -24766
rect -78199 -24810 -78155 -24766
rect -78099 -24810 -78055 -24766
rect -77999 -24810 -77955 -24766
rect -77899 -24810 -77855 -24766
rect -77799 -24810 -77755 -24766
rect -77699 -24810 -77655 -24766
rect -77599 -24810 -77555 -24766
rect -77499 -24810 -77455 -24766
rect -77399 -24810 -77355 -24766
rect -77299 -24810 -77255 -24766
rect -76799 -24810 -76755 -24766
rect -76699 -24810 -76655 -24766
rect -76599 -24810 -76555 -24766
rect -76499 -24810 -76455 -24766
rect -76399 -24810 -76355 -24766
rect -76299 -24810 -76255 -24766
rect -76199 -24810 -76155 -24766
rect -76099 -24810 -76055 -24766
rect -75999 -24810 -75955 -24766
rect -75899 -24810 -75855 -24766
rect -75799 -24810 -75755 -24766
rect -75699 -24810 -75655 -24766
rect -75599 -24810 -75555 -24766
rect -75499 -24810 -75455 -24766
rect -75399 -24810 -75355 -24766
rect -75299 -24810 -75255 -24766
rect 80849 -24770 80893 -24726
rect 80949 -24770 80993 -24726
rect 81049 -24770 81093 -24726
rect 81149 -24770 81193 -24726
rect 81249 -24770 81293 -24726
rect 81349 -24770 81393 -24726
rect 81449 -24770 81493 -24726
rect 81549 -24770 81593 -24726
rect 81649 -24770 81693 -24726
rect 81749 -24770 81793 -24726
rect 81849 -24770 81893 -24726
rect 81949 -24770 81993 -24726
rect 82049 -24770 82093 -24726
rect 82149 -24770 82193 -24726
rect 82249 -24770 82293 -24726
rect 82349 -24770 82393 -24726
rect 82849 -24770 82893 -24726
rect 82949 -24770 82993 -24726
rect 83049 -24770 83093 -24726
rect 83149 -24770 83193 -24726
rect 83249 -24770 83293 -24726
rect 83349 -24770 83393 -24726
rect 83449 -24770 83493 -24726
rect 83549 -24770 83593 -24726
rect 83649 -24770 83693 -24726
rect 83749 -24770 83793 -24726
rect 83849 -24770 83893 -24726
rect 83949 -24770 83993 -24726
rect 84049 -24770 84093 -24726
rect 84149 -24770 84193 -24726
rect 84249 -24770 84293 -24726
rect 84349 -24770 84393 -24726
rect 84849 -24770 84893 -24726
rect 84949 -24770 84993 -24726
rect 85049 -24770 85093 -24726
rect 85149 -24770 85193 -24726
rect 85249 -24770 85293 -24726
rect 85349 -24770 85393 -24726
rect 85449 -24770 85493 -24726
rect 85549 -24770 85593 -24726
rect 85649 -24770 85693 -24726
rect 85749 -24770 85793 -24726
rect 85849 -24770 85893 -24726
rect 85949 -24770 85993 -24726
rect 86049 -24770 86093 -24726
rect 86149 -24770 86193 -24726
rect 86249 -24770 86293 -24726
rect 86349 -24770 86393 -24726
rect 86849 -24770 86893 -24726
rect 86949 -24770 86993 -24726
rect 87049 -24770 87093 -24726
rect 87149 -24770 87193 -24726
rect 87249 -24770 87293 -24726
rect 87349 -24770 87393 -24726
rect 87449 -24770 87493 -24726
rect 87549 -24770 87593 -24726
rect 87649 -24770 87693 -24726
rect 87749 -24770 87793 -24726
rect 87849 -24770 87893 -24726
rect 87949 -24770 87993 -24726
rect 88049 -24770 88093 -24726
rect 88149 -24770 88193 -24726
rect 88249 -24770 88293 -24726
rect 88349 -24770 88393 -24726
rect 109104 -24739 109148 -24695
rect 109204 -24739 109248 -24695
rect 109304 -24739 109348 -24695
rect 109404 -24739 109448 -24695
rect 109504 -24739 109548 -24695
rect 109604 -24739 109648 -24695
rect 109704 -24739 109748 -24695
rect 109804 -24739 109848 -24695
rect 109904 -24739 109948 -24695
rect 110004 -24739 110048 -24695
rect 110104 -24739 110148 -24695
rect 110204 -24739 110248 -24695
rect 110304 -24739 110348 -24695
rect 110404 -24739 110448 -24695
rect 110504 -24739 110548 -24695
rect 110604 -24739 110648 -24695
rect 111104 -24739 111148 -24695
rect 111204 -24739 111248 -24695
rect 111304 -24739 111348 -24695
rect 111404 -24739 111448 -24695
rect 111504 -24739 111548 -24695
rect 111604 -24739 111648 -24695
rect 111704 -24739 111748 -24695
rect 111804 -24739 111848 -24695
rect 111904 -24739 111948 -24695
rect 112004 -24739 112048 -24695
rect 112104 -24739 112148 -24695
rect 112204 -24739 112248 -24695
rect 112304 -24739 112348 -24695
rect 112404 -24739 112448 -24695
rect 112504 -24739 112548 -24695
rect 112604 -24739 112648 -24695
rect 113104 -24739 113148 -24695
rect 113204 -24739 113248 -24695
rect 113304 -24739 113348 -24695
rect 113404 -24739 113448 -24695
rect 113504 -24739 113548 -24695
rect 113604 -24739 113648 -24695
rect 113704 -24739 113748 -24695
rect 113804 -24739 113848 -24695
rect 113904 -24739 113948 -24695
rect 114004 -24739 114048 -24695
rect 114104 -24739 114148 -24695
rect 114204 -24739 114248 -24695
rect 114304 -24739 114348 -24695
rect 114404 -24739 114448 -24695
rect 114504 -24739 114548 -24695
rect 114604 -24739 114648 -24695
rect 115104 -24739 115148 -24695
rect 115204 -24739 115248 -24695
rect 115304 -24739 115348 -24695
rect 115404 -24739 115448 -24695
rect 115504 -24739 115548 -24695
rect 115604 -24739 115648 -24695
rect 115704 -24739 115748 -24695
rect 115804 -24739 115848 -24695
rect 115904 -24739 115948 -24695
rect 116004 -24739 116048 -24695
rect 116104 -24739 116148 -24695
rect 116204 -24739 116248 -24695
rect 116304 -24739 116348 -24695
rect 116404 -24739 116448 -24695
rect 116504 -24739 116548 -24695
rect 116604 -24739 116648 -24695
rect -82799 -24910 -82755 -24866
rect -82699 -24910 -82655 -24866
rect -82599 -24910 -82555 -24866
rect -82499 -24910 -82455 -24866
rect -82399 -24910 -82355 -24866
rect -82299 -24910 -82255 -24866
rect -82199 -24910 -82155 -24866
rect -82099 -24910 -82055 -24866
rect -81999 -24910 -81955 -24866
rect -81899 -24910 -81855 -24866
rect -81799 -24910 -81755 -24866
rect -81699 -24910 -81655 -24866
rect -81599 -24910 -81555 -24866
rect -81499 -24910 -81455 -24866
rect -81399 -24910 -81355 -24866
rect -81299 -24910 -81255 -24866
rect -80799 -24910 -80755 -24866
rect -80699 -24910 -80655 -24866
rect -80599 -24910 -80555 -24866
rect -80499 -24910 -80455 -24866
rect -80399 -24910 -80355 -24866
rect -80299 -24910 -80255 -24866
rect -80199 -24910 -80155 -24866
rect -80099 -24910 -80055 -24866
rect -79999 -24910 -79955 -24866
rect -79899 -24910 -79855 -24866
rect -79799 -24910 -79755 -24866
rect -79699 -24910 -79655 -24866
rect -79599 -24910 -79555 -24866
rect -79499 -24910 -79455 -24866
rect -79399 -24910 -79355 -24866
rect -79299 -24910 -79255 -24866
rect -78799 -24910 -78755 -24866
rect -78699 -24910 -78655 -24866
rect -78599 -24910 -78555 -24866
rect -78499 -24910 -78455 -24866
rect -78399 -24910 -78355 -24866
rect -78299 -24910 -78255 -24866
rect -78199 -24910 -78155 -24866
rect -78099 -24910 -78055 -24866
rect -77999 -24910 -77955 -24866
rect -77899 -24910 -77855 -24866
rect -77799 -24910 -77755 -24866
rect -77699 -24910 -77655 -24866
rect -77599 -24910 -77555 -24866
rect -77499 -24910 -77455 -24866
rect -77399 -24910 -77355 -24866
rect -77299 -24910 -77255 -24866
rect -76799 -24910 -76755 -24866
rect -76699 -24910 -76655 -24866
rect -76599 -24910 -76555 -24866
rect -76499 -24910 -76455 -24866
rect -76399 -24910 -76355 -24866
rect -76299 -24910 -76255 -24866
rect -76199 -24910 -76155 -24866
rect -76099 -24910 -76055 -24866
rect -75999 -24910 -75955 -24866
rect -75899 -24910 -75855 -24866
rect -75799 -24910 -75755 -24866
rect -75699 -24910 -75655 -24866
rect -75599 -24910 -75555 -24866
rect -75499 -24910 -75455 -24866
rect -75399 -24910 -75355 -24866
rect -75299 -24910 -75255 -24866
rect 80849 -24870 80893 -24826
rect 80949 -24870 80993 -24826
rect 81049 -24870 81093 -24826
rect 81149 -24870 81193 -24826
rect 81249 -24870 81293 -24826
rect 81349 -24870 81393 -24826
rect 81449 -24870 81493 -24826
rect 81549 -24870 81593 -24826
rect 81649 -24870 81693 -24826
rect 81749 -24870 81793 -24826
rect 81849 -24870 81893 -24826
rect 81949 -24870 81993 -24826
rect 82049 -24870 82093 -24826
rect 82149 -24870 82193 -24826
rect 82249 -24870 82293 -24826
rect 82349 -24870 82393 -24826
rect 82849 -24870 82893 -24826
rect 82949 -24870 82993 -24826
rect 83049 -24870 83093 -24826
rect 83149 -24870 83193 -24826
rect 83249 -24870 83293 -24826
rect 83349 -24870 83393 -24826
rect 83449 -24870 83493 -24826
rect 83549 -24870 83593 -24826
rect 83649 -24870 83693 -24826
rect 83749 -24870 83793 -24826
rect 83849 -24870 83893 -24826
rect 83949 -24870 83993 -24826
rect 84049 -24870 84093 -24826
rect 84149 -24870 84193 -24826
rect 84249 -24870 84293 -24826
rect 84349 -24870 84393 -24826
rect 84849 -24870 84893 -24826
rect 84949 -24870 84993 -24826
rect 85049 -24870 85093 -24826
rect 85149 -24870 85193 -24826
rect 85249 -24870 85293 -24826
rect 85349 -24870 85393 -24826
rect 85449 -24870 85493 -24826
rect 85549 -24870 85593 -24826
rect 85649 -24870 85693 -24826
rect 85749 -24870 85793 -24826
rect 85849 -24870 85893 -24826
rect 85949 -24870 85993 -24826
rect 86049 -24870 86093 -24826
rect 86149 -24870 86193 -24826
rect 86249 -24870 86293 -24826
rect 86349 -24870 86393 -24826
rect 86849 -24870 86893 -24826
rect 86949 -24870 86993 -24826
rect 87049 -24870 87093 -24826
rect 87149 -24870 87193 -24826
rect 87249 -24870 87293 -24826
rect 87349 -24870 87393 -24826
rect 87449 -24870 87493 -24826
rect 87549 -24870 87593 -24826
rect 87649 -24870 87693 -24826
rect 87749 -24870 87793 -24826
rect 87849 -24870 87893 -24826
rect 87949 -24870 87993 -24826
rect 88049 -24870 88093 -24826
rect 88149 -24870 88193 -24826
rect 88249 -24870 88293 -24826
rect 88349 -24870 88393 -24826
rect 109104 -24839 109148 -24795
rect 109204 -24839 109248 -24795
rect 109304 -24839 109348 -24795
rect 109404 -24839 109448 -24795
rect 109504 -24839 109548 -24795
rect 109604 -24839 109648 -24795
rect 109704 -24839 109748 -24795
rect 109804 -24839 109848 -24795
rect 109904 -24839 109948 -24795
rect 110004 -24839 110048 -24795
rect 110104 -24839 110148 -24795
rect 110204 -24839 110248 -24795
rect 110304 -24839 110348 -24795
rect 110404 -24839 110448 -24795
rect 110504 -24839 110548 -24795
rect 110604 -24839 110648 -24795
rect 111104 -24839 111148 -24795
rect 111204 -24839 111248 -24795
rect 111304 -24839 111348 -24795
rect 111404 -24839 111448 -24795
rect 111504 -24839 111548 -24795
rect 111604 -24839 111648 -24795
rect 111704 -24839 111748 -24795
rect 111804 -24839 111848 -24795
rect 111904 -24839 111948 -24795
rect 112004 -24839 112048 -24795
rect 112104 -24839 112148 -24795
rect 112204 -24839 112248 -24795
rect 112304 -24839 112348 -24795
rect 112404 -24839 112448 -24795
rect 112504 -24839 112548 -24795
rect 112604 -24839 112648 -24795
rect 113104 -24839 113148 -24795
rect 113204 -24839 113248 -24795
rect 113304 -24839 113348 -24795
rect 113404 -24839 113448 -24795
rect 113504 -24839 113548 -24795
rect 113604 -24839 113648 -24795
rect 113704 -24839 113748 -24795
rect 113804 -24839 113848 -24795
rect 113904 -24839 113948 -24795
rect 114004 -24839 114048 -24795
rect 114104 -24839 114148 -24795
rect 114204 -24839 114248 -24795
rect 114304 -24839 114348 -24795
rect 114404 -24839 114448 -24795
rect 114504 -24839 114548 -24795
rect 114604 -24839 114648 -24795
rect 115104 -24839 115148 -24795
rect 115204 -24839 115248 -24795
rect 115304 -24839 115348 -24795
rect 115404 -24839 115448 -24795
rect 115504 -24839 115548 -24795
rect 115604 -24839 115648 -24795
rect 115704 -24839 115748 -24795
rect 115804 -24839 115848 -24795
rect 115904 -24839 115948 -24795
rect 116004 -24839 116048 -24795
rect 116104 -24839 116148 -24795
rect 116204 -24839 116248 -24795
rect 116304 -24839 116348 -24795
rect 116404 -24839 116448 -24795
rect 116504 -24839 116548 -24795
rect 116604 -24839 116648 -24795
rect -82799 -25010 -82755 -24966
rect -82699 -25010 -82655 -24966
rect -82599 -25010 -82555 -24966
rect -82499 -25010 -82455 -24966
rect -82399 -25010 -82355 -24966
rect -82299 -25010 -82255 -24966
rect -82199 -25010 -82155 -24966
rect -82099 -25010 -82055 -24966
rect -81999 -25010 -81955 -24966
rect -81899 -25010 -81855 -24966
rect -81799 -25010 -81755 -24966
rect -81699 -25010 -81655 -24966
rect -81599 -25010 -81555 -24966
rect -81499 -25010 -81455 -24966
rect -81399 -25010 -81355 -24966
rect -81299 -25010 -81255 -24966
rect -80799 -25010 -80755 -24966
rect -80699 -25010 -80655 -24966
rect -80599 -25010 -80555 -24966
rect -80499 -25010 -80455 -24966
rect -80399 -25010 -80355 -24966
rect -80299 -25010 -80255 -24966
rect -80199 -25010 -80155 -24966
rect -80099 -25010 -80055 -24966
rect -79999 -25010 -79955 -24966
rect -79899 -25010 -79855 -24966
rect -79799 -25010 -79755 -24966
rect -79699 -25010 -79655 -24966
rect -79599 -25010 -79555 -24966
rect -79499 -25010 -79455 -24966
rect -79399 -25010 -79355 -24966
rect -79299 -25010 -79255 -24966
rect -78799 -25010 -78755 -24966
rect -78699 -25010 -78655 -24966
rect -78599 -25010 -78555 -24966
rect -78499 -25010 -78455 -24966
rect -78399 -25010 -78355 -24966
rect -78299 -25010 -78255 -24966
rect -78199 -25010 -78155 -24966
rect -78099 -25010 -78055 -24966
rect -77999 -25010 -77955 -24966
rect -77899 -25010 -77855 -24966
rect -77799 -25010 -77755 -24966
rect -77699 -25010 -77655 -24966
rect -77599 -25010 -77555 -24966
rect -77499 -25010 -77455 -24966
rect -77399 -25010 -77355 -24966
rect -77299 -25010 -77255 -24966
rect -76799 -25010 -76755 -24966
rect -76699 -25010 -76655 -24966
rect -76599 -25010 -76555 -24966
rect -76499 -25010 -76455 -24966
rect -76399 -25010 -76355 -24966
rect -76299 -25010 -76255 -24966
rect -76199 -25010 -76155 -24966
rect -76099 -25010 -76055 -24966
rect -75999 -25010 -75955 -24966
rect -75899 -25010 -75855 -24966
rect -75799 -25010 -75755 -24966
rect -75699 -25010 -75655 -24966
rect -75599 -25010 -75555 -24966
rect -75499 -25010 -75455 -24966
rect -75399 -25010 -75355 -24966
rect -75299 -25010 -75255 -24966
rect 80849 -24970 80893 -24926
rect 80949 -24970 80993 -24926
rect 81049 -24970 81093 -24926
rect 81149 -24970 81193 -24926
rect 81249 -24970 81293 -24926
rect 81349 -24970 81393 -24926
rect 81449 -24970 81493 -24926
rect 81549 -24970 81593 -24926
rect 81649 -24970 81693 -24926
rect 81749 -24970 81793 -24926
rect 81849 -24970 81893 -24926
rect 81949 -24970 81993 -24926
rect 82049 -24970 82093 -24926
rect 82149 -24970 82193 -24926
rect 82249 -24970 82293 -24926
rect 82349 -24970 82393 -24926
rect 82849 -24970 82893 -24926
rect 82949 -24970 82993 -24926
rect 83049 -24970 83093 -24926
rect 83149 -24970 83193 -24926
rect 83249 -24970 83293 -24926
rect 83349 -24970 83393 -24926
rect 83449 -24970 83493 -24926
rect 83549 -24970 83593 -24926
rect 83649 -24970 83693 -24926
rect 83749 -24970 83793 -24926
rect 83849 -24970 83893 -24926
rect 83949 -24970 83993 -24926
rect 84049 -24970 84093 -24926
rect 84149 -24970 84193 -24926
rect 84249 -24970 84293 -24926
rect 84349 -24970 84393 -24926
rect 84849 -24970 84893 -24926
rect 84949 -24970 84993 -24926
rect 85049 -24970 85093 -24926
rect 85149 -24970 85193 -24926
rect 85249 -24970 85293 -24926
rect 85349 -24970 85393 -24926
rect 85449 -24970 85493 -24926
rect 85549 -24970 85593 -24926
rect 85649 -24970 85693 -24926
rect 85749 -24970 85793 -24926
rect 85849 -24970 85893 -24926
rect 85949 -24970 85993 -24926
rect 86049 -24970 86093 -24926
rect 86149 -24970 86193 -24926
rect 86249 -24970 86293 -24926
rect 86349 -24970 86393 -24926
rect 86849 -24970 86893 -24926
rect 86949 -24970 86993 -24926
rect 87049 -24970 87093 -24926
rect 87149 -24970 87193 -24926
rect 87249 -24970 87293 -24926
rect 87349 -24970 87393 -24926
rect 87449 -24970 87493 -24926
rect 87549 -24970 87593 -24926
rect 87649 -24970 87693 -24926
rect 87749 -24970 87793 -24926
rect 87849 -24970 87893 -24926
rect 87949 -24970 87993 -24926
rect 88049 -24970 88093 -24926
rect 88149 -24970 88193 -24926
rect 88249 -24970 88293 -24926
rect 88349 -24970 88393 -24926
rect 109104 -24939 109148 -24895
rect 109204 -24939 109248 -24895
rect 109304 -24939 109348 -24895
rect 109404 -24939 109448 -24895
rect 109504 -24939 109548 -24895
rect 109604 -24939 109648 -24895
rect 109704 -24939 109748 -24895
rect 109804 -24939 109848 -24895
rect 109904 -24939 109948 -24895
rect 110004 -24939 110048 -24895
rect 110104 -24939 110148 -24895
rect 110204 -24939 110248 -24895
rect 110304 -24939 110348 -24895
rect 110404 -24939 110448 -24895
rect 110504 -24939 110548 -24895
rect 110604 -24939 110648 -24895
rect 111104 -24939 111148 -24895
rect 111204 -24939 111248 -24895
rect 111304 -24939 111348 -24895
rect 111404 -24939 111448 -24895
rect 111504 -24939 111548 -24895
rect 111604 -24939 111648 -24895
rect 111704 -24939 111748 -24895
rect 111804 -24939 111848 -24895
rect 111904 -24939 111948 -24895
rect 112004 -24939 112048 -24895
rect 112104 -24939 112148 -24895
rect 112204 -24939 112248 -24895
rect 112304 -24939 112348 -24895
rect 112404 -24939 112448 -24895
rect 112504 -24939 112548 -24895
rect 112604 -24939 112648 -24895
rect 113104 -24939 113148 -24895
rect 113204 -24939 113248 -24895
rect 113304 -24939 113348 -24895
rect 113404 -24939 113448 -24895
rect 113504 -24939 113548 -24895
rect 113604 -24939 113648 -24895
rect 113704 -24939 113748 -24895
rect 113804 -24939 113848 -24895
rect 113904 -24939 113948 -24895
rect 114004 -24939 114048 -24895
rect 114104 -24939 114148 -24895
rect 114204 -24939 114248 -24895
rect 114304 -24939 114348 -24895
rect 114404 -24939 114448 -24895
rect 114504 -24939 114548 -24895
rect 114604 -24939 114648 -24895
rect 115104 -24939 115148 -24895
rect 115204 -24939 115248 -24895
rect 115304 -24939 115348 -24895
rect 115404 -24939 115448 -24895
rect 115504 -24939 115548 -24895
rect 115604 -24939 115648 -24895
rect 115704 -24939 115748 -24895
rect 115804 -24939 115848 -24895
rect 115904 -24939 115948 -24895
rect 116004 -24939 116048 -24895
rect 116104 -24939 116148 -24895
rect 116204 -24939 116248 -24895
rect 116304 -24939 116348 -24895
rect 116404 -24939 116448 -24895
rect 116504 -24939 116548 -24895
rect 116604 -24939 116648 -24895
rect -82799 -25110 -82755 -25066
rect -82699 -25110 -82655 -25066
rect -82599 -25110 -82555 -25066
rect -82499 -25110 -82455 -25066
rect -82399 -25110 -82355 -25066
rect -82299 -25110 -82255 -25066
rect -82199 -25110 -82155 -25066
rect -82099 -25110 -82055 -25066
rect -81999 -25110 -81955 -25066
rect -81899 -25110 -81855 -25066
rect -81799 -25110 -81755 -25066
rect -81699 -25110 -81655 -25066
rect -81599 -25110 -81555 -25066
rect -81499 -25110 -81455 -25066
rect -81399 -25110 -81355 -25066
rect -81299 -25110 -81255 -25066
rect -80799 -25110 -80755 -25066
rect -80699 -25110 -80655 -25066
rect -80599 -25110 -80555 -25066
rect -80499 -25110 -80455 -25066
rect -80399 -25110 -80355 -25066
rect -80299 -25110 -80255 -25066
rect -80199 -25110 -80155 -25066
rect -80099 -25110 -80055 -25066
rect -79999 -25110 -79955 -25066
rect -79899 -25110 -79855 -25066
rect -79799 -25110 -79755 -25066
rect -79699 -25110 -79655 -25066
rect -79599 -25110 -79555 -25066
rect -79499 -25110 -79455 -25066
rect -79399 -25110 -79355 -25066
rect -79299 -25110 -79255 -25066
rect -78799 -25110 -78755 -25066
rect -78699 -25110 -78655 -25066
rect -78599 -25110 -78555 -25066
rect -78499 -25110 -78455 -25066
rect -78399 -25110 -78355 -25066
rect -78299 -25110 -78255 -25066
rect -78199 -25110 -78155 -25066
rect -78099 -25110 -78055 -25066
rect -77999 -25110 -77955 -25066
rect -77899 -25110 -77855 -25066
rect -77799 -25110 -77755 -25066
rect -77699 -25110 -77655 -25066
rect -77599 -25110 -77555 -25066
rect -77499 -25110 -77455 -25066
rect -77399 -25110 -77355 -25066
rect -77299 -25110 -77255 -25066
rect -76799 -25110 -76755 -25066
rect -76699 -25110 -76655 -25066
rect -76599 -25110 -76555 -25066
rect -76499 -25110 -76455 -25066
rect -76399 -25110 -76355 -25066
rect -76299 -25110 -76255 -25066
rect -76199 -25110 -76155 -25066
rect -76099 -25110 -76055 -25066
rect -75999 -25110 -75955 -25066
rect -75899 -25110 -75855 -25066
rect -75799 -25110 -75755 -25066
rect -75699 -25110 -75655 -25066
rect -75599 -25110 -75555 -25066
rect -75499 -25110 -75455 -25066
rect -75399 -25110 -75355 -25066
rect -75299 -25110 -75255 -25066
rect 80849 -25070 80893 -25026
rect 80949 -25070 80993 -25026
rect 81049 -25070 81093 -25026
rect 81149 -25070 81193 -25026
rect 81249 -25070 81293 -25026
rect 81349 -25070 81393 -25026
rect 81449 -25070 81493 -25026
rect 81549 -25070 81593 -25026
rect 81649 -25070 81693 -25026
rect 81749 -25070 81793 -25026
rect 81849 -25070 81893 -25026
rect 81949 -25070 81993 -25026
rect 82049 -25070 82093 -25026
rect 82149 -25070 82193 -25026
rect 82249 -25070 82293 -25026
rect 82349 -25070 82393 -25026
rect 82849 -25070 82893 -25026
rect 82949 -25070 82993 -25026
rect 83049 -25070 83093 -25026
rect 83149 -25070 83193 -25026
rect 83249 -25070 83293 -25026
rect 83349 -25070 83393 -25026
rect 83449 -25070 83493 -25026
rect 83549 -25070 83593 -25026
rect 83649 -25070 83693 -25026
rect 83749 -25070 83793 -25026
rect 83849 -25070 83893 -25026
rect 83949 -25070 83993 -25026
rect 84049 -25070 84093 -25026
rect 84149 -25070 84193 -25026
rect 84249 -25070 84293 -25026
rect 84349 -25070 84393 -25026
rect 84849 -25070 84893 -25026
rect 84949 -25070 84993 -25026
rect 85049 -25070 85093 -25026
rect 85149 -25070 85193 -25026
rect 85249 -25070 85293 -25026
rect 85349 -25070 85393 -25026
rect 85449 -25070 85493 -25026
rect 85549 -25070 85593 -25026
rect 85649 -25070 85693 -25026
rect 85749 -25070 85793 -25026
rect 85849 -25070 85893 -25026
rect 85949 -25070 85993 -25026
rect 86049 -25070 86093 -25026
rect 86149 -25070 86193 -25026
rect 86249 -25070 86293 -25026
rect 86349 -25070 86393 -25026
rect 86849 -25070 86893 -25026
rect 86949 -25070 86993 -25026
rect 87049 -25070 87093 -25026
rect 87149 -25070 87193 -25026
rect 87249 -25070 87293 -25026
rect 87349 -25070 87393 -25026
rect 87449 -25070 87493 -25026
rect 87549 -25070 87593 -25026
rect 87649 -25070 87693 -25026
rect 87749 -25070 87793 -25026
rect 87849 -25070 87893 -25026
rect 87949 -25070 87993 -25026
rect 88049 -25070 88093 -25026
rect 88149 -25070 88193 -25026
rect 88249 -25070 88293 -25026
rect 88349 -25070 88393 -25026
rect 109104 -25039 109148 -24995
rect 109204 -25039 109248 -24995
rect 109304 -25039 109348 -24995
rect 109404 -25039 109448 -24995
rect 109504 -25039 109548 -24995
rect 109604 -25039 109648 -24995
rect 109704 -25039 109748 -24995
rect 109804 -25039 109848 -24995
rect 109904 -25039 109948 -24995
rect 110004 -25039 110048 -24995
rect 110104 -25039 110148 -24995
rect 110204 -25039 110248 -24995
rect 110304 -25039 110348 -24995
rect 110404 -25039 110448 -24995
rect 110504 -25039 110548 -24995
rect 110604 -25039 110648 -24995
rect 111104 -25039 111148 -24995
rect 111204 -25039 111248 -24995
rect 111304 -25039 111348 -24995
rect 111404 -25039 111448 -24995
rect 111504 -25039 111548 -24995
rect 111604 -25039 111648 -24995
rect 111704 -25039 111748 -24995
rect 111804 -25039 111848 -24995
rect 111904 -25039 111948 -24995
rect 112004 -25039 112048 -24995
rect 112104 -25039 112148 -24995
rect 112204 -25039 112248 -24995
rect 112304 -25039 112348 -24995
rect 112404 -25039 112448 -24995
rect 112504 -25039 112548 -24995
rect 112604 -25039 112648 -24995
rect 113104 -25039 113148 -24995
rect 113204 -25039 113248 -24995
rect 113304 -25039 113348 -24995
rect 113404 -25039 113448 -24995
rect 113504 -25039 113548 -24995
rect 113604 -25039 113648 -24995
rect 113704 -25039 113748 -24995
rect 113804 -25039 113848 -24995
rect 113904 -25039 113948 -24995
rect 114004 -25039 114048 -24995
rect 114104 -25039 114148 -24995
rect 114204 -25039 114248 -24995
rect 114304 -25039 114348 -24995
rect 114404 -25039 114448 -24995
rect 114504 -25039 114548 -24995
rect 114604 -25039 114648 -24995
rect 115104 -25039 115148 -24995
rect 115204 -25039 115248 -24995
rect 115304 -25039 115348 -24995
rect 115404 -25039 115448 -24995
rect 115504 -25039 115548 -24995
rect 115604 -25039 115648 -24995
rect 115704 -25039 115748 -24995
rect 115804 -25039 115848 -24995
rect 115904 -25039 115948 -24995
rect 116004 -25039 116048 -24995
rect 116104 -25039 116148 -24995
rect 116204 -25039 116248 -24995
rect 116304 -25039 116348 -24995
rect 116404 -25039 116448 -24995
rect 116504 -25039 116548 -24995
rect 116604 -25039 116648 -24995
rect -82799 -25210 -82755 -25166
rect -82699 -25210 -82655 -25166
rect -82599 -25210 -82555 -25166
rect -82499 -25210 -82455 -25166
rect -82399 -25210 -82355 -25166
rect -82299 -25210 -82255 -25166
rect -82199 -25210 -82155 -25166
rect -82099 -25210 -82055 -25166
rect -81999 -25210 -81955 -25166
rect -81899 -25210 -81855 -25166
rect -81799 -25210 -81755 -25166
rect -81699 -25210 -81655 -25166
rect -81599 -25210 -81555 -25166
rect -81499 -25210 -81455 -25166
rect -81399 -25210 -81355 -25166
rect -81299 -25210 -81255 -25166
rect -80799 -25210 -80755 -25166
rect -80699 -25210 -80655 -25166
rect -80599 -25210 -80555 -25166
rect -80499 -25210 -80455 -25166
rect -80399 -25210 -80355 -25166
rect -80299 -25210 -80255 -25166
rect -80199 -25210 -80155 -25166
rect -80099 -25210 -80055 -25166
rect -79999 -25210 -79955 -25166
rect -79899 -25210 -79855 -25166
rect -79799 -25210 -79755 -25166
rect -79699 -25210 -79655 -25166
rect -79599 -25210 -79555 -25166
rect -79499 -25210 -79455 -25166
rect -79399 -25210 -79355 -25166
rect -79299 -25210 -79255 -25166
rect -78799 -25210 -78755 -25166
rect -78699 -25210 -78655 -25166
rect -78599 -25210 -78555 -25166
rect -78499 -25210 -78455 -25166
rect -78399 -25210 -78355 -25166
rect -78299 -25210 -78255 -25166
rect -78199 -25210 -78155 -25166
rect -78099 -25210 -78055 -25166
rect -77999 -25210 -77955 -25166
rect -77899 -25210 -77855 -25166
rect -77799 -25210 -77755 -25166
rect -77699 -25210 -77655 -25166
rect -77599 -25210 -77555 -25166
rect -77499 -25210 -77455 -25166
rect -77399 -25210 -77355 -25166
rect -77299 -25210 -77255 -25166
rect -76799 -25210 -76755 -25166
rect -76699 -25210 -76655 -25166
rect -76599 -25210 -76555 -25166
rect -76499 -25210 -76455 -25166
rect -76399 -25210 -76355 -25166
rect -76299 -25210 -76255 -25166
rect -76199 -25210 -76155 -25166
rect -76099 -25210 -76055 -25166
rect -75999 -25210 -75955 -25166
rect -75899 -25210 -75855 -25166
rect -75799 -25210 -75755 -25166
rect -75699 -25210 -75655 -25166
rect -75599 -25210 -75555 -25166
rect -75499 -25210 -75455 -25166
rect -75399 -25210 -75355 -25166
rect -75299 -25210 -75255 -25166
rect 80849 -25170 80893 -25126
rect 80949 -25170 80993 -25126
rect 81049 -25170 81093 -25126
rect 81149 -25170 81193 -25126
rect 81249 -25170 81293 -25126
rect 81349 -25170 81393 -25126
rect 81449 -25170 81493 -25126
rect 81549 -25170 81593 -25126
rect 81649 -25170 81693 -25126
rect 81749 -25170 81793 -25126
rect 81849 -25170 81893 -25126
rect 81949 -25170 81993 -25126
rect 82049 -25170 82093 -25126
rect 82149 -25170 82193 -25126
rect 82249 -25170 82293 -25126
rect 82349 -25170 82393 -25126
rect 82849 -25170 82893 -25126
rect 82949 -25170 82993 -25126
rect 83049 -25170 83093 -25126
rect 83149 -25170 83193 -25126
rect 83249 -25170 83293 -25126
rect 83349 -25170 83393 -25126
rect 83449 -25170 83493 -25126
rect 83549 -25170 83593 -25126
rect 83649 -25170 83693 -25126
rect 83749 -25170 83793 -25126
rect 83849 -25170 83893 -25126
rect 83949 -25170 83993 -25126
rect 84049 -25170 84093 -25126
rect 84149 -25170 84193 -25126
rect 84249 -25170 84293 -25126
rect 84349 -25170 84393 -25126
rect 84849 -25170 84893 -25126
rect 84949 -25170 84993 -25126
rect 85049 -25170 85093 -25126
rect 85149 -25170 85193 -25126
rect 85249 -25170 85293 -25126
rect 85349 -25170 85393 -25126
rect 85449 -25170 85493 -25126
rect 85549 -25170 85593 -25126
rect 85649 -25170 85693 -25126
rect 85749 -25170 85793 -25126
rect 85849 -25170 85893 -25126
rect 85949 -25170 85993 -25126
rect 86049 -25170 86093 -25126
rect 86149 -25170 86193 -25126
rect 86249 -25170 86293 -25126
rect 86349 -25170 86393 -25126
rect 86849 -25170 86893 -25126
rect 86949 -25170 86993 -25126
rect 87049 -25170 87093 -25126
rect 87149 -25170 87193 -25126
rect 87249 -25170 87293 -25126
rect 87349 -25170 87393 -25126
rect 87449 -25170 87493 -25126
rect 87549 -25170 87593 -25126
rect 87649 -25170 87693 -25126
rect 87749 -25170 87793 -25126
rect 87849 -25170 87893 -25126
rect 87949 -25170 87993 -25126
rect 88049 -25170 88093 -25126
rect 88149 -25170 88193 -25126
rect 88249 -25170 88293 -25126
rect 88349 -25170 88393 -25126
rect 109104 -25139 109148 -25095
rect 109204 -25139 109248 -25095
rect 109304 -25139 109348 -25095
rect 109404 -25139 109448 -25095
rect 109504 -25139 109548 -25095
rect 109604 -25139 109648 -25095
rect 109704 -25139 109748 -25095
rect 109804 -25139 109848 -25095
rect 109904 -25139 109948 -25095
rect 110004 -25139 110048 -25095
rect 110104 -25139 110148 -25095
rect 110204 -25139 110248 -25095
rect 110304 -25139 110348 -25095
rect 110404 -25139 110448 -25095
rect 110504 -25139 110548 -25095
rect 110604 -25139 110648 -25095
rect 111104 -25139 111148 -25095
rect 111204 -25139 111248 -25095
rect 111304 -25139 111348 -25095
rect 111404 -25139 111448 -25095
rect 111504 -25139 111548 -25095
rect 111604 -25139 111648 -25095
rect 111704 -25139 111748 -25095
rect 111804 -25139 111848 -25095
rect 111904 -25139 111948 -25095
rect 112004 -25139 112048 -25095
rect 112104 -25139 112148 -25095
rect 112204 -25139 112248 -25095
rect 112304 -25139 112348 -25095
rect 112404 -25139 112448 -25095
rect 112504 -25139 112548 -25095
rect 112604 -25139 112648 -25095
rect 113104 -25139 113148 -25095
rect 113204 -25139 113248 -25095
rect 113304 -25139 113348 -25095
rect 113404 -25139 113448 -25095
rect 113504 -25139 113548 -25095
rect 113604 -25139 113648 -25095
rect 113704 -25139 113748 -25095
rect 113804 -25139 113848 -25095
rect 113904 -25139 113948 -25095
rect 114004 -25139 114048 -25095
rect 114104 -25139 114148 -25095
rect 114204 -25139 114248 -25095
rect 114304 -25139 114348 -25095
rect 114404 -25139 114448 -25095
rect 114504 -25139 114548 -25095
rect 114604 -25139 114648 -25095
rect 115104 -25139 115148 -25095
rect 115204 -25139 115248 -25095
rect 115304 -25139 115348 -25095
rect 115404 -25139 115448 -25095
rect 115504 -25139 115548 -25095
rect 115604 -25139 115648 -25095
rect 115704 -25139 115748 -25095
rect 115804 -25139 115848 -25095
rect 115904 -25139 115948 -25095
rect 116004 -25139 116048 -25095
rect 116104 -25139 116148 -25095
rect 116204 -25139 116248 -25095
rect 116304 -25139 116348 -25095
rect 116404 -25139 116448 -25095
rect 116504 -25139 116548 -25095
rect 116604 -25139 116648 -25095
rect -82799 -25310 -82755 -25266
rect -82699 -25310 -82655 -25266
rect -82599 -25310 -82555 -25266
rect -82499 -25310 -82455 -25266
rect -82399 -25310 -82355 -25266
rect -82299 -25310 -82255 -25266
rect -82199 -25310 -82155 -25266
rect -82099 -25310 -82055 -25266
rect -81999 -25310 -81955 -25266
rect -81899 -25310 -81855 -25266
rect -81799 -25310 -81755 -25266
rect -81699 -25310 -81655 -25266
rect -81599 -25310 -81555 -25266
rect -81499 -25310 -81455 -25266
rect -81399 -25310 -81355 -25266
rect -81299 -25310 -81255 -25266
rect -80799 -25310 -80755 -25266
rect -80699 -25310 -80655 -25266
rect -80599 -25310 -80555 -25266
rect -80499 -25310 -80455 -25266
rect -80399 -25310 -80355 -25266
rect -80299 -25310 -80255 -25266
rect -80199 -25310 -80155 -25266
rect -80099 -25310 -80055 -25266
rect -79999 -25310 -79955 -25266
rect -79899 -25310 -79855 -25266
rect -79799 -25310 -79755 -25266
rect -79699 -25310 -79655 -25266
rect -79599 -25310 -79555 -25266
rect -79499 -25310 -79455 -25266
rect -79399 -25310 -79355 -25266
rect -79299 -25310 -79255 -25266
rect -78799 -25310 -78755 -25266
rect -78699 -25310 -78655 -25266
rect -78599 -25310 -78555 -25266
rect -78499 -25310 -78455 -25266
rect -78399 -25310 -78355 -25266
rect -78299 -25310 -78255 -25266
rect -78199 -25310 -78155 -25266
rect -78099 -25310 -78055 -25266
rect -77999 -25310 -77955 -25266
rect -77899 -25310 -77855 -25266
rect -77799 -25310 -77755 -25266
rect -77699 -25310 -77655 -25266
rect -77599 -25310 -77555 -25266
rect -77499 -25310 -77455 -25266
rect -77399 -25310 -77355 -25266
rect -77299 -25310 -77255 -25266
rect -76799 -25310 -76755 -25266
rect -76699 -25310 -76655 -25266
rect -76599 -25310 -76555 -25266
rect -76499 -25310 -76455 -25266
rect -76399 -25310 -76355 -25266
rect -76299 -25310 -76255 -25266
rect -76199 -25310 -76155 -25266
rect -76099 -25310 -76055 -25266
rect -75999 -25310 -75955 -25266
rect -75899 -25310 -75855 -25266
rect -75799 -25310 -75755 -25266
rect -75699 -25310 -75655 -25266
rect -75599 -25310 -75555 -25266
rect -75499 -25310 -75455 -25266
rect -75399 -25310 -75355 -25266
rect -75299 -25310 -75255 -25266
rect 80849 -25270 80893 -25226
rect 80949 -25270 80993 -25226
rect 81049 -25270 81093 -25226
rect 81149 -25270 81193 -25226
rect 81249 -25270 81293 -25226
rect 81349 -25270 81393 -25226
rect 81449 -25270 81493 -25226
rect 81549 -25270 81593 -25226
rect 81649 -25270 81693 -25226
rect 81749 -25270 81793 -25226
rect 81849 -25270 81893 -25226
rect 81949 -25270 81993 -25226
rect 82049 -25270 82093 -25226
rect 82149 -25270 82193 -25226
rect 82249 -25270 82293 -25226
rect 82349 -25270 82393 -25226
rect 82849 -25270 82893 -25226
rect 82949 -25270 82993 -25226
rect 83049 -25270 83093 -25226
rect 83149 -25270 83193 -25226
rect 83249 -25270 83293 -25226
rect 83349 -25270 83393 -25226
rect 83449 -25270 83493 -25226
rect 83549 -25270 83593 -25226
rect 83649 -25270 83693 -25226
rect 83749 -25270 83793 -25226
rect 83849 -25270 83893 -25226
rect 83949 -25270 83993 -25226
rect 84049 -25270 84093 -25226
rect 84149 -25270 84193 -25226
rect 84249 -25270 84293 -25226
rect 84349 -25270 84393 -25226
rect 84849 -25270 84893 -25226
rect 84949 -25270 84993 -25226
rect 85049 -25270 85093 -25226
rect 85149 -25270 85193 -25226
rect 85249 -25270 85293 -25226
rect 85349 -25270 85393 -25226
rect 85449 -25270 85493 -25226
rect 85549 -25270 85593 -25226
rect 85649 -25270 85693 -25226
rect 85749 -25270 85793 -25226
rect 85849 -25270 85893 -25226
rect 85949 -25270 85993 -25226
rect 86049 -25270 86093 -25226
rect 86149 -25270 86193 -25226
rect 86249 -25270 86293 -25226
rect 86349 -25270 86393 -25226
rect 86849 -25270 86893 -25226
rect 86949 -25270 86993 -25226
rect 87049 -25270 87093 -25226
rect 87149 -25270 87193 -25226
rect 87249 -25270 87293 -25226
rect 87349 -25270 87393 -25226
rect 87449 -25270 87493 -25226
rect 87549 -25270 87593 -25226
rect 87649 -25270 87693 -25226
rect 87749 -25270 87793 -25226
rect 87849 -25270 87893 -25226
rect 87949 -25270 87993 -25226
rect 88049 -25270 88093 -25226
rect 88149 -25270 88193 -25226
rect 88249 -25270 88293 -25226
rect 88349 -25270 88393 -25226
rect 109104 -25239 109148 -25195
rect 109204 -25239 109248 -25195
rect 109304 -25239 109348 -25195
rect 109404 -25239 109448 -25195
rect 109504 -25239 109548 -25195
rect 109604 -25239 109648 -25195
rect 109704 -25239 109748 -25195
rect 109804 -25239 109848 -25195
rect 109904 -25239 109948 -25195
rect 110004 -25239 110048 -25195
rect 110104 -25239 110148 -25195
rect 110204 -25239 110248 -25195
rect 110304 -25239 110348 -25195
rect 110404 -25239 110448 -25195
rect 110504 -25239 110548 -25195
rect 110604 -25239 110648 -25195
rect 111104 -25239 111148 -25195
rect 111204 -25239 111248 -25195
rect 111304 -25239 111348 -25195
rect 111404 -25239 111448 -25195
rect 111504 -25239 111548 -25195
rect 111604 -25239 111648 -25195
rect 111704 -25239 111748 -25195
rect 111804 -25239 111848 -25195
rect 111904 -25239 111948 -25195
rect 112004 -25239 112048 -25195
rect 112104 -25239 112148 -25195
rect 112204 -25239 112248 -25195
rect 112304 -25239 112348 -25195
rect 112404 -25239 112448 -25195
rect 112504 -25239 112548 -25195
rect 112604 -25239 112648 -25195
rect 113104 -25239 113148 -25195
rect 113204 -25239 113248 -25195
rect 113304 -25239 113348 -25195
rect 113404 -25239 113448 -25195
rect 113504 -25239 113548 -25195
rect 113604 -25239 113648 -25195
rect 113704 -25239 113748 -25195
rect 113804 -25239 113848 -25195
rect 113904 -25239 113948 -25195
rect 114004 -25239 114048 -25195
rect 114104 -25239 114148 -25195
rect 114204 -25239 114248 -25195
rect 114304 -25239 114348 -25195
rect 114404 -25239 114448 -25195
rect 114504 -25239 114548 -25195
rect 114604 -25239 114648 -25195
rect 115104 -25239 115148 -25195
rect 115204 -25239 115248 -25195
rect 115304 -25239 115348 -25195
rect 115404 -25239 115448 -25195
rect 115504 -25239 115548 -25195
rect 115604 -25239 115648 -25195
rect 115704 -25239 115748 -25195
rect 115804 -25239 115848 -25195
rect 115904 -25239 115948 -25195
rect 116004 -25239 116048 -25195
rect 116104 -25239 116148 -25195
rect 116204 -25239 116248 -25195
rect 116304 -25239 116348 -25195
rect 116404 -25239 116448 -25195
rect 116504 -25239 116548 -25195
rect 116604 -25239 116648 -25195
rect -82799 -25410 -82755 -25366
rect -82699 -25410 -82655 -25366
rect -82599 -25410 -82555 -25366
rect -82499 -25410 -82455 -25366
rect -82399 -25410 -82355 -25366
rect -82299 -25410 -82255 -25366
rect -82199 -25410 -82155 -25366
rect -82099 -25410 -82055 -25366
rect -81999 -25410 -81955 -25366
rect -81899 -25410 -81855 -25366
rect -81799 -25410 -81755 -25366
rect -81699 -25410 -81655 -25366
rect -81599 -25410 -81555 -25366
rect -81499 -25410 -81455 -25366
rect -81399 -25410 -81355 -25366
rect -81299 -25410 -81255 -25366
rect -80799 -25410 -80755 -25366
rect -80699 -25410 -80655 -25366
rect -80599 -25410 -80555 -25366
rect -80499 -25410 -80455 -25366
rect -80399 -25410 -80355 -25366
rect -80299 -25410 -80255 -25366
rect -80199 -25410 -80155 -25366
rect -80099 -25410 -80055 -25366
rect -79999 -25410 -79955 -25366
rect -79899 -25410 -79855 -25366
rect -79799 -25410 -79755 -25366
rect -79699 -25410 -79655 -25366
rect -79599 -25410 -79555 -25366
rect -79499 -25410 -79455 -25366
rect -79399 -25410 -79355 -25366
rect -79299 -25410 -79255 -25366
rect -78799 -25410 -78755 -25366
rect -78699 -25410 -78655 -25366
rect -78599 -25410 -78555 -25366
rect -78499 -25410 -78455 -25366
rect -78399 -25410 -78355 -25366
rect -78299 -25410 -78255 -25366
rect -78199 -25410 -78155 -25366
rect -78099 -25410 -78055 -25366
rect -77999 -25410 -77955 -25366
rect -77899 -25410 -77855 -25366
rect -77799 -25410 -77755 -25366
rect -77699 -25410 -77655 -25366
rect -77599 -25410 -77555 -25366
rect -77499 -25410 -77455 -25366
rect -77399 -25410 -77355 -25366
rect -77299 -25410 -77255 -25366
rect -76799 -25410 -76755 -25366
rect -76699 -25410 -76655 -25366
rect -76599 -25410 -76555 -25366
rect -76499 -25410 -76455 -25366
rect -76399 -25410 -76355 -25366
rect -76299 -25410 -76255 -25366
rect -76199 -25410 -76155 -25366
rect -76099 -25410 -76055 -25366
rect -75999 -25410 -75955 -25366
rect -75899 -25410 -75855 -25366
rect -75799 -25410 -75755 -25366
rect -75699 -25410 -75655 -25366
rect -75599 -25410 -75555 -25366
rect -75499 -25410 -75455 -25366
rect -75399 -25410 -75355 -25366
rect -75299 -25410 -75255 -25366
rect 80849 -25370 80893 -25326
rect 80949 -25370 80993 -25326
rect 81049 -25370 81093 -25326
rect 81149 -25370 81193 -25326
rect 81249 -25370 81293 -25326
rect 81349 -25370 81393 -25326
rect 81449 -25370 81493 -25326
rect 81549 -25370 81593 -25326
rect 81649 -25370 81693 -25326
rect 81749 -25370 81793 -25326
rect 81849 -25370 81893 -25326
rect 81949 -25370 81993 -25326
rect 82049 -25370 82093 -25326
rect 82149 -25370 82193 -25326
rect 82249 -25370 82293 -25326
rect 82349 -25370 82393 -25326
rect 82849 -25370 82893 -25326
rect 82949 -25370 82993 -25326
rect 83049 -25370 83093 -25326
rect 83149 -25370 83193 -25326
rect 83249 -25370 83293 -25326
rect 83349 -25370 83393 -25326
rect 83449 -25370 83493 -25326
rect 83549 -25370 83593 -25326
rect 83649 -25370 83693 -25326
rect 83749 -25370 83793 -25326
rect 83849 -25370 83893 -25326
rect 83949 -25370 83993 -25326
rect 84049 -25370 84093 -25326
rect 84149 -25370 84193 -25326
rect 84249 -25370 84293 -25326
rect 84349 -25370 84393 -25326
rect 84849 -25370 84893 -25326
rect 84949 -25370 84993 -25326
rect 85049 -25370 85093 -25326
rect 85149 -25370 85193 -25326
rect 85249 -25370 85293 -25326
rect 85349 -25370 85393 -25326
rect 85449 -25370 85493 -25326
rect 85549 -25370 85593 -25326
rect 85649 -25370 85693 -25326
rect 85749 -25370 85793 -25326
rect 85849 -25370 85893 -25326
rect 85949 -25370 85993 -25326
rect 86049 -25370 86093 -25326
rect 86149 -25370 86193 -25326
rect 86249 -25370 86293 -25326
rect 86349 -25370 86393 -25326
rect 86849 -25370 86893 -25326
rect 86949 -25370 86993 -25326
rect 87049 -25370 87093 -25326
rect 87149 -25370 87193 -25326
rect 87249 -25370 87293 -25326
rect 87349 -25370 87393 -25326
rect 87449 -25370 87493 -25326
rect 87549 -25370 87593 -25326
rect 87649 -25370 87693 -25326
rect 87749 -25370 87793 -25326
rect 87849 -25370 87893 -25326
rect 87949 -25370 87993 -25326
rect 88049 -25370 88093 -25326
rect 88149 -25370 88193 -25326
rect 88249 -25370 88293 -25326
rect 88349 -25370 88393 -25326
rect 109104 -25339 109148 -25295
rect 109204 -25339 109248 -25295
rect 109304 -25339 109348 -25295
rect 109404 -25339 109448 -25295
rect 109504 -25339 109548 -25295
rect 109604 -25339 109648 -25295
rect 109704 -25339 109748 -25295
rect 109804 -25339 109848 -25295
rect 109904 -25339 109948 -25295
rect 110004 -25339 110048 -25295
rect 110104 -25339 110148 -25295
rect 110204 -25339 110248 -25295
rect 110304 -25339 110348 -25295
rect 110404 -25339 110448 -25295
rect 110504 -25339 110548 -25295
rect 110604 -25339 110648 -25295
rect 111104 -25339 111148 -25295
rect 111204 -25339 111248 -25295
rect 111304 -25339 111348 -25295
rect 111404 -25339 111448 -25295
rect 111504 -25339 111548 -25295
rect 111604 -25339 111648 -25295
rect 111704 -25339 111748 -25295
rect 111804 -25339 111848 -25295
rect 111904 -25339 111948 -25295
rect 112004 -25339 112048 -25295
rect 112104 -25339 112148 -25295
rect 112204 -25339 112248 -25295
rect 112304 -25339 112348 -25295
rect 112404 -25339 112448 -25295
rect 112504 -25339 112548 -25295
rect 112604 -25339 112648 -25295
rect 113104 -25339 113148 -25295
rect 113204 -25339 113248 -25295
rect 113304 -25339 113348 -25295
rect 113404 -25339 113448 -25295
rect 113504 -25339 113548 -25295
rect 113604 -25339 113648 -25295
rect 113704 -25339 113748 -25295
rect 113804 -25339 113848 -25295
rect 113904 -25339 113948 -25295
rect 114004 -25339 114048 -25295
rect 114104 -25339 114148 -25295
rect 114204 -25339 114248 -25295
rect 114304 -25339 114348 -25295
rect 114404 -25339 114448 -25295
rect 114504 -25339 114548 -25295
rect 114604 -25339 114648 -25295
rect 115104 -25339 115148 -25295
rect 115204 -25339 115248 -25295
rect 115304 -25339 115348 -25295
rect 115404 -25339 115448 -25295
rect 115504 -25339 115548 -25295
rect 115604 -25339 115648 -25295
rect 115704 -25339 115748 -25295
rect 115804 -25339 115848 -25295
rect 115904 -25339 115948 -25295
rect 116004 -25339 116048 -25295
rect 116104 -25339 116148 -25295
rect 116204 -25339 116248 -25295
rect 116304 -25339 116348 -25295
rect 116404 -25339 116448 -25295
rect 116504 -25339 116548 -25295
rect 116604 -25339 116648 -25295
rect -82799 -25510 -82755 -25466
rect -82699 -25510 -82655 -25466
rect -82599 -25510 -82555 -25466
rect -82499 -25510 -82455 -25466
rect -82399 -25510 -82355 -25466
rect -82299 -25510 -82255 -25466
rect -82199 -25510 -82155 -25466
rect -82099 -25510 -82055 -25466
rect -81999 -25510 -81955 -25466
rect -81899 -25510 -81855 -25466
rect -81799 -25510 -81755 -25466
rect -81699 -25510 -81655 -25466
rect -81599 -25510 -81555 -25466
rect -81499 -25510 -81455 -25466
rect -81399 -25510 -81355 -25466
rect -81299 -25510 -81255 -25466
rect -80799 -25510 -80755 -25466
rect -80699 -25510 -80655 -25466
rect -80599 -25510 -80555 -25466
rect -80499 -25510 -80455 -25466
rect -80399 -25510 -80355 -25466
rect -80299 -25510 -80255 -25466
rect -80199 -25510 -80155 -25466
rect -80099 -25510 -80055 -25466
rect -79999 -25510 -79955 -25466
rect -79899 -25510 -79855 -25466
rect -79799 -25510 -79755 -25466
rect -79699 -25510 -79655 -25466
rect -79599 -25510 -79555 -25466
rect -79499 -25510 -79455 -25466
rect -79399 -25510 -79355 -25466
rect -79299 -25510 -79255 -25466
rect -78799 -25510 -78755 -25466
rect -78699 -25510 -78655 -25466
rect -78599 -25510 -78555 -25466
rect -78499 -25510 -78455 -25466
rect -78399 -25510 -78355 -25466
rect -78299 -25510 -78255 -25466
rect -78199 -25510 -78155 -25466
rect -78099 -25510 -78055 -25466
rect -77999 -25510 -77955 -25466
rect -77899 -25510 -77855 -25466
rect -77799 -25510 -77755 -25466
rect -77699 -25510 -77655 -25466
rect -77599 -25510 -77555 -25466
rect -77499 -25510 -77455 -25466
rect -77399 -25510 -77355 -25466
rect -77299 -25510 -77255 -25466
rect -76799 -25510 -76755 -25466
rect -76699 -25510 -76655 -25466
rect -76599 -25510 -76555 -25466
rect -76499 -25510 -76455 -25466
rect -76399 -25510 -76355 -25466
rect -76299 -25510 -76255 -25466
rect -76199 -25510 -76155 -25466
rect -76099 -25510 -76055 -25466
rect -75999 -25510 -75955 -25466
rect -75899 -25510 -75855 -25466
rect -75799 -25510 -75755 -25466
rect -75699 -25510 -75655 -25466
rect -75599 -25510 -75555 -25466
rect -75499 -25510 -75455 -25466
rect -75399 -25510 -75355 -25466
rect -75299 -25510 -75255 -25466
rect 80849 -25470 80893 -25426
rect 80949 -25470 80993 -25426
rect 81049 -25470 81093 -25426
rect 81149 -25470 81193 -25426
rect 81249 -25470 81293 -25426
rect 81349 -25470 81393 -25426
rect 81449 -25470 81493 -25426
rect 81549 -25470 81593 -25426
rect 81649 -25470 81693 -25426
rect 81749 -25470 81793 -25426
rect 81849 -25470 81893 -25426
rect 81949 -25470 81993 -25426
rect 82049 -25470 82093 -25426
rect 82149 -25470 82193 -25426
rect 82249 -25470 82293 -25426
rect 82349 -25470 82393 -25426
rect 82849 -25470 82893 -25426
rect 82949 -25470 82993 -25426
rect 83049 -25470 83093 -25426
rect 83149 -25470 83193 -25426
rect 83249 -25470 83293 -25426
rect 83349 -25470 83393 -25426
rect 83449 -25470 83493 -25426
rect 83549 -25470 83593 -25426
rect 83649 -25470 83693 -25426
rect 83749 -25470 83793 -25426
rect 83849 -25470 83893 -25426
rect 83949 -25470 83993 -25426
rect 84049 -25470 84093 -25426
rect 84149 -25470 84193 -25426
rect 84249 -25470 84293 -25426
rect 84349 -25470 84393 -25426
rect 84849 -25470 84893 -25426
rect 84949 -25470 84993 -25426
rect 85049 -25470 85093 -25426
rect 85149 -25470 85193 -25426
rect 85249 -25470 85293 -25426
rect 85349 -25470 85393 -25426
rect 85449 -25470 85493 -25426
rect 85549 -25470 85593 -25426
rect 85649 -25470 85693 -25426
rect 85749 -25470 85793 -25426
rect 85849 -25470 85893 -25426
rect 85949 -25470 85993 -25426
rect 86049 -25470 86093 -25426
rect 86149 -25470 86193 -25426
rect 86249 -25470 86293 -25426
rect 86349 -25470 86393 -25426
rect 86849 -25470 86893 -25426
rect 86949 -25470 86993 -25426
rect 87049 -25470 87093 -25426
rect 87149 -25470 87193 -25426
rect 87249 -25470 87293 -25426
rect 87349 -25470 87393 -25426
rect 87449 -25470 87493 -25426
rect 87549 -25470 87593 -25426
rect 87649 -25470 87693 -25426
rect 87749 -25470 87793 -25426
rect 87849 -25470 87893 -25426
rect 87949 -25470 87993 -25426
rect 88049 -25470 88093 -25426
rect 88149 -25470 88193 -25426
rect 88249 -25470 88293 -25426
rect 88349 -25470 88393 -25426
rect 109104 -25439 109148 -25395
rect 109204 -25439 109248 -25395
rect 109304 -25439 109348 -25395
rect 109404 -25439 109448 -25395
rect 109504 -25439 109548 -25395
rect 109604 -25439 109648 -25395
rect 109704 -25439 109748 -25395
rect 109804 -25439 109848 -25395
rect 109904 -25439 109948 -25395
rect 110004 -25439 110048 -25395
rect 110104 -25439 110148 -25395
rect 110204 -25439 110248 -25395
rect 110304 -25439 110348 -25395
rect 110404 -25439 110448 -25395
rect 110504 -25439 110548 -25395
rect 110604 -25439 110648 -25395
rect 111104 -25439 111148 -25395
rect 111204 -25439 111248 -25395
rect 111304 -25439 111348 -25395
rect 111404 -25439 111448 -25395
rect 111504 -25439 111548 -25395
rect 111604 -25439 111648 -25395
rect 111704 -25439 111748 -25395
rect 111804 -25439 111848 -25395
rect 111904 -25439 111948 -25395
rect 112004 -25439 112048 -25395
rect 112104 -25439 112148 -25395
rect 112204 -25439 112248 -25395
rect 112304 -25439 112348 -25395
rect 112404 -25439 112448 -25395
rect 112504 -25439 112548 -25395
rect 112604 -25439 112648 -25395
rect 113104 -25439 113148 -25395
rect 113204 -25439 113248 -25395
rect 113304 -25439 113348 -25395
rect 113404 -25439 113448 -25395
rect 113504 -25439 113548 -25395
rect 113604 -25439 113648 -25395
rect 113704 -25439 113748 -25395
rect 113804 -25439 113848 -25395
rect 113904 -25439 113948 -25395
rect 114004 -25439 114048 -25395
rect 114104 -25439 114148 -25395
rect 114204 -25439 114248 -25395
rect 114304 -25439 114348 -25395
rect 114404 -25439 114448 -25395
rect 114504 -25439 114548 -25395
rect 114604 -25439 114648 -25395
rect 115104 -25439 115148 -25395
rect 115204 -25439 115248 -25395
rect 115304 -25439 115348 -25395
rect 115404 -25439 115448 -25395
rect 115504 -25439 115548 -25395
rect 115604 -25439 115648 -25395
rect 115704 -25439 115748 -25395
rect 115804 -25439 115848 -25395
rect 115904 -25439 115948 -25395
rect 116004 -25439 116048 -25395
rect 116104 -25439 116148 -25395
rect 116204 -25439 116248 -25395
rect 116304 -25439 116348 -25395
rect 116404 -25439 116448 -25395
rect 116504 -25439 116548 -25395
rect 116604 -25439 116648 -25395
rect -82799 -25610 -82755 -25566
rect -82699 -25610 -82655 -25566
rect -82599 -25610 -82555 -25566
rect -82499 -25610 -82455 -25566
rect -82399 -25610 -82355 -25566
rect -82299 -25610 -82255 -25566
rect -82199 -25610 -82155 -25566
rect -82099 -25610 -82055 -25566
rect -81999 -25610 -81955 -25566
rect -81899 -25610 -81855 -25566
rect -81799 -25610 -81755 -25566
rect -81699 -25610 -81655 -25566
rect -81599 -25610 -81555 -25566
rect -81499 -25610 -81455 -25566
rect -81399 -25610 -81355 -25566
rect -81299 -25610 -81255 -25566
rect -80799 -25610 -80755 -25566
rect -80699 -25610 -80655 -25566
rect -80599 -25610 -80555 -25566
rect -80499 -25610 -80455 -25566
rect -80399 -25610 -80355 -25566
rect -80299 -25610 -80255 -25566
rect -80199 -25610 -80155 -25566
rect -80099 -25610 -80055 -25566
rect -79999 -25610 -79955 -25566
rect -79899 -25610 -79855 -25566
rect -79799 -25610 -79755 -25566
rect -79699 -25610 -79655 -25566
rect -79599 -25610 -79555 -25566
rect -79499 -25610 -79455 -25566
rect -79399 -25610 -79355 -25566
rect -79299 -25610 -79255 -25566
rect -78799 -25610 -78755 -25566
rect -78699 -25610 -78655 -25566
rect -78599 -25610 -78555 -25566
rect -78499 -25610 -78455 -25566
rect -78399 -25610 -78355 -25566
rect -78299 -25610 -78255 -25566
rect -78199 -25610 -78155 -25566
rect -78099 -25610 -78055 -25566
rect -77999 -25610 -77955 -25566
rect -77899 -25610 -77855 -25566
rect -77799 -25610 -77755 -25566
rect -77699 -25610 -77655 -25566
rect -77599 -25610 -77555 -25566
rect -77499 -25610 -77455 -25566
rect -77399 -25610 -77355 -25566
rect -77299 -25610 -77255 -25566
rect -76799 -25610 -76755 -25566
rect -76699 -25610 -76655 -25566
rect -76599 -25610 -76555 -25566
rect -76499 -25610 -76455 -25566
rect -76399 -25610 -76355 -25566
rect -76299 -25610 -76255 -25566
rect -76199 -25610 -76155 -25566
rect -76099 -25610 -76055 -25566
rect -75999 -25610 -75955 -25566
rect -75899 -25610 -75855 -25566
rect -75799 -25610 -75755 -25566
rect -75699 -25610 -75655 -25566
rect -75599 -25610 -75555 -25566
rect -75499 -25610 -75455 -25566
rect -75399 -25610 -75355 -25566
rect -75299 -25610 -75255 -25566
rect 80849 -25570 80893 -25526
rect 80949 -25570 80993 -25526
rect 81049 -25570 81093 -25526
rect 81149 -25570 81193 -25526
rect 81249 -25570 81293 -25526
rect 81349 -25570 81393 -25526
rect 81449 -25570 81493 -25526
rect 81549 -25570 81593 -25526
rect 81649 -25570 81693 -25526
rect 81749 -25570 81793 -25526
rect 81849 -25570 81893 -25526
rect 81949 -25570 81993 -25526
rect 82049 -25570 82093 -25526
rect 82149 -25570 82193 -25526
rect 82249 -25570 82293 -25526
rect 82349 -25570 82393 -25526
rect 82849 -25570 82893 -25526
rect 82949 -25570 82993 -25526
rect 83049 -25570 83093 -25526
rect 83149 -25570 83193 -25526
rect 83249 -25570 83293 -25526
rect 83349 -25570 83393 -25526
rect 83449 -25570 83493 -25526
rect 83549 -25570 83593 -25526
rect 83649 -25570 83693 -25526
rect 83749 -25570 83793 -25526
rect 83849 -25570 83893 -25526
rect 83949 -25570 83993 -25526
rect 84049 -25570 84093 -25526
rect 84149 -25570 84193 -25526
rect 84249 -25570 84293 -25526
rect 84349 -25570 84393 -25526
rect 84849 -25570 84893 -25526
rect 84949 -25570 84993 -25526
rect 85049 -25570 85093 -25526
rect 85149 -25570 85193 -25526
rect 85249 -25570 85293 -25526
rect 85349 -25570 85393 -25526
rect 85449 -25570 85493 -25526
rect 85549 -25570 85593 -25526
rect 85649 -25570 85693 -25526
rect 85749 -25570 85793 -25526
rect 85849 -25570 85893 -25526
rect 85949 -25570 85993 -25526
rect 86049 -25570 86093 -25526
rect 86149 -25570 86193 -25526
rect 86249 -25570 86293 -25526
rect 86349 -25570 86393 -25526
rect 86849 -25570 86893 -25526
rect 86949 -25570 86993 -25526
rect 87049 -25570 87093 -25526
rect 87149 -25570 87193 -25526
rect 87249 -25570 87293 -25526
rect 87349 -25570 87393 -25526
rect 87449 -25570 87493 -25526
rect 87549 -25570 87593 -25526
rect 87649 -25570 87693 -25526
rect 87749 -25570 87793 -25526
rect 87849 -25570 87893 -25526
rect 87949 -25570 87993 -25526
rect 88049 -25570 88093 -25526
rect 88149 -25570 88193 -25526
rect 88249 -25570 88293 -25526
rect 88349 -25570 88393 -25526
rect 109104 -25539 109148 -25495
rect 109204 -25539 109248 -25495
rect 109304 -25539 109348 -25495
rect 109404 -25539 109448 -25495
rect 109504 -25539 109548 -25495
rect 109604 -25539 109648 -25495
rect 109704 -25539 109748 -25495
rect 109804 -25539 109848 -25495
rect 109904 -25539 109948 -25495
rect 110004 -25539 110048 -25495
rect 110104 -25539 110148 -25495
rect 110204 -25539 110248 -25495
rect 110304 -25539 110348 -25495
rect 110404 -25539 110448 -25495
rect 110504 -25539 110548 -25495
rect 110604 -25539 110648 -25495
rect 111104 -25539 111148 -25495
rect 111204 -25539 111248 -25495
rect 111304 -25539 111348 -25495
rect 111404 -25539 111448 -25495
rect 111504 -25539 111548 -25495
rect 111604 -25539 111648 -25495
rect 111704 -25539 111748 -25495
rect 111804 -25539 111848 -25495
rect 111904 -25539 111948 -25495
rect 112004 -25539 112048 -25495
rect 112104 -25539 112148 -25495
rect 112204 -25539 112248 -25495
rect 112304 -25539 112348 -25495
rect 112404 -25539 112448 -25495
rect 112504 -25539 112548 -25495
rect 112604 -25539 112648 -25495
rect 113104 -25539 113148 -25495
rect 113204 -25539 113248 -25495
rect 113304 -25539 113348 -25495
rect 113404 -25539 113448 -25495
rect 113504 -25539 113548 -25495
rect 113604 -25539 113648 -25495
rect 113704 -25539 113748 -25495
rect 113804 -25539 113848 -25495
rect 113904 -25539 113948 -25495
rect 114004 -25539 114048 -25495
rect 114104 -25539 114148 -25495
rect 114204 -25539 114248 -25495
rect 114304 -25539 114348 -25495
rect 114404 -25539 114448 -25495
rect 114504 -25539 114548 -25495
rect 114604 -25539 114648 -25495
rect 115104 -25539 115148 -25495
rect 115204 -25539 115248 -25495
rect 115304 -25539 115348 -25495
rect 115404 -25539 115448 -25495
rect 115504 -25539 115548 -25495
rect 115604 -25539 115648 -25495
rect 115704 -25539 115748 -25495
rect 115804 -25539 115848 -25495
rect 115904 -25539 115948 -25495
rect 116004 -25539 116048 -25495
rect 116104 -25539 116148 -25495
rect 116204 -25539 116248 -25495
rect 116304 -25539 116348 -25495
rect 116404 -25539 116448 -25495
rect 116504 -25539 116548 -25495
rect 116604 -25539 116648 -25495
rect 109104 -25639 109148 -25595
rect 109204 -25639 109248 -25595
rect 109304 -25639 109348 -25595
rect 109404 -25639 109448 -25595
rect 109504 -25639 109548 -25595
rect 109604 -25639 109648 -25595
rect 109704 -25639 109748 -25595
rect 109804 -25639 109848 -25595
rect 109904 -25639 109948 -25595
rect 110004 -25639 110048 -25595
rect 110104 -25639 110148 -25595
rect 110204 -25639 110248 -25595
rect 110304 -25639 110348 -25595
rect 110404 -25639 110448 -25595
rect 110504 -25639 110548 -25595
rect 110604 -25639 110648 -25595
rect 111104 -25639 111148 -25595
rect 111204 -25639 111248 -25595
rect 111304 -25639 111348 -25595
rect 111404 -25639 111448 -25595
rect 111504 -25639 111548 -25595
rect 111604 -25639 111648 -25595
rect 111704 -25639 111748 -25595
rect 111804 -25639 111848 -25595
rect 111904 -25639 111948 -25595
rect 112004 -25639 112048 -25595
rect 112104 -25639 112148 -25595
rect 112204 -25639 112248 -25595
rect 112304 -25639 112348 -25595
rect 112404 -25639 112448 -25595
rect 112504 -25639 112548 -25595
rect 112604 -25639 112648 -25595
rect 113104 -25639 113148 -25595
rect 113204 -25639 113248 -25595
rect 113304 -25639 113348 -25595
rect 113404 -25639 113448 -25595
rect 113504 -25639 113548 -25595
rect 113604 -25639 113648 -25595
rect 113704 -25639 113748 -25595
rect 113804 -25639 113848 -25595
rect 113904 -25639 113948 -25595
rect 114004 -25639 114048 -25595
rect 114104 -25639 114148 -25595
rect 114204 -25639 114248 -25595
rect 114304 -25639 114348 -25595
rect 114404 -25639 114448 -25595
rect 114504 -25639 114548 -25595
rect 114604 -25639 114648 -25595
rect 115104 -25639 115148 -25595
rect 115204 -25639 115248 -25595
rect 115304 -25639 115348 -25595
rect 115404 -25639 115448 -25595
rect 115504 -25639 115548 -25595
rect 115604 -25639 115648 -25595
rect 115704 -25639 115748 -25595
rect 115804 -25639 115848 -25595
rect 115904 -25639 115948 -25595
rect 116004 -25639 116048 -25595
rect 116104 -25639 116148 -25595
rect 116204 -25639 116248 -25595
rect 116304 -25639 116348 -25595
rect 116404 -25639 116448 -25595
rect 116504 -25639 116548 -25595
rect 116604 -25639 116648 -25595
rect -82799 -25710 -82755 -25666
rect -82699 -25710 -82655 -25666
rect -82599 -25710 -82555 -25666
rect -82499 -25710 -82455 -25666
rect -82399 -25710 -82355 -25666
rect -82299 -25710 -82255 -25666
rect -82199 -25710 -82155 -25666
rect -82099 -25710 -82055 -25666
rect -81999 -25710 -81955 -25666
rect -81899 -25710 -81855 -25666
rect -81799 -25710 -81755 -25666
rect -81699 -25710 -81655 -25666
rect -81599 -25710 -81555 -25666
rect -81499 -25710 -81455 -25666
rect -81399 -25710 -81355 -25666
rect -81299 -25710 -81255 -25666
rect -80799 -25710 -80755 -25666
rect -80699 -25710 -80655 -25666
rect -80599 -25710 -80555 -25666
rect -80499 -25710 -80455 -25666
rect -80399 -25710 -80355 -25666
rect -80299 -25710 -80255 -25666
rect -80199 -25710 -80155 -25666
rect -80099 -25710 -80055 -25666
rect -79999 -25710 -79955 -25666
rect -79899 -25710 -79855 -25666
rect -79799 -25710 -79755 -25666
rect -79699 -25710 -79655 -25666
rect -79599 -25710 -79555 -25666
rect -79499 -25710 -79455 -25666
rect -79399 -25710 -79355 -25666
rect -79299 -25710 -79255 -25666
rect -78799 -25710 -78755 -25666
rect -78699 -25710 -78655 -25666
rect -78599 -25710 -78555 -25666
rect -78499 -25710 -78455 -25666
rect -78399 -25710 -78355 -25666
rect -78299 -25710 -78255 -25666
rect -78199 -25710 -78155 -25666
rect -78099 -25710 -78055 -25666
rect -77999 -25710 -77955 -25666
rect -77899 -25710 -77855 -25666
rect -77799 -25710 -77755 -25666
rect -77699 -25710 -77655 -25666
rect -77599 -25710 -77555 -25666
rect -77499 -25710 -77455 -25666
rect -77399 -25710 -77355 -25666
rect -77299 -25710 -77255 -25666
rect -76799 -25710 -76755 -25666
rect -76699 -25710 -76655 -25666
rect -76599 -25710 -76555 -25666
rect -76499 -25710 -76455 -25666
rect -76399 -25710 -76355 -25666
rect -76299 -25710 -76255 -25666
rect -76199 -25710 -76155 -25666
rect -76099 -25710 -76055 -25666
rect -75999 -25710 -75955 -25666
rect -75899 -25710 -75855 -25666
rect -75799 -25710 -75755 -25666
rect -75699 -25710 -75655 -25666
rect -75599 -25710 -75555 -25666
rect -75499 -25710 -75455 -25666
rect -75399 -25710 -75355 -25666
rect -75299 -25710 -75255 -25666
rect 109104 -25739 109148 -25695
rect 109204 -25739 109248 -25695
rect 109304 -25739 109348 -25695
rect 109404 -25739 109448 -25695
rect 109504 -25739 109548 -25695
rect 109604 -25739 109648 -25695
rect 109704 -25739 109748 -25695
rect 109804 -25739 109848 -25695
rect 109904 -25739 109948 -25695
rect 110004 -25739 110048 -25695
rect 110104 -25739 110148 -25695
rect 110204 -25739 110248 -25695
rect 110304 -25739 110348 -25695
rect 110404 -25739 110448 -25695
rect 110504 -25739 110548 -25695
rect 110604 -25739 110648 -25695
rect 111104 -25739 111148 -25695
rect 111204 -25739 111248 -25695
rect 111304 -25739 111348 -25695
rect 111404 -25739 111448 -25695
rect 111504 -25739 111548 -25695
rect 111604 -25739 111648 -25695
rect 111704 -25739 111748 -25695
rect 111804 -25739 111848 -25695
rect 111904 -25739 111948 -25695
rect 112004 -25739 112048 -25695
rect 112104 -25739 112148 -25695
rect 112204 -25739 112248 -25695
rect 112304 -25739 112348 -25695
rect 112404 -25739 112448 -25695
rect 112504 -25739 112548 -25695
rect 112604 -25739 112648 -25695
rect 113104 -25739 113148 -25695
rect 113204 -25739 113248 -25695
rect 113304 -25739 113348 -25695
rect 113404 -25739 113448 -25695
rect 113504 -25739 113548 -25695
rect 113604 -25739 113648 -25695
rect 113704 -25739 113748 -25695
rect 113804 -25739 113848 -25695
rect 113904 -25739 113948 -25695
rect 114004 -25739 114048 -25695
rect 114104 -25739 114148 -25695
rect 114204 -25739 114248 -25695
rect 114304 -25739 114348 -25695
rect 114404 -25739 114448 -25695
rect 114504 -25739 114548 -25695
rect 114604 -25739 114648 -25695
rect 115104 -25739 115148 -25695
rect 115204 -25739 115248 -25695
rect 115304 -25739 115348 -25695
rect 115404 -25739 115448 -25695
rect 115504 -25739 115548 -25695
rect 115604 -25739 115648 -25695
rect 115704 -25739 115748 -25695
rect 115804 -25739 115848 -25695
rect 115904 -25739 115948 -25695
rect 116004 -25739 116048 -25695
rect 116104 -25739 116148 -25695
rect 116204 -25739 116248 -25695
rect 116304 -25739 116348 -25695
rect 116404 -25739 116448 -25695
rect 116504 -25739 116548 -25695
rect 116604 -25739 116648 -25695
rect -82799 -25810 -82755 -25766
rect -82699 -25810 -82655 -25766
rect -82599 -25810 -82555 -25766
rect -82499 -25810 -82455 -25766
rect -82399 -25810 -82355 -25766
rect -82299 -25810 -82255 -25766
rect -82199 -25810 -82155 -25766
rect -82099 -25810 -82055 -25766
rect -81999 -25810 -81955 -25766
rect -81899 -25810 -81855 -25766
rect -81799 -25810 -81755 -25766
rect -81699 -25810 -81655 -25766
rect -81599 -25810 -81555 -25766
rect -81499 -25810 -81455 -25766
rect -81399 -25810 -81355 -25766
rect -81299 -25810 -81255 -25766
rect -80799 -25810 -80755 -25766
rect -80699 -25810 -80655 -25766
rect -80599 -25810 -80555 -25766
rect -80499 -25810 -80455 -25766
rect -80399 -25810 -80355 -25766
rect -80299 -25810 -80255 -25766
rect -80199 -25810 -80155 -25766
rect -80099 -25810 -80055 -25766
rect -79999 -25810 -79955 -25766
rect -79899 -25810 -79855 -25766
rect -79799 -25810 -79755 -25766
rect -79699 -25810 -79655 -25766
rect -79599 -25810 -79555 -25766
rect -79499 -25810 -79455 -25766
rect -79399 -25810 -79355 -25766
rect -79299 -25810 -79255 -25766
rect -78799 -25810 -78755 -25766
rect -78699 -25810 -78655 -25766
rect -78599 -25810 -78555 -25766
rect -78499 -25810 -78455 -25766
rect -78399 -25810 -78355 -25766
rect -78299 -25810 -78255 -25766
rect -78199 -25810 -78155 -25766
rect -78099 -25810 -78055 -25766
rect -77999 -25810 -77955 -25766
rect -77899 -25810 -77855 -25766
rect -77799 -25810 -77755 -25766
rect -77699 -25810 -77655 -25766
rect -77599 -25810 -77555 -25766
rect -77499 -25810 -77455 -25766
rect -77399 -25810 -77355 -25766
rect -77299 -25810 -77255 -25766
rect -76799 -25810 -76755 -25766
rect -76699 -25810 -76655 -25766
rect -76599 -25810 -76555 -25766
rect -76499 -25810 -76455 -25766
rect -76399 -25810 -76355 -25766
rect -76299 -25810 -76255 -25766
rect -76199 -25810 -76155 -25766
rect -76099 -25810 -76055 -25766
rect -75999 -25810 -75955 -25766
rect -75899 -25810 -75855 -25766
rect -75799 -25810 -75755 -25766
rect -75699 -25810 -75655 -25766
rect -75599 -25810 -75555 -25766
rect -75499 -25810 -75455 -25766
rect -75399 -25810 -75355 -25766
rect -75299 -25810 -75255 -25766
rect -82799 -25910 -82755 -25866
rect -82699 -25910 -82655 -25866
rect -82599 -25910 -82555 -25866
rect -82499 -25910 -82455 -25866
rect -82399 -25910 -82355 -25866
rect -82299 -25910 -82255 -25866
rect -82199 -25910 -82155 -25866
rect -82099 -25910 -82055 -25866
rect -81999 -25910 -81955 -25866
rect -81899 -25910 -81855 -25866
rect -81799 -25910 -81755 -25866
rect -81699 -25910 -81655 -25866
rect -81599 -25910 -81555 -25866
rect -81499 -25910 -81455 -25866
rect -81399 -25910 -81355 -25866
rect -81299 -25910 -81255 -25866
rect -80799 -25910 -80755 -25866
rect -80699 -25910 -80655 -25866
rect -80599 -25910 -80555 -25866
rect -80499 -25910 -80455 -25866
rect -80399 -25910 -80355 -25866
rect -80299 -25910 -80255 -25866
rect -80199 -25910 -80155 -25866
rect -80099 -25910 -80055 -25866
rect -79999 -25910 -79955 -25866
rect -79899 -25910 -79855 -25866
rect -79799 -25910 -79755 -25866
rect -79699 -25910 -79655 -25866
rect -79599 -25910 -79555 -25866
rect -79499 -25910 -79455 -25866
rect -79399 -25910 -79355 -25866
rect -79299 -25910 -79255 -25866
rect -78799 -25910 -78755 -25866
rect -78699 -25910 -78655 -25866
rect -78599 -25910 -78555 -25866
rect -78499 -25910 -78455 -25866
rect -78399 -25910 -78355 -25866
rect -78299 -25910 -78255 -25866
rect -78199 -25910 -78155 -25866
rect -78099 -25910 -78055 -25866
rect -77999 -25910 -77955 -25866
rect -77899 -25910 -77855 -25866
rect -77799 -25910 -77755 -25866
rect -77699 -25910 -77655 -25866
rect -77599 -25910 -77555 -25866
rect -77499 -25910 -77455 -25866
rect -77399 -25910 -77355 -25866
rect -77299 -25910 -77255 -25866
rect -76799 -25910 -76755 -25866
rect -76699 -25910 -76655 -25866
rect -76599 -25910 -76555 -25866
rect -76499 -25910 -76455 -25866
rect -76399 -25910 -76355 -25866
rect -76299 -25910 -76255 -25866
rect -76199 -25910 -76155 -25866
rect -76099 -25910 -76055 -25866
rect -75999 -25910 -75955 -25866
rect -75899 -25910 -75855 -25866
rect -75799 -25910 -75755 -25866
rect -75699 -25910 -75655 -25866
rect -75599 -25910 -75555 -25866
rect -75499 -25910 -75455 -25866
rect -75399 -25910 -75355 -25866
rect -75299 -25910 -75255 -25866
rect 109305 -51181 109349 -51137
rect 109405 -51181 109449 -51137
rect 109505 -51181 109549 -51137
rect 109605 -51181 109649 -51137
rect 109705 -51181 109749 -51137
rect 109805 -51181 109849 -51137
rect 109905 -51181 109949 -51137
rect 110005 -51181 110049 -51137
rect 110105 -51181 110149 -51137
rect 110205 -51181 110249 -51137
rect 110305 -51181 110349 -51137
rect 110405 -51181 110449 -51137
rect 110505 -51181 110549 -51137
rect 110605 -51181 110649 -51137
rect 110705 -51181 110749 -51137
rect 110805 -51181 110849 -51137
rect 111305 -51181 111349 -51137
rect 111405 -51181 111449 -51137
rect 111505 -51181 111549 -51137
rect 111605 -51181 111649 -51137
rect 111705 -51181 111749 -51137
rect 111805 -51181 111849 -51137
rect 111905 -51181 111949 -51137
rect 112005 -51181 112049 -51137
rect 112105 -51181 112149 -51137
rect 112205 -51181 112249 -51137
rect 112305 -51181 112349 -51137
rect 112405 -51181 112449 -51137
rect 112505 -51181 112549 -51137
rect 112605 -51181 112649 -51137
rect 112705 -51181 112749 -51137
rect 112805 -51181 112849 -51137
rect 113305 -51181 113349 -51137
rect 113405 -51181 113449 -51137
rect 113505 -51181 113549 -51137
rect 113605 -51181 113649 -51137
rect 113705 -51181 113749 -51137
rect 113805 -51181 113849 -51137
rect 113905 -51181 113949 -51137
rect 114005 -51181 114049 -51137
rect 114105 -51181 114149 -51137
rect 114205 -51181 114249 -51137
rect 114305 -51181 114349 -51137
rect 114405 -51181 114449 -51137
rect 114505 -51181 114549 -51137
rect 114605 -51181 114649 -51137
rect 114705 -51181 114749 -51137
rect 114805 -51181 114849 -51137
rect 115305 -51181 115349 -51137
rect 115405 -51181 115449 -51137
rect 115505 -51181 115549 -51137
rect 115605 -51181 115649 -51137
rect 115705 -51181 115749 -51137
rect 115805 -51181 115849 -51137
rect 115905 -51181 115949 -51137
rect 116005 -51181 116049 -51137
rect 116105 -51181 116149 -51137
rect 116205 -51181 116249 -51137
rect 116305 -51181 116349 -51137
rect 116405 -51181 116449 -51137
rect 116505 -51181 116549 -51137
rect 116605 -51181 116649 -51137
rect 116705 -51181 116749 -51137
rect 116805 -51181 116849 -51137
rect 109305 -51281 109349 -51237
rect 109405 -51281 109449 -51237
rect 109505 -51281 109549 -51237
rect 109605 -51281 109649 -51237
rect 109705 -51281 109749 -51237
rect 109805 -51281 109849 -51237
rect 109905 -51281 109949 -51237
rect 110005 -51281 110049 -51237
rect 110105 -51281 110149 -51237
rect 110205 -51281 110249 -51237
rect 110305 -51281 110349 -51237
rect 110405 -51281 110449 -51237
rect 110505 -51281 110549 -51237
rect 110605 -51281 110649 -51237
rect 110705 -51281 110749 -51237
rect 110805 -51281 110849 -51237
rect 111305 -51281 111349 -51237
rect 111405 -51281 111449 -51237
rect 111505 -51281 111549 -51237
rect 111605 -51281 111649 -51237
rect 111705 -51281 111749 -51237
rect 111805 -51281 111849 -51237
rect 111905 -51281 111949 -51237
rect 112005 -51281 112049 -51237
rect 112105 -51281 112149 -51237
rect 112205 -51281 112249 -51237
rect 112305 -51281 112349 -51237
rect 112405 -51281 112449 -51237
rect 112505 -51281 112549 -51237
rect 112605 -51281 112649 -51237
rect 112705 -51281 112749 -51237
rect 112805 -51281 112849 -51237
rect 113305 -51281 113349 -51237
rect 113405 -51281 113449 -51237
rect 113505 -51281 113549 -51237
rect 113605 -51281 113649 -51237
rect 113705 -51281 113749 -51237
rect 113805 -51281 113849 -51237
rect 113905 -51281 113949 -51237
rect 114005 -51281 114049 -51237
rect 114105 -51281 114149 -51237
rect 114205 -51281 114249 -51237
rect 114305 -51281 114349 -51237
rect 114405 -51281 114449 -51237
rect 114505 -51281 114549 -51237
rect 114605 -51281 114649 -51237
rect 114705 -51281 114749 -51237
rect 114805 -51281 114849 -51237
rect 115305 -51281 115349 -51237
rect 115405 -51281 115449 -51237
rect 115505 -51281 115549 -51237
rect 115605 -51281 115649 -51237
rect 115705 -51281 115749 -51237
rect 115805 -51281 115849 -51237
rect 115905 -51281 115949 -51237
rect 116005 -51281 116049 -51237
rect 116105 -51281 116149 -51237
rect 116205 -51281 116249 -51237
rect 116305 -51281 116349 -51237
rect 116405 -51281 116449 -51237
rect 116505 -51281 116549 -51237
rect 116605 -51281 116649 -51237
rect 116705 -51281 116749 -51237
rect 116805 -51281 116849 -51237
rect 109305 -51381 109349 -51337
rect 109405 -51381 109449 -51337
rect 109505 -51381 109549 -51337
rect 109605 -51381 109649 -51337
rect 109705 -51381 109749 -51337
rect 109805 -51381 109849 -51337
rect 109905 -51381 109949 -51337
rect 110005 -51381 110049 -51337
rect 110105 -51381 110149 -51337
rect 110205 -51381 110249 -51337
rect 110305 -51381 110349 -51337
rect 110405 -51381 110449 -51337
rect 110505 -51381 110549 -51337
rect 110605 -51381 110649 -51337
rect 110705 -51381 110749 -51337
rect 110805 -51381 110849 -51337
rect 111305 -51381 111349 -51337
rect 111405 -51381 111449 -51337
rect 111505 -51381 111549 -51337
rect 111605 -51381 111649 -51337
rect 111705 -51381 111749 -51337
rect 111805 -51381 111849 -51337
rect 111905 -51381 111949 -51337
rect 112005 -51381 112049 -51337
rect 112105 -51381 112149 -51337
rect 112205 -51381 112249 -51337
rect 112305 -51381 112349 -51337
rect 112405 -51381 112449 -51337
rect 112505 -51381 112549 -51337
rect 112605 -51381 112649 -51337
rect 112705 -51381 112749 -51337
rect 112805 -51381 112849 -51337
rect 113305 -51381 113349 -51337
rect 113405 -51381 113449 -51337
rect 113505 -51381 113549 -51337
rect 113605 -51381 113649 -51337
rect 113705 -51381 113749 -51337
rect 113805 -51381 113849 -51337
rect 113905 -51381 113949 -51337
rect 114005 -51381 114049 -51337
rect 114105 -51381 114149 -51337
rect 114205 -51381 114249 -51337
rect 114305 -51381 114349 -51337
rect 114405 -51381 114449 -51337
rect 114505 -51381 114549 -51337
rect 114605 -51381 114649 -51337
rect 114705 -51381 114749 -51337
rect 114805 -51381 114849 -51337
rect 115305 -51381 115349 -51337
rect 115405 -51381 115449 -51337
rect 115505 -51381 115549 -51337
rect 115605 -51381 115649 -51337
rect 115705 -51381 115749 -51337
rect 115805 -51381 115849 -51337
rect 115905 -51381 115949 -51337
rect 116005 -51381 116049 -51337
rect 116105 -51381 116149 -51337
rect 116205 -51381 116249 -51337
rect 116305 -51381 116349 -51337
rect 116405 -51381 116449 -51337
rect 116505 -51381 116549 -51337
rect 116605 -51381 116649 -51337
rect 116705 -51381 116749 -51337
rect 116805 -51381 116849 -51337
rect 109305 -51481 109349 -51437
rect 109405 -51481 109449 -51437
rect 109505 -51481 109549 -51437
rect 109605 -51481 109649 -51437
rect 109705 -51481 109749 -51437
rect 109805 -51481 109849 -51437
rect 109905 -51481 109949 -51437
rect 110005 -51481 110049 -51437
rect 110105 -51481 110149 -51437
rect 110205 -51481 110249 -51437
rect 110305 -51481 110349 -51437
rect 110405 -51481 110449 -51437
rect 110505 -51481 110549 -51437
rect 110605 -51481 110649 -51437
rect 110705 -51481 110749 -51437
rect 110805 -51481 110849 -51437
rect 111305 -51481 111349 -51437
rect 111405 -51481 111449 -51437
rect 111505 -51481 111549 -51437
rect 111605 -51481 111649 -51437
rect 111705 -51481 111749 -51437
rect 111805 -51481 111849 -51437
rect 111905 -51481 111949 -51437
rect 112005 -51481 112049 -51437
rect 112105 -51481 112149 -51437
rect 112205 -51481 112249 -51437
rect 112305 -51481 112349 -51437
rect 112405 -51481 112449 -51437
rect 112505 -51481 112549 -51437
rect 112605 -51481 112649 -51437
rect 112705 -51481 112749 -51437
rect 112805 -51481 112849 -51437
rect 113305 -51481 113349 -51437
rect 113405 -51481 113449 -51437
rect 113505 -51481 113549 -51437
rect 113605 -51481 113649 -51437
rect 113705 -51481 113749 -51437
rect 113805 -51481 113849 -51437
rect 113905 -51481 113949 -51437
rect 114005 -51481 114049 -51437
rect 114105 -51481 114149 -51437
rect 114205 -51481 114249 -51437
rect 114305 -51481 114349 -51437
rect 114405 -51481 114449 -51437
rect 114505 -51481 114549 -51437
rect 114605 -51481 114649 -51437
rect 114705 -51481 114749 -51437
rect 114805 -51481 114849 -51437
rect 115305 -51481 115349 -51437
rect 115405 -51481 115449 -51437
rect 115505 -51481 115549 -51437
rect 115605 -51481 115649 -51437
rect 115705 -51481 115749 -51437
rect 115805 -51481 115849 -51437
rect 115905 -51481 115949 -51437
rect 116005 -51481 116049 -51437
rect 116105 -51481 116149 -51437
rect 116205 -51481 116249 -51437
rect 116305 -51481 116349 -51437
rect 116405 -51481 116449 -51437
rect 116505 -51481 116549 -51437
rect 116605 -51481 116649 -51437
rect 116705 -51481 116749 -51437
rect 116805 -51481 116849 -51437
rect 109305 -51581 109349 -51537
rect 109405 -51581 109449 -51537
rect 109505 -51581 109549 -51537
rect 109605 -51581 109649 -51537
rect 109705 -51581 109749 -51537
rect 109805 -51581 109849 -51537
rect 109905 -51581 109949 -51537
rect 110005 -51581 110049 -51537
rect 110105 -51581 110149 -51537
rect 110205 -51581 110249 -51537
rect 110305 -51581 110349 -51537
rect 110405 -51581 110449 -51537
rect 110505 -51581 110549 -51537
rect 110605 -51581 110649 -51537
rect 110705 -51581 110749 -51537
rect 110805 -51581 110849 -51537
rect 111305 -51581 111349 -51537
rect 111405 -51581 111449 -51537
rect 111505 -51581 111549 -51537
rect 111605 -51581 111649 -51537
rect 111705 -51581 111749 -51537
rect 111805 -51581 111849 -51537
rect 111905 -51581 111949 -51537
rect 112005 -51581 112049 -51537
rect 112105 -51581 112149 -51537
rect 112205 -51581 112249 -51537
rect 112305 -51581 112349 -51537
rect 112405 -51581 112449 -51537
rect 112505 -51581 112549 -51537
rect 112605 -51581 112649 -51537
rect 112705 -51581 112749 -51537
rect 112805 -51581 112849 -51537
rect 113305 -51581 113349 -51537
rect 113405 -51581 113449 -51537
rect 113505 -51581 113549 -51537
rect 113605 -51581 113649 -51537
rect 113705 -51581 113749 -51537
rect 113805 -51581 113849 -51537
rect 113905 -51581 113949 -51537
rect 114005 -51581 114049 -51537
rect 114105 -51581 114149 -51537
rect 114205 -51581 114249 -51537
rect 114305 -51581 114349 -51537
rect 114405 -51581 114449 -51537
rect 114505 -51581 114549 -51537
rect 114605 -51581 114649 -51537
rect 114705 -51581 114749 -51537
rect 114805 -51581 114849 -51537
rect 115305 -51581 115349 -51537
rect 115405 -51581 115449 -51537
rect 115505 -51581 115549 -51537
rect 115605 -51581 115649 -51537
rect 115705 -51581 115749 -51537
rect 115805 -51581 115849 -51537
rect 115905 -51581 115949 -51537
rect 116005 -51581 116049 -51537
rect 116105 -51581 116149 -51537
rect 116205 -51581 116249 -51537
rect 116305 -51581 116349 -51537
rect 116405 -51581 116449 -51537
rect 116505 -51581 116549 -51537
rect 116605 -51581 116649 -51537
rect 116705 -51581 116749 -51537
rect 116805 -51581 116849 -51537
rect 109305 -51681 109349 -51637
rect 109405 -51681 109449 -51637
rect 109505 -51681 109549 -51637
rect 109605 -51681 109649 -51637
rect 109705 -51681 109749 -51637
rect 109805 -51681 109849 -51637
rect 109905 -51681 109949 -51637
rect 110005 -51681 110049 -51637
rect 110105 -51681 110149 -51637
rect 110205 -51681 110249 -51637
rect 110305 -51681 110349 -51637
rect 110405 -51681 110449 -51637
rect 110505 -51681 110549 -51637
rect 110605 -51681 110649 -51637
rect 110705 -51681 110749 -51637
rect 110805 -51681 110849 -51637
rect 111305 -51681 111349 -51637
rect 111405 -51681 111449 -51637
rect 111505 -51681 111549 -51637
rect 111605 -51681 111649 -51637
rect 111705 -51681 111749 -51637
rect 111805 -51681 111849 -51637
rect 111905 -51681 111949 -51637
rect 112005 -51681 112049 -51637
rect 112105 -51681 112149 -51637
rect 112205 -51681 112249 -51637
rect 112305 -51681 112349 -51637
rect 112405 -51681 112449 -51637
rect 112505 -51681 112549 -51637
rect 112605 -51681 112649 -51637
rect 112705 -51681 112749 -51637
rect 112805 -51681 112849 -51637
rect 113305 -51681 113349 -51637
rect 113405 -51681 113449 -51637
rect 113505 -51681 113549 -51637
rect 113605 -51681 113649 -51637
rect 113705 -51681 113749 -51637
rect 113805 -51681 113849 -51637
rect 113905 -51681 113949 -51637
rect 114005 -51681 114049 -51637
rect 114105 -51681 114149 -51637
rect 114205 -51681 114249 -51637
rect 114305 -51681 114349 -51637
rect 114405 -51681 114449 -51637
rect 114505 -51681 114549 -51637
rect 114605 -51681 114649 -51637
rect 114705 -51681 114749 -51637
rect 114805 -51681 114849 -51637
rect 115305 -51681 115349 -51637
rect 115405 -51681 115449 -51637
rect 115505 -51681 115549 -51637
rect 115605 -51681 115649 -51637
rect 115705 -51681 115749 -51637
rect 115805 -51681 115849 -51637
rect 115905 -51681 115949 -51637
rect 116005 -51681 116049 -51637
rect 116105 -51681 116149 -51637
rect 116205 -51681 116249 -51637
rect 116305 -51681 116349 -51637
rect 116405 -51681 116449 -51637
rect 116505 -51681 116549 -51637
rect 116605 -51681 116649 -51637
rect 116705 -51681 116749 -51637
rect 116805 -51681 116849 -51637
rect 109305 -51781 109349 -51737
rect 109405 -51781 109449 -51737
rect 109505 -51781 109549 -51737
rect 109605 -51781 109649 -51737
rect 109705 -51781 109749 -51737
rect 109805 -51781 109849 -51737
rect 109905 -51781 109949 -51737
rect 110005 -51781 110049 -51737
rect 110105 -51781 110149 -51737
rect 110205 -51781 110249 -51737
rect 110305 -51781 110349 -51737
rect 110405 -51781 110449 -51737
rect 110505 -51781 110549 -51737
rect 110605 -51781 110649 -51737
rect 110705 -51781 110749 -51737
rect 110805 -51781 110849 -51737
rect 111305 -51781 111349 -51737
rect 111405 -51781 111449 -51737
rect 111505 -51781 111549 -51737
rect 111605 -51781 111649 -51737
rect 111705 -51781 111749 -51737
rect 111805 -51781 111849 -51737
rect 111905 -51781 111949 -51737
rect 112005 -51781 112049 -51737
rect 112105 -51781 112149 -51737
rect 112205 -51781 112249 -51737
rect 112305 -51781 112349 -51737
rect 112405 -51781 112449 -51737
rect 112505 -51781 112549 -51737
rect 112605 -51781 112649 -51737
rect 112705 -51781 112749 -51737
rect 112805 -51781 112849 -51737
rect 113305 -51781 113349 -51737
rect 113405 -51781 113449 -51737
rect 113505 -51781 113549 -51737
rect 113605 -51781 113649 -51737
rect 113705 -51781 113749 -51737
rect 113805 -51781 113849 -51737
rect 113905 -51781 113949 -51737
rect 114005 -51781 114049 -51737
rect 114105 -51781 114149 -51737
rect 114205 -51781 114249 -51737
rect 114305 -51781 114349 -51737
rect 114405 -51781 114449 -51737
rect 114505 -51781 114549 -51737
rect 114605 -51781 114649 -51737
rect 114705 -51781 114749 -51737
rect 114805 -51781 114849 -51737
rect 115305 -51781 115349 -51737
rect 115405 -51781 115449 -51737
rect 115505 -51781 115549 -51737
rect 115605 -51781 115649 -51737
rect 115705 -51781 115749 -51737
rect 115805 -51781 115849 -51737
rect 115905 -51781 115949 -51737
rect 116005 -51781 116049 -51737
rect 116105 -51781 116149 -51737
rect 116205 -51781 116249 -51737
rect 116305 -51781 116349 -51737
rect 116405 -51781 116449 -51737
rect 116505 -51781 116549 -51737
rect 116605 -51781 116649 -51737
rect 116705 -51781 116749 -51737
rect 116805 -51781 116849 -51737
rect 109305 -51881 109349 -51837
rect 109405 -51881 109449 -51837
rect 109505 -51881 109549 -51837
rect 109605 -51881 109649 -51837
rect 109705 -51881 109749 -51837
rect 109805 -51881 109849 -51837
rect 109905 -51881 109949 -51837
rect 110005 -51881 110049 -51837
rect 110105 -51881 110149 -51837
rect 110205 -51881 110249 -51837
rect 110305 -51881 110349 -51837
rect 110405 -51881 110449 -51837
rect 110505 -51881 110549 -51837
rect 110605 -51881 110649 -51837
rect 110705 -51881 110749 -51837
rect 110805 -51881 110849 -51837
rect 111305 -51881 111349 -51837
rect 111405 -51881 111449 -51837
rect 111505 -51881 111549 -51837
rect 111605 -51881 111649 -51837
rect 111705 -51881 111749 -51837
rect 111805 -51881 111849 -51837
rect 111905 -51881 111949 -51837
rect 112005 -51881 112049 -51837
rect 112105 -51881 112149 -51837
rect 112205 -51881 112249 -51837
rect 112305 -51881 112349 -51837
rect 112405 -51881 112449 -51837
rect 112505 -51881 112549 -51837
rect 112605 -51881 112649 -51837
rect 112705 -51881 112749 -51837
rect 112805 -51881 112849 -51837
rect 113305 -51881 113349 -51837
rect 113405 -51881 113449 -51837
rect 113505 -51881 113549 -51837
rect 113605 -51881 113649 -51837
rect 113705 -51881 113749 -51837
rect 113805 -51881 113849 -51837
rect 113905 -51881 113949 -51837
rect 114005 -51881 114049 -51837
rect 114105 -51881 114149 -51837
rect 114205 -51881 114249 -51837
rect 114305 -51881 114349 -51837
rect 114405 -51881 114449 -51837
rect 114505 -51881 114549 -51837
rect 114605 -51881 114649 -51837
rect 114705 -51881 114749 -51837
rect 114805 -51881 114849 -51837
rect 115305 -51881 115349 -51837
rect 115405 -51881 115449 -51837
rect 115505 -51881 115549 -51837
rect 115605 -51881 115649 -51837
rect 115705 -51881 115749 -51837
rect 115805 -51881 115849 -51837
rect 115905 -51881 115949 -51837
rect 116005 -51881 116049 -51837
rect 116105 -51881 116149 -51837
rect 116205 -51881 116249 -51837
rect 116305 -51881 116349 -51837
rect 116405 -51881 116449 -51837
rect 116505 -51881 116549 -51837
rect 116605 -51881 116649 -51837
rect 116705 -51881 116749 -51837
rect 116805 -51881 116849 -51837
rect 109305 -51981 109349 -51937
rect 109405 -51981 109449 -51937
rect 109505 -51981 109549 -51937
rect 109605 -51981 109649 -51937
rect 109705 -51981 109749 -51937
rect 109805 -51981 109849 -51937
rect 109905 -51981 109949 -51937
rect 110005 -51981 110049 -51937
rect 110105 -51981 110149 -51937
rect 110205 -51981 110249 -51937
rect 110305 -51981 110349 -51937
rect 110405 -51981 110449 -51937
rect 110505 -51981 110549 -51937
rect 110605 -51981 110649 -51937
rect 110705 -51981 110749 -51937
rect 110805 -51981 110849 -51937
rect 111305 -51981 111349 -51937
rect 111405 -51981 111449 -51937
rect 111505 -51981 111549 -51937
rect 111605 -51981 111649 -51937
rect 111705 -51981 111749 -51937
rect 111805 -51981 111849 -51937
rect 111905 -51981 111949 -51937
rect 112005 -51981 112049 -51937
rect 112105 -51981 112149 -51937
rect 112205 -51981 112249 -51937
rect 112305 -51981 112349 -51937
rect 112405 -51981 112449 -51937
rect 112505 -51981 112549 -51937
rect 112605 -51981 112649 -51937
rect 112705 -51981 112749 -51937
rect 112805 -51981 112849 -51937
rect 113305 -51981 113349 -51937
rect 113405 -51981 113449 -51937
rect 113505 -51981 113549 -51937
rect 113605 -51981 113649 -51937
rect 113705 -51981 113749 -51937
rect 113805 -51981 113849 -51937
rect 113905 -51981 113949 -51937
rect 114005 -51981 114049 -51937
rect 114105 -51981 114149 -51937
rect 114205 -51981 114249 -51937
rect 114305 -51981 114349 -51937
rect 114405 -51981 114449 -51937
rect 114505 -51981 114549 -51937
rect 114605 -51981 114649 -51937
rect 114705 -51981 114749 -51937
rect 114805 -51981 114849 -51937
rect 115305 -51981 115349 -51937
rect 115405 -51981 115449 -51937
rect 115505 -51981 115549 -51937
rect 115605 -51981 115649 -51937
rect 115705 -51981 115749 -51937
rect 115805 -51981 115849 -51937
rect 115905 -51981 115949 -51937
rect 116005 -51981 116049 -51937
rect 116105 -51981 116149 -51937
rect 116205 -51981 116249 -51937
rect 116305 -51981 116349 -51937
rect 116405 -51981 116449 -51937
rect 116505 -51981 116549 -51937
rect 116605 -51981 116649 -51937
rect 116705 -51981 116749 -51937
rect 116805 -51981 116849 -51937
rect 109305 -52081 109349 -52037
rect 109405 -52081 109449 -52037
rect 109505 -52081 109549 -52037
rect 109605 -52081 109649 -52037
rect 109705 -52081 109749 -52037
rect 109805 -52081 109849 -52037
rect 109905 -52081 109949 -52037
rect 110005 -52081 110049 -52037
rect 110105 -52081 110149 -52037
rect 110205 -52081 110249 -52037
rect 110305 -52081 110349 -52037
rect 110405 -52081 110449 -52037
rect 110505 -52081 110549 -52037
rect 110605 -52081 110649 -52037
rect 110705 -52081 110749 -52037
rect 110805 -52081 110849 -52037
rect 111305 -52081 111349 -52037
rect 111405 -52081 111449 -52037
rect 111505 -52081 111549 -52037
rect 111605 -52081 111649 -52037
rect 111705 -52081 111749 -52037
rect 111805 -52081 111849 -52037
rect 111905 -52081 111949 -52037
rect 112005 -52081 112049 -52037
rect 112105 -52081 112149 -52037
rect 112205 -52081 112249 -52037
rect 112305 -52081 112349 -52037
rect 112405 -52081 112449 -52037
rect 112505 -52081 112549 -52037
rect 112605 -52081 112649 -52037
rect 112705 -52081 112749 -52037
rect 112805 -52081 112849 -52037
rect 113305 -52081 113349 -52037
rect 113405 -52081 113449 -52037
rect 113505 -52081 113549 -52037
rect 113605 -52081 113649 -52037
rect 113705 -52081 113749 -52037
rect 113805 -52081 113849 -52037
rect 113905 -52081 113949 -52037
rect 114005 -52081 114049 -52037
rect 114105 -52081 114149 -52037
rect 114205 -52081 114249 -52037
rect 114305 -52081 114349 -52037
rect 114405 -52081 114449 -52037
rect 114505 -52081 114549 -52037
rect 114605 -52081 114649 -52037
rect 114705 -52081 114749 -52037
rect 114805 -52081 114849 -52037
rect 115305 -52081 115349 -52037
rect 115405 -52081 115449 -52037
rect 115505 -52081 115549 -52037
rect 115605 -52081 115649 -52037
rect 115705 -52081 115749 -52037
rect 115805 -52081 115849 -52037
rect 115905 -52081 115949 -52037
rect 116005 -52081 116049 -52037
rect 116105 -52081 116149 -52037
rect 116205 -52081 116249 -52037
rect 116305 -52081 116349 -52037
rect 116405 -52081 116449 -52037
rect 116505 -52081 116549 -52037
rect 116605 -52081 116649 -52037
rect 116705 -52081 116749 -52037
rect 116805 -52081 116849 -52037
rect 109305 -52181 109349 -52137
rect 109405 -52181 109449 -52137
rect 109505 -52181 109549 -52137
rect 109605 -52181 109649 -52137
rect 109705 -52181 109749 -52137
rect 109805 -52181 109849 -52137
rect 109905 -52181 109949 -52137
rect 110005 -52181 110049 -52137
rect 110105 -52181 110149 -52137
rect 110205 -52181 110249 -52137
rect 110305 -52181 110349 -52137
rect 110405 -52181 110449 -52137
rect 110505 -52181 110549 -52137
rect 110605 -52181 110649 -52137
rect 110705 -52181 110749 -52137
rect 110805 -52181 110849 -52137
rect 111305 -52181 111349 -52137
rect 111405 -52181 111449 -52137
rect 111505 -52181 111549 -52137
rect 111605 -52181 111649 -52137
rect 111705 -52181 111749 -52137
rect 111805 -52181 111849 -52137
rect 111905 -52181 111949 -52137
rect 112005 -52181 112049 -52137
rect 112105 -52181 112149 -52137
rect 112205 -52181 112249 -52137
rect 112305 -52181 112349 -52137
rect 112405 -52181 112449 -52137
rect 112505 -52181 112549 -52137
rect 112605 -52181 112649 -52137
rect 112705 -52181 112749 -52137
rect 112805 -52181 112849 -52137
rect 113305 -52181 113349 -52137
rect 113405 -52181 113449 -52137
rect 113505 -52181 113549 -52137
rect 113605 -52181 113649 -52137
rect 113705 -52181 113749 -52137
rect 113805 -52181 113849 -52137
rect 113905 -52181 113949 -52137
rect 114005 -52181 114049 -52137
rect 114105 -52181 114149 -52137
rect 114205 -52181 114249 -52137
rect 114305 -52181 114349 -52137
rect 114405 -52181 114449 -52137
rect 114505 -52181 114549 -52137
rect 114605 -52181 114649 -52137
rect 114705 -52181 114749 -52137
rect 114805 -52181 114849 -52137
rect 115305 -52181 115349 -52137
rect 115405 -52181 115449 -52137
rect 115505 -52181 115549 -52137
rect 115605 -52181 115649 -52137
rect 115705 -52181 115749 -52137
rect 115805 -52181 115849 -52137
rect 115905 -52181 115949 -52137
rect 116005 -52181 116049 -52137
rect 116105 -52181 116149 -52137
rect 116205 -52181 116249 -52137
rect 116305 -52181 116349 -52137
rect 116405 -52181 116449 -52137
rect 116505 -52181 116549 -52137
rect 116605 -52181 116649 -52137
rect 116705 -52181 116749 -52137
rect 116805 -52181 116849 -52137
rect 109305 -52281 109349 -52237
rect 109405 -52281 109449 -52237
rect 109505 -52281 109549 -52237
rect 109605 -52281 109649 -52237
rect 109705 -52281 109749 -52237
rect 109805 -52281 109849 -52237
rect 109905 -52281 109949 -52237
rect 110005 -52281 110049 -52237
rect 110105 -52281 110149 -52237
rect 110205 -52281 110249 -52237
rect 110305 -52281 110349 -52237
rect 110405 -52281 110449 -52237
rect 110505 -52281 110549 -52237
rect 110605 -52281 110649 -52237
rect 110705 -52281 110749 -52237
rect 110805 -52281 110849 -52237
rect 111305 -52281 111349 -52237
rect 111405 -52281 111449 -52237
rect 111505 -52281 111549 -52237
rect 111605 -52281 111649 -52237
rect 111705 -52281 111749 -52237
rect 111805 -52281 111849 -52237
rect 111905 -52281 111949 -52237
rect 112005 -52281 112049 -52237
rect 112105 -52281 112149 -52237
rect 112205 -52281 112249 -52237
rect 112305 -52281 112349 -52237
rect 112405 -52281 112449 -52237
rect 112505 -52281 112549 -52237
rect 112605 -52281 112649 -52237
rect 112705 -52281 112749 -52237
rect 112805 -52281 112849 -52237
rect 113305 -52281 113349 -52237
rect 113405 -52281 113449 -52237
rect 113505 -52281 113549 -52237
rect 113605 -52281 113649 -52237
rect 113705 -52281 113749 -52237
rect 113805 -52281 113849 -52237
rect 113905 -52281 113949 -52237
rect 114005 -52281 114049 -52237
rect 114105 -52281 114149 -52237
rect 114205 -52281 114249 -52237
rect 114305 -52281 114349 -52237
rect 114405 -52281 114449 -52237
rect 114505 -52281 114549 -52237
rect 114605 -52281 114649 -52237
rect 114705 -52281 114749 -52237
rect 114805 -52281 114849 -52237
rect 115305 -52281 115349 -52237
rect 115405 -52281 115449 -52237
rect 115505 -52281 115549 -52237
rect 115605 -52281 115649 -52237
rect 115705 -52281 115749 -52237
rect 115805 -52281 115849 -52237
rect 115905 -52281 115949 -52237
rect 116005 -52281 116049 -52237
rect 116105 -52281 116149 -52237
rect 116205 -52281 116249 -52237
rect 116305 -52281 116349 -52237
rect 116405 -52281 116449 -52237
rect 116505 -52281 116549 -52237
rect 116605 -52281 116649 -52237
rect 116705 -52281 116749 -52237
rect 116805 -52281 116849 -52237
rect 109305 -52381 109349 -52337
rect 109405 -52381 109449 -52337
rect 109505 -52381 109549 -52337
rect 109605 -52381 109649 -52337
rect 109705 -52381 109749 -52337
rect 109805 -52381 109849 -52337
rect 109905 -52381 109949 -52337
rect 110005 -52381 110049 -52337
rect 110105 -52381 110149 -52337
rect 110205 -52381 110249 -52337
rect 110305 -52381 110349 -52337
rect 110405 -52381 110449 -52337
rect 110505 -52381 110549 -52337
rect 110605 -52381 110649 -52337
rect 110705 -52381 110749 -52337
rect 110805 -52381 110849 -52337
rect 111305 -52381 111349 -52337
rect 111405 -52381 111449 -52337
rect 111505 -52381 111549 -52337
rect 111605 -52381 111649 -52337
rect 111705 -52381 111749 -52337
rect 111805 -52381 111849 -52337
rect 111905 -52381 111949 -52337
rect 112005 -52381 112049 -52337
rect 112105 -52381 112149 -52337
rect 112205 -52381 112249 -52337
rect 112305 -52381 112349 -52337
rect 112405 -52381 112449 -52337
rect 112505 -52381 112549 -52337
rect 112605 -52381 112649 -52337
rect 112705 -52381 112749 -52337
rect 112805 -52381 112849 -52337
rect 113305 -52381 113349 -52337
rect 113405 -52381 113449 -52337
rect 113505 -52381 113549 -52337
rect 113605 -52381 113649 -52337
rect 113705 -52381 113749 -52337
rect 113805 -52381 113849 -52337
rect 113905 -52381 113949 -52337
rect 114005 -52381 114049 -52337
rect 114105 -52381 114149 -52337
rect 114205 -52381 114249 -52337
rect 114305 -52381 114349 -52337
rect 114405 -52381 114449 -52337
rect 114505 -52381 114549 -52337
rect 114605 -52381 114649 -52337
rect 114705 -52381 114749 -52337
rect 114805 -52381 114849 -52337
rect 115305 -52381 115349 -52337
rect 115405 -52381 115449 -52337
rect 115505 -52381 115549 -52337
rect 115605 -52381 115649 -52337
rect 115705 -52381 115749 -52337
rect 115805 -52381 115849 -52337
rect 115905 -52381 115949 -52337
rect 116005 -52381 116049 -52337
rect 116105 -52381 116149 -52337
rect 116205 -52381 116249 -52337
rect 116305 -52381 116349 -52337
rect 116405 -52381 116449 -52337
rect 116505 -52381 116549 -52337
rect 116605 -52381 116649 -52337
rect 116705 -52381 116749 -52337
rect 116805 -52381 116849 -52337
rect 109305 -52481 109349 -52437
rect 109405 -52481 109449 -52437
rect 109505 -52481 109549 -52437
rect 109605 -52481 109649 -52437
rect 109705 -52481 109749 -52437
rect 109805 -52481 109849 -52437
rect 109905 -52481 109949 -52437
rect 110005 -52481 110049 -52437
rect 110105 -52481 110149 -52437
rect 110205 -52481 110249 -52437
rect 110305 -52481 110349 -52437
rect 110405 -52481 110449 -52437
rect 110505 -52481 110549 -52437
rect 110605 -52481 110649 -52437
rect 110705 -52481 110749 -52437
rect 110805 -52481 110849 -52437
rect 111305 -52481 111349 -52437
rect 111405 -52481 111449 -52437
rect 111505 -52481 111549 -52437
rect 111605 -52481 111649 -52437
rect 111705 -52481 111749 -52437
rect 111805 -52481 111849 -52437
rect 111905 -52481 111949 -52437
rect 112005 -52481 112049 -52437
rect 112105 -52481 112149 -52437
rect 112205 -52481 112249 -52437
rect 112305 -52481 112349 -52437
rect 112405 -52481 112449 -52437
rect 112505 -52481 112549 -52437
rect 112605 -52481 112649 -52437
rect 112705 -52481 112749 -52437
rect 112805 -52481 112849 -52437
rect 113305 -52481 113349 -52437
rect 113405 -52481 113449 -52437
rect 113505 -52481 113549 -52437
rect 113605 -52481 113649 -52437
rect 113705 -52481 113749 -52437
rect 113805 -52481 113849 -52437
rect 113905 -52481 113949 -52437
rect 114005 -52481 114049 -52437
rect 114105 -52481 114149 -52437
rect 114205 -52481 114249 -52437
rect 114305 -52481 114349 -52437
rect 114405 -52481 114449 -52437
rect 114505 -52481 114549 -52437
rect 114605 -52481 114649 -52437
rect 114705 -52481 114749 -52437
rect 114805 -52481 114849 -52437
rect 115305 -52481 115349 -52437
rect 115405 -52481 115449 -52437
rect 115505 -52481 115549 -52437
rect 115605 -52481 115649 -52437
rect 115705 -52481 115749 -52437
rect 115805 -52481 115849 -52437
rect 115905 -52481 115949 -52437
rect 116005 -52481 116049 -52437
rect 116105 -52481 116149 -52437
rect 116205 -52481 116249 -52437
rect 116305 -52481 116349 -52437
rect 116405 -52481 116449 -52437
rect 116505 -52481 116549 -52437
rect 116605 -52481 116649 -52437
rect 116705 -52481 116749 -52437
rect 116805 -52481 116849 -52437
rect 109305 -52581 109349 -52537
rect 109405 -52581 109449 -52537
rect 109505 -52581 109549 -52537
rect 109605 -52581 109649 -52537
rect 109705 -52581 109749 -52537
rect 109805 -52581 109849 -52537
rect 109905 -52581 109949 -52537
rect 110005 -52581 110049 -52537
rect 110105 -52581 110149 -52537
rect 110205 -52581 110249 -52537
rect 110305 -52581 110349 -52537
rect 110405 -52581 110449 -52537
rect 110505 -52581 110549 -52537
rect 110605 -52581 110649 -52537
rect 110705 -52581 110749 -52537
rect 110805 -52581 110849 -52537
rect 111305 -52581 111349 -52537
rect 111405 -52581 111449 -52537
rect 111505 -52581 111549 -52537
rect 111605 -52581 111649 -52537
rect 111705 -52581 111749 -52537
rect 111805 -52581 111849 -52537
rect 111905 -52581 111949 -52537
rect 112005 -52581 112049 -52537
rect 112105 -52581 112149 -52537
rect 112205 -52581 112249 -52537
rect 112305 -52581 112349 -52537
rect 112405 -52581 112449 -52537
rect 112505 -52581 112549 -52537
rect 112605 -52581 112649 -52537
rect 112705 -52581 112749 -52537
rect 112805 -52581 112849 -52537
rect 113305 -52581 113349 -52537
rect 113405 -52581 113449 -52537
rect 113505 -52581 113549 -52537
rect 113605 -52581 113649 -52537
rect 113705 -52581 113749 -52537
rect 113805 -52581 113849 -52537
rect 113905 -52581 113949 -52537
rect 114005 -52581 114049 -52537
rect 114105 -52581 114149 -52537
rect 114205 -52581 114249 -52537
rect 114305 -52581 114349 -52537
rect 114405 -52581 114449 -52537
rect 114505 -52581 114549 -52537
rect 114605 -52581 114649 -52537
rect 114705 -52581 114749 -52537
rect 114805 -52581 114849 -52537
rect 115305 -52581 115349 -52537
rect 115405 -52581 115449 -52537
rect 115505 -52581 115549 -52537
rect 115605 -52581 115649 -52537
rect 115705 -52581 115749 -52537
rect 115805 -52581 115849 -52537
rect 115905 -52581 115949 -52537
rect 116005 -52581 116049 -52537
rect 116105 -52581 116149 -52537
rect 116205 -52581 116249 -52537
rect 116305 -52581 116349 -52537
rect 116405 -52581 116449 -52537
rect 116505 -52581 116549 -52537
rect 116605 -52581 116649 -52537
rect 116705 -52581 116749 -52537
rect 116805 -52581 116849 -52537
rect 109305 -52681 109349 -52637
rect 109405 -52681 109449 -52637
rect 109505 -52681 109549 -52637
rect 109605 -52681 109649 -52637
rect 109705 -52681 109749 -52637
rect 109805 -52681 109849 -52637
rect 109905 -52681 109949 -52637
rect 110005 -52681 110049 -52637
rect 110105 -52681 110149 -52637
rect 110205 -52681 110249 -52637
rect 110305 -52681 110349 -52637
rect 110405 -52681 110449 -52637
rect 110505 -52681 110549 -52637
rect 110605 -52681 110649 -52637
rect 110705 -52681 110749 -52637
rect 110805 -52681 110849 -52637
rect 111305 -52681 111349 -52637
rect 111405 -52681 111449 -52637
rect 111505 -52681 111549 -52637
rect 111605 -52681 111649 -52637
rect 111705 -52681 111749 -52637
rect 111805 -52681 111849 -52637
rect 111905 -52681 111949 -52637
rect 112005 -52681 112049 -52637
rect 112105 -52681 112149 -52637
rect 112205 -52681 112249 -52637
rect 112305 -52681 112349 -52637
rect 112405 -52681 112449 -52637
rect 112505 -52681 112549 -52637
rect 112605 -52681 112649 -52637
rect 112705 -52681 112749 -52637
rect 112805 -52681 112849 -52637
rect 113305 -52681 113349 -52637
rect 113405 -52681 113449 -52637
rect 113505 -52681 113549 -52637
rect 113605 -52681 113649 -52637
rect 113705 -52681 113749 -52637
rect 113805 -52681 113849 -52637
rect 113905 -52681 113949 -52637
rect 114005 -52681 114049 -52637
rect 114105 -52681 114149 -52637
rect 114205 -52681 114249 -52637
rect 114305 -52681 114349 -52637
rect 114405 -52681 114449 -52637
rect 114505 -52681 114549 -52637
rect 114605 -52681 114649 -52637
rect 114705 -52681 114749 -52637
rect 114805 -52681 114849 -52637
rect 115305 -52681 115349 -52637
rect 115405 -52681 115449 -52637
rect 115505 -52681 115549 -52637
rect 115605 -52681 115649 -52637
rect 115705 -52681 115749 -52637
rect 115805 -52681 115849 -52637
rect 115905 -52681 115949 -52637
rect 116005 -52681 116049 -52637
rect 116105 -52681 116149 -52637
rect 116205 -52681 116249 -52637
rect 116305 -52681 116349 -52637
rect 116405 -52681 116449 -52637
rect 116505 -52681 116549 -52637
rect 116605 -52681 116649 -52637
rect 116705 -52681 116749 -52637
rect 116805 -52681 116849 -52637
rect 9236 -75232 9280 -75188
rect 9336 -75232 9380 -75188
rect 9436 -75232 9480 -75188
rect 9536 -75232 9580 -75188
rect 9636 -75232 9680 -75188
rect 9736 -75232 9780 -75188
rect 9836 -75232 9880 -75188
rect 9936 -75232 9980 -75188
rect 10036 -75232 10080 -75188
rect 10136 -75232 10180 -75188
rect 10236 -75232 10280 -75188
rect 10336 -75232 10380 -75188
rect 10436 -75232 10480 -75188
rect 10536 -75232 10580 -75188
rect 10636 -75232 10680 -75188
rect 10736 -75232 10780 -75188
rect 11236 -75232 11280 -75188
rect 11336 -75232 11380 -75188
rect 11436 -75232 11480 -75188
rect 11536 -75232 11580 -75188
rect 11636 -75232 11680 -75188
rect 11736 -75232 11780 -75188
rect 11836 -75232 11880 -75188
rect 11936 -75232 11980 -75188
rect 12036 -75232 12080 -75188
rect 12136 -75232 12180 -75188
rect 12236 -75232 12280 -75188
rect 12336 -75232 12380 -75188
rect 12436 -75232 12480 -75188
rect 12536 -75232 12580 -75188
rect 12636 -75232 12680 -75188
rect 12736 -75232 12780 -75188
rect 13236 -75232 13280 -75188
rect 13336 -75232 13380 -75188
rect 13436 -75232 13480 -75188
rect 13536 -75232 13580 -75188
rect 13636 -75232 13680 -75188
rect 13736 -75232 13780 -75188
rect 13836 -75232 13880 -75188
rect 13936 -75232 13980 -75188
rect 14036 -75232 14080 -75188
rect 14136 -75232 14180 -75188
rect 14236 -75232 14280 -75188
rect 14336 -75232 14380 -75188
rect 14436 -75232 14480 -75188
rect 14536 -75232 14580 -75188
rect 14636 -75232 14680 -75188
rect 14736 -75232 14780 -75188
rect 15236 -75232 15280 -75188
rect 15336 -75232 15380 -75188
rect 15436 -75232 15480 -75188
rect 15536 -75232 15580 -75188
rect 15636 -75232 15680 -75188
rect 15736 -75232 15780 -75188
rect 15836 -75232 15880 -75188
rect 15936 -75232 15980 -75188
rect 16036 -75232 16080 -75188
rect 16136 -75232 16180 -75188
rect 16236 -75232 16280 -75188
rect 16336 -75232 16380 -75188
rect 16436 -75232 16480 -75188
rect 16536 -75232 16580 -75188
rect 16636 -75232 16680 -75188
rect 16736 -75232 16780 -75188
rect 9236 -75332 9280 -75288
rect 9336 -75332 9380 -75288
rect 9436 -75332 9480 -75288
rect 9536 -75332 9580 -75288
rect 9636 -75332 9680 -75288
rect 9736 -75332 9780 -75288
rect 9836 -75332 9880 -75288
rect 9936 -75332 9980 -75288
rect 10036 -75332 10080 -75288
rect 10136 -75332 10180 -75288
rect 10236 -75332 10280 -75288
rect 10336 -75332 10380 -75288
rect 10436 -75332 10480 -75288
rect 10536 -75332 10580 -75288
rect 10636 -75332 10680 -75288
rect 10736 -75332 10780 -75288
rect 11236 -75332 11280 -75288
rect 11336 -75332 11380 -75288
rect 11436 -75332 11480 -75288
rect 11536 -75332 11580 -75288
rect 11636 -75332 11680 -75288
rect 11736 -75332 11780 -75288
rect 11836 -75332 11880 -75288
rect 11936 -75332 11980 -75288
rect 12036 -75332 12080 -75288
rect 12136 -75332 12180 -75288
rect 12236 -75332 12280 -75288
rect 12336 -75332 12380 -75288
rect 12436 -75332 12480 -75288
rect 12536 -75332 12580 -75288
rect 12636 -75332 12680 -75288
rect 12736 -75332 12780 -75288
rect 13236 -75332 13280 -75288
rect 13336 -75332 13380 -75288
rect 13436 -75332 13480 -75288
rect 13536 -75332 13580 -75288
rect 13636 -75332 13680 -75288
rect 13736 -75332 13780 -75288
rect 13836 -75332 13880 -75288
rect 13936 -75332 13980 -75288
rect 14036 -75332 14080 -75288
rect 14136 -75332 14180 -75288
rect 14236 -75332 14280 -75288
rect 14336 -75332 14380 -75288
rect 14436 -75332 14480 -75288
rect 14536 -75332 14580 -75288
rect 14636 -75332 14680 -75288
rect 14736 -75332 14780 -75288
rect 15236 -75332 15280 -75288
rect 15336 -75332 15380 -75288
rect 15436 -75332 15480 -75288
rect 15536 -75332 15580 -75288
rect 15636 -75332 15680 -75288
rect 15736 -75332 15780 -75288
rect 15836 -75332 15880 -75288
rect 15936 -75332 15980 -75288
rect 16036 -75332 16080 -75288
rect 16136 -75332 16180 -75288
rect 16236 -75332 16280 -75288
rect 16336 -75332 16380 -75288
rect 16436 -75332 16480 -75288
rect 16536 -75332 16580 -75288
rect 16636 -75332 16680 -75288
rect 16736 -75332 16780 -75288
rect 9236 -75432 9280 -75388
rect 9336 -75432 9380 -75388
rect 9436 -75432 9480 -75388
rect 9536 -75432 9580 -75388
rect 9636 -75432 9680 -75388
rect 9736 -75432 9780 -75388
rect 9836 -75432 9880 -75388
rect 9936 -75432 9980 -75388
rect 10036 -75432 10080 -75388
rect 10136 -75432 10180 -75388
rect 10236 -75432 10280 -75388
rect 10336 -75432 10380 -75388
rect 10436 -75432 10480 -75388
rect 10536 -75432 10580 -75388
rect 10636 -75432 10680 -75388
rect 10736 -75432 10780 -75388
rect 11236 -75432 11280 -75388
rect 11336 -75432 11380 -75388
rect 11436 -75432 11480 -75388
rect 11536 -75432 11580 -75388
rect 11636 -75432 11680 -75388
rect 11736 -75432 11780 -75388
rect 11836 -75432 11880 -75388
rect 11936 -75432 11980 -75388
rect 12036 -75432 12080 -75388
rect 12136 -75432 12180 -75388
rect 12236 -75432 12280 -75388
rect 12336 -75432 12380 -75388
rect 12436 -75432 12480 -75388
rect 12536 -75432 12580 -75388
rect 12636 -75432 12680 -75388
rect 12736 -75432 12780 -75388
rect 13236 -75432 13280 -75388
rect 13336 -75432 13380 -75388
rect 13436 -75432 13480 -75388
rect 13536 -75432 13580 -75388
rect 13636 -75432 13680 -75388
rect 13736 -75432 13780 -75388
rect 13836 -75432 13880 -75388
rect 13936 -75432 13980 -75388
rect 14036 -75432 14080 -75388
rect 14136 -75432 14180 -75388
rect 14236 -75432 14280 -75388
rect 14336 -75432 14380 -75388
rect 14436 -75432 14480 -75388
rect 14536 -75432 14580 -75388
rect 14636 -75432 14680 -75388
rect 14736 -75432 14780 -75388
rect 15236 -75432 15280 -75388
rect 15336 -75432 15380 -75388
rect 15436 -75432 15480 -75388
rect 15536 -75432 15580 -75388
rect 15636 -75432 15680 -75388
rect 15736 -75432 15780 -75388
rect 15836 -75432 15880 -75388
rect 15936 -75432 15980 -75388
rect 16036 -75432 16080 -75388
rect 16136 -75432 16180 -75388
rect 16236 -75432 16280 -75388
rect 16336 -75432 16380 -75388
rect 16436 -75432 16480 -75388
rect 16536 -75432 16580 -75388
rect 16636 -75432 16680 -75388
rect 16736 -75432 16780 -75388
rect 9236 -75532 9280 -75488
rect 9336 -75532 9380 -75488
rect 9436 -75532 9480 -75488
rect 9536 -75532 9580 -75488
rect 9636 -75532 9680 -75488
rect 9736 -75532 9780 -75488
rect 9836 -75532 9880 -75488
rect 9936 -75532 9980 -75488
rect 10036 -75532 10080 -75488
rect 10136 -75532 10180 -75488
rect 10236 -75532 10280 -75488
rect 10336 -75532 10380 -75488
rect 10436 -75532 10480 -75488
rect 10536 -75532 10580 -75488
rect 10636 -75532 10680 -75488
rect 10736 -75532 10780 -75488
rect 11236 -75532 11280 -75488
rect 11336 -75532 11380 -75488
rect 11436 -75532 11480 -75488
rect 11536 -75532 11580 -75488
rect 11636 -75532 11680 -75488
rect 11736 -75532 11780 -75488
rect 11836 -75532 11880 -75488
rect 11936 -75532 11980 -75488
rect 12036 -75532 12080 -75488
rect 12136 -75532 12180 -75488
rect 12236 -75532 12280 -75488
rect 12336 -75532 12380 -75488
rect 12436 -75532 12480 -75488
rect 12536 -75532 12580 -75488
rect 12636 -75532 12680 -75488
rect 12736 -75532 12780 -75488
rect 13236 -75532 13280 -75488
rect 13336 -75532 13380 -75488
rect 13436 -75532 13480 -75488
rect 13536 -75532 13580 -75488
rect 13636 -75532 13680 -75488
rect 13736 -75532 13780 -75488
rect 13836 -75532 13880 -75488
rect 13936 -75532 13980 -75488
rect 14036 -75532 14080 -75488
rect 14136 -75532 14180 -75488
rect 14236 -75532 14280 -75488
rect 14336 -75532 14380 -75488
rect 14436 -75532 14480 -75488
rect 14536 -75532 14580 -75488
rect 14636 -75532 14680 -75488
rect 14736 -75532 14780 -75488
rect 15236 -75532 15280 -75488
rect 15336 -75532 15380 -75488
rect 15436 -75532 15480 -75488
rect 15536 -75532 15580 -75488
rect 15636 -75532 15680 -75488
rect 15736 -75532 15780 -75488
rect 15836 -75532 15880 -75488
rect 15936 -75532 15980 -75488
rect 16036 -75532 16080 -75488
rect 16136 -75532 16180 -75488
rect 16236 -75532 16280 -75488
rect 16336 -75532 16380 -75488
rect 16436 -75532 16480 -75488
rect 16536 -75532 16580 -75488
rect 16636 -75532 16680 -75488
rect 16736 -75532 16780 -75488
rect 9236 -75632 9280 -75588
rect 9336 -75632 9380 -75588
rect 9436 -75632 9480 -75588
rect 9536 -75632 9580 -75588
rect 9636 -75632 9680 -75588
rect 9736 -75632 9780 -75588
rect 9836 -75632 9880 -75588
rect 9936 -75632 9980 -75588
rect 10036 -75632 10080 -75588
rect 10136 -75632 10180 -75588
rect 10236 -75632 10280 -75588
rect 10336 -75632 10380 -75588
rect 10436 -75632 10480 -75588
rect 10536 -75632 10580 -75588
rect 10636 -75632 10680 -75588
rect 10736 -75632 10780 -75588
rect 11236 -75632 11280 -75588
rect 11336 -75632 11380 -75588
rect 11436 -75632 11480 -75588
rect 11536 -75632 11580 -75588
rect 11636 -75632 11680 -75588
rect 11736 -75632 11780 -75588
rect 11836 -75632 11880 -75588
rect 11936 -75632 11980 -75588
rect 12036 -75632 12080 -75588
rect 12136 -75632 12180 -75588
rect 12236 -75632 12280 -75588
rect 12336 -75632 12380 -75588
rect 12436 -75632 12480 -75588
rect 12536 -75632 12580 -75588
rect 12636 -75632 12680 -75588
rect 12736 -75632 12780 -75588
rect 13236 -75632 13280 -75588
rect 13336 -75632 13380 -75588
rect 13436 -75632 13480 -75588
rect 13536 -75632 13580 -75588
rect 13636 -75632 13680 -75588
rect 13736 -75632 13780 -75588
rect 13836 -75632 13880 -75588
rect 13936 -75632 13980 -75588
rect 14036 -75632 14080 -75588
rect 14136 -75632 14180 -75588
rect 14236 -75632 14280 -75588
rect 14336 -75632 14380 -75588
rect 14436 -75632 14480 -75588
rect 14536 -75632 14580 -75588
rect 14636 -75632 14680 -75588
rect 14736 -75632 14780 -75588
rect 15236 -75632 15280 -75588
rect 15336 -75632 15380 -75588
rect 15436 -75632 15480 -75588
rect 15536 -75632 15580 -75588
rect 15636 -75632 15680 -75588
rect 15736 -75632 15780 -75588
rect 15836 -75632 15880 -75588
rect 15936 -75632 15980 -75588
rect 16036 -75632 16080 -75588
rect 16136 -75632 16180 -75588
rect 16236 -75632 16280 -75588
rect 16336 -75632 16380 -75588
rect 16436 -75632 16480 -75588
rect 16536 -75632 16580 -75588
rect 16636 -75632 16680 -75588
rect 16736 -75632 16780 -75588
rect 9236 -75732 9280 -75688
rect 9336 -75732 9380 -75688
rect 9436 -75732 9480 -75688
rect 9536 -75732 9580 -75688
rect 9636 -75732 9680 -75688
rect 9736 -75732 9780 -75688
rect 9836 -75732 9880 -75688
rect 9936 -75732 9980 -75688
rect 10036 -75732 10080 -75688
rect 10136 -75732 10180 -75688
rect 10236 -75732 10280 -75688
rect 10336 -75732 10380 -75688
rect 10436 -75732 10480 -75688
rect 10536 -75732 10580 -75688
rect 10636 -75732 10680 -75688
rect 10736 -75732 10780 -75688
rect 11236 -75732 11280 -75688
rect 11336 -75732 11380 -75688
rect 11436 -75732 11480 -75688
rect 11536 -75732 11580 -75688
rect 11636 -75732 11680 -75688
rect 11736 -75732 11780 -75688
rect 11836 -75732 11880 -75688
rect 11936 -75732 11980 -75688
rect 12036 -75732 12080 -75688
rect 12136 -75732 12180 -75688
rect 12236 -75732 12280 -75688
rect 12336 -75732 12380 -75688
rect 12436 -75732 12480 -75688
rect 12536 -75732 12580 -75688
rect 12636 -75732 12680 -75688
rect 12736 -75732 12780 -75688
rect 13236 -75732 13280 -75688
rect 13336 -75732 13380 -75688
rect 13436 -75732 13480 -75688
rect 13536 -75732 13580 -75688
rect 13636 -75732 13680 -75688
rect 13736 -75732 13780 -75688
rect 13836 -75732 13880 -75688
rect 13936 -75732 13980 -75688
rect 14036 -75732 14080 -75688
rect 14136 -75732 14180 -75688
rect 14236 -75732 14280 -75688
rect 14336 -75732 14380 -75688
rect 14436 -75732 14480 -75688
rect 14536 -75732 14580 -75688
rect 14636 -75732 14680 -75688
rect 14736 -75732 14780 -75688
rect 15236 -75732 15280 -75688
rect 15336 -75732 15380 -75688
rect 15436 -75732 15480 -75688
rect 15536 -75732 15580 -75688
rect 15636 -75732 15680 -75688
rect 15736 -75732 15780 -75688
rect 15836 -75732 15880 -75688
rect 15936 -75732 15980 -75688
rect 16036 -75732 16080 -75688
rect 16136 -75732 16180 -75688
rect 16236 -75732 16280 -75688
rect 16336 -75732 16380 -75688
rect 16436 -75732 16480 -75688
rect 16536 -75732 16580 -75688
rect 16636 -75732 16680 -75688
rect 16736 -75732 16780 -75688
rect 9236 -75832 9280 -75788
rect 9336 -75832 9380 -75788
rect 9436 -75832 9480 -75788
rect 9536 -75832 9580 -75788
rect 9636 -75832 9680 -75788
rect 9736 -75832 9780 -75788
rect 9836 -75832 9880 -75788
rect 9936 -75832 9980 -75788
rect 10036 -75832 10080 -75788
rect 10136 -75832 10180 -75788
rect 10236 -75832 10280 -75788
rect 10336 -75832 10380 -75788
rect 10436 -75832 10480 -75788
rect 10536 -75832 10580 -75788
rect 10636 -75832 10680 -75788
rect 10736 -75832 10780 -75788
rect 11236 -75832 11280 -75788
rect 11336 -75832 11380 -75788
rect 11436 -75832 11480 -75788
rect 11536 -75832 11580 -75788
rect 11636 -75832 11680 -75788
rect 11736 -75832 11780 -75788
rect 11836 -75832 11880 -75788
rect 11936 -75832 11980 -75788
rect 12036 -75832 12080 -75788
rect 12136 -75832 12180 -75788
rect 12236 -75832 12280 -75788
rect 12336 -75832 12380 -75788
rect 12436 -75832 12480 -75788
rect 12536 -75832 12580 -75788
rect 12636 -75832 12680 -75788
rect 12736 -75832 12780 -75788
rect 13236 -75832 13280 -75788
rect 13336 -75832 13380 -75788
rect 13436 -75832 13480 -75788
rect 13536 -75832 13580 -75788
rect 13636 -75832 13680 -75788
rect 13736 -75832 13780 -75788
rect 13836 -75832 13880 -75788
rect 13936 -75832 13980 -75788
rect 14036 -75832 14080 -75788
rect 14136 -75832 14180 -75788
rect 14236 -75832 14280 -75788
rect 14336 -75832 14380 -75788
rect 14436 -75832 14480 -75788
rect 14536 -75832 14580 -75788
rect 14636 -75832 14680 -75788
rect 14736 -75832 14780 -75788
rect 15236 -75832 15280 -75788
rect 15336 -75832 15380 -75788
rect 15436 -75832 15480 -75788
rect 15536 -75832 15580 -75788
rect 15636 -75832 15680 -75788
rect 15736 -75832 15780 -75788
rect 15836 -75832 15880 -75788
rect 15936 -75832 15980 -75788
rect 16036 -75832 16080 -75788
rect 16136 -75832 16180 -75788
rect 16236 -75832 16280 -75788
rect 16336 -75832 16380 -75788
rect 16436 -75832 16480 -75788
rect 16536 -75832 16580 -75788
rect 16636 -75832 16680 -75788
rect 16736 -75832 16780 -75788
rect 9236 -75932 9280 -75888
rect 9336 -75932 9380 -75888
rect 9436 -75932 9480 -75888
rect 9536 -75932 9580 -75888
rect 9636 -75932 9680 -75888
rect 9736 -75932 9780 -75888
rect 9836 -75932 9880 -75888
rect 9936 -75932 9980 -75888
rect 10036 -75932 10080 -75888
rect 10136 -75932 10180 -75888
rect 10236 -75932 10280 -75888
rect 10336 -75932 10380 -75888
rect 10436 -75932 10480 -75888
rect 10536 -75932 10580 -75888
rect 10636 -75932 10680 -75888
rect 10736 -75932 10780 -75888
rect 11236 -75932 11280 -75888
rect 11336 -75932 11380 -75888
rect 11436 -75932 11480 -75888
rect 11536 -75932 11580 -75888
rect 11636 -75932 11680 -75888
rect 11736 -75932 11780 -75888
rect 11836 -75932 11880 -75888
rect 11936 -75932 11980 -75888
rect 12036 -75932 12080 -75888
rect 12136 -75932 12180 -75888
rect 12236 -75932 12280 -75888
rect 12336 -75932 12380 -75888
rect 12436 -75932 12480 -75888
rect 12536 -75932 12580 -75888
rect 12636 -75932 12680 -75888
rect 12736 -75932 12780 -75888
rect 13236 -75932 13280 -75888
rect 13336 -75932 13380 -75888
rect 13436 -75932 13480 -75888
rect 13536 -75932 13580 -75888
rect 13636 -75932 13680 -75888
rect 13736 -75932 13780 -75888
rect 13836 -75932 13880 -75888
rect 13936 -75932 13980 -75888
rect 14036 -75932 14080 -75888
rect 14136 -75932 14180 -75888
rect 14236 -75932 14280 -75888
rect 14336 -75932 14380 -75888
rect 14436 -75932 14480 -75888
rect 14536 -75932 14580 -75888
rect 14636 -75932 14680 -75888
rect 14736 -75932 14780 -75888
rect 15236 -75932 15280 -75888
rect 15336 -75932 15380 -75888
rect 15436 -75932 15480 -75888
rect 15536 -75932 15580 -75888
rect 15636 -75932 15680 -75888
rect 15736 -75932 15780 -75888
rect 15836 -75932 15880 -75888
rect 15936 -75932 15980 -75888
rect 16036 -75932 16080 -75888
rect 16136 -75932 16180 -75888
rect 16236 -75932 16280 -75888
rect 16336 -75932 16380 -75888
rect 16436 -75932 16480 -75888
rect 16536 -75932 16580 -75888
rect 16636 -75932 16680 -75888
rect 16736 -75932 16780 -75888
rect 9236 -76032 9280 -75988
rect 9336 -76032 9380 -75988
rect 9436 -76032 9480 -75988
rect 9536 -76032 9580 -75988
rect 9636 -76032 9680 -75988
rect 9736 -76032 9780 -75988
rect 9836 -76032 9880 -75988
rect 9936 -76032 9980 -75988
rect 10036 -76032 10080 -75988
rect 10136 -76032 10180 -75988
rect 10236 -76032 10280 -75988
rect 10336 -76032 10380 -75988
rect 10436 -76032 10480 -75988
rect 10536 -76032 10580 -75988
rect 10636 -76032 10680 -75988
rect 10736 -76032 10780 -75988
rect 11236 -76032 11280 -75988
rect 11336 -76032 11380 -75988
rect 11436 -76032 11480 -75988
rect 11536 -76032 11580 -75988
rect 11636 -76032 11680 -75988
rect 11736 -76032 11780 -75988
rect 11836 -76032 11880 -75988
rect 11936 -76032 11980 -75988
rect 12036 -76032 12080 -75988
rect 12136 -76032 12180 -75988
rect 12236 -76032 12280 -75988
rect 12336 -76032 12380 -75988
rect 12436 -76032 12480 -75988
rect 12536 -76032 12580 -75988
rect 12636 -76032 12680 -75988
rect 12736 -76032 12780 -75988
rect 13236 -76032 13280 -75988
rect 13336 -76032 13380 -75988
rect 13436 -76032 13480 -75988
rect 13536 -76032 13580 -75988
rect 13636 -76032 13680 -75988
rect 13736 -76032 13780 -75988
rect 13836 -76032 13880 -75988
rect 13936 -76032 13980 -75988
rect 14036 -76032 14080 -75988
rect 14136 -76032 14180 -75988
rect 14236 -76032 14280 -75988
rect 14336 -76032 14380 -75988
rect 14436 -76032 14480 -75988
rect 14536 -76032 14580 -75988
rect 14636 -76032 14680 -75988
rect 14736 -76032 14780 -75988
rect 15236 -76032 15280 -75988
rect 15336 -76032 15380 -75988
rect 15436 -76032 15480 -75988
rect 15536 -76032 15580 -75988
rect 15636 -76032 15680 -75988
rect 15736 -76032 15780 -75988
rect 15836 -76032 15880 -75988
rect 15936 -76032 15980 -75988
rect 16036 -76032 16080 -75988
rect 16136 -76032 16180 -75988
rect 16236 -76032 16280 -75988
rect 16336 -76032 16380 -75988
rect 16436 -76032 16480 -75988
rect 16536 -76032 16580 -75988
rect 16636 -76032 16680 -75988
rect 16736 -76032 16780 -75988
rect 9236 -76132 9280 -76088
rect 9336 -76132 9380 -76088
rect 9436 -76132 9480 -76088
rect 9536 -76132 9580 -76088
rect 9636 -76132 9680 -76088
rect 9736 -76132 9780 -76088
rect 9836 -76132 9880 -76088
rect 9936 -76132 9980 -76088
rect 10036 -76132 10080 -76088
rect 10136 -76132 10180 -76088
rect 10236 -76132 10280 -76088
rect 10336 -76132 10380 -76088
rect 10436 -76132 10480 -76088
rect 10536 -76132 10580 -76088
rect 10636 -76132 10680 -76088
rect 10736 -76132 10780 -76088
rect 11236 -76132 11280 -76088
rect 11336 -76132 11380 -76088
rect 11436 -76132 11480 -76088
rect 11536 -76132 11580 -76088
rect 11636 -76132 11680 -76088
rect 11736 -76132 11780 -76088
rect 11836 -76132 11880 -76088
rect 11936 -76132 11980 -76088
rect 12036 -76132 12080 -76088
rect 12136 -76132 12180 -76088
rect 12236 -76132 12280 -76088
rect 12336 -76132 12380 -76088
rect 12436 -76132 12480 -76088
rect 12536 -76132 12580 -76088
rect 12636 -76132 12680 -76088
rect 12736 -76132 12780 -76088
rect 13236 -76132 13280 -76088
rect 13336 -76132 13380 -76088
rect 13436 -76132 13480 -76088
rect 13536 -76132 13580 -76088
rect 13636 -76132 13680 -76088
rect 13736 -76132 13780 -76088
rect 13836 -76132 13880 -76088
rect 13936 -76132 13980 -76088
rect 14036 -76132 14080 -76088
rect 14136 -76132 14180 -76088
rect 14236 -76132 14280 -76088
rect 14336 -76132 14380 -76088
rect 14436 -76132 14480 -76088
rect 14536 -76132 14580 -76088
rect 14636 -76132 14680 -76088
rect 14736 -76132 14780 -76088
rect 15236 -76132 15280 -76088
rect 15336 -76132 15380 -76088
rect 15436 -76132 15480 -76088
rect 15536 -76132 15580 -76088
rect 15636 -76132 15680 -76088
rect 15736 -76132 15780 -76088
rect 15836 -76132 15880 -76088
rect 15936 -76132 15980 -76088
rect 16036 -76132 16080 -76088
rect 16136 -76132 16180 -76088
rect 16236 -76132 16280 -76088
rect 16336 -76132 16380 -76088
rect 16436 -76132 16480 -76088
rect 16536 -76132 16580 -76088
rect 16636 -76132 16680 -76088
rect 16736 -76132 16780 -76088
rect 9236 -76232 9280 -76188
rect 9336 -76232 9380 -76188
rect 9436 -76232 9480 -76188
rect 9536 -76232 9580 -76188
rect 9636 -76232 9680 -76188
rect 9736 -76232 9780 -76188
rect 9836 -76232 9880 -76188
rect 9936 -76232 9980 -76188
rect 10036 -76232 10080 -76188
rect 10136 -76232 10180 -76188
rect 10236 -76232 10280 -76188
rect 10336 -76232 10380 -76188
rect 10436 -76232 10480 -76188
rect 10536 -76232 10580 -76188
rect 10636 -76232 10680 -76188
rect 10736 -76232 10780 -76188
rect 11236 -76232 11280 -76188
rect 11336 -76232 11380 -76188
rect 11436 -76232 11480 -76188
rect 11536 -76232 11580 -76188
rect 11636 -76232 11680 -76188
rect 11736 -76232 11780 -76188
rect 11836 -76232 11880 -76188
rect 11936 -76232 11980 -76188
rect 12036 -76232 12080 -76188
rect 12136 -76232 12180 -76188
rect 12236 -76232 12280 -76188
rect 12336 -76232 12380 -76188
rect 12436 -76232 12480 -76188
rect 12536 -76232 12580 -76188
rect 12636 -76232 12680 -76188
rect 12736 -76232 12780 -76188
rect 13236 -76232 13280 -76188
rect 13336 -76232 13380 -76188
rect 13436 -76232 13480 -76188
rect 13536 -76232 13580 -76188
rect 13636 -76232 13680 -76188
rect 13736 -76232 13780 -76188
rect 13836 -76232 13880 -76188
rect 13936 -76232 13980 -76188
rect 14036 -76232 14080 -76188
rect 14136 -76232 14180 -76188
rect 14236 -76232 14280 -76188
rect 14336 -76232 14380 -76188
rect 14436 -76232 14480 -76188
rect 14536 -76232 14580 -76188
rect 14636 -76232 14680 -76188
rect 14736 -76232 14780 -76188
rect 15236 -76232 15280 -76188
rect 15336 -76232 15380 -76188
rect 15436 -76232 15480 -76188
rect 15536 -76232 15580 -76188
rect 15636 -76232 15680 -76188
rect 15736 -76232 15780 -76188
rect 15836 -76232 15880 -76188
rect 15936 -76232 15980 -76188
rect 16036 -76232 16080 -76188
rect 16136 -76232 16180 -76188
rect 16236 -76232 16280 -76188
rect 16336 -76232 16380 -76188
rect 16436 -76232 16480 -76188
rect 16536 -76232 16580 -76188
rect 16636 -76232 16680 -76188
rect 16736 -76232 16780 -76188
rect 9236 -76332 9280 -76288
rect 9336 -76332 9380 -76288
rect 9436 -76332 9480 -76288
rect 9536 -76332 9580 -76288
rect 9636 -76332 9680 -76288
rect 9736 -76332 9780 -76288
rect 9836 -76332 9880 -76288
rect 9936 -76332 9980 -76288
rect 10036 -76332 10080 -76288
rect 10136 -76332 10180 -76288
rect 10236 -76332 10280 -76288
rect 10336 -76332 10380 -76288
rect 10436 -76332 10480 -76288
rect 10536 -76332 10580 -76288
rect 10636 -76332 10680 -76288
rect 10736 -76332 10780 -76288
rect 11236 -76332 11280 -76288
rect 11336 -76332 11380 -76288
rect 11436 -76332 11480 -76288
rect 11536 -76332 11580 -76288
rect 11636 -76332 11680 -76288
rect 11736 -76332 11780 -76288
rect 11836 -76332 11880 -76288
rect 11936 -76332 11980 -76288
rect 12036 -76332 12080 -76288
rect 12136 -76332 12180 -76288
rect 12236 -76332 12280 -76288
rect 12336 -76332 12380 -76288
rect 12436 -76332 12480 -76288
rect 12536 -76332 12580 -76288
rect 12636 -76332 12680 -76288
rect 12736 -76332 12780 -76288
rect 13236 -76332 13280 -76288
rect 13336 -76332 13380 -76288
rect 13436 -76332 13480 -76288
rect 13536 -76332 13580 -76288
rect 13636 -76332 13680 -76288
rect 13736 -76332 13780 -76288
rect 13836 -76332 13880 -76288
rect 13936 -76332 13980 -76288
rect 14036 -76332 14080 -76288
rect 14136 -76332 14180 -76288
rect 14236 -76332 14280 -76288
rect 14336 -76332 14380 -76288
rect 14436 -76332 14480 -76288
rect 14536 -76332 14580 -76288
rect 14636 -76332 14680 -76288
rect 14736 -76332 14780 -76288
rect 15236 -76332 15280 -76288
rect 15336 -76332 15380 -76288
rect 15436 -76332 15480 -76288
rect 15536 -76332 15580 -76288
rect 15636 -76332 15680 -76288
rect 15736 -76332 15780 -76288
rect 15836 -76332 15880 -76288
rect 15936 -76332 15980 -76288
rect 16036 -76332 16080 -76288
rect 16136 -76332 16180 -76288
rect 16236 -76332 16280 -76288
rect 16336 -76332 16380 -76288
rect 16436 -76332 16480 -76288
rect 16536 -76332 16580 -76288
rect 16636 -76332 16680 -76288
rect 16736 -76332 16780 -76288
rect 9236 -76432 9280 -76388
rect 9336 -76432 9380 -76388
rect 9436 -76432 9480 -76388
rect 9536 -76432 9580 -76388
rect 9636 -76432 9680 -76388
rect 9736 -76432 9780 -76388
rect 9836 -76432 9880 -76388
rect 9936 -76432 9980 -76388
rect 10036 -76432 10080 -76388
rect 10136 -76432 10180 -76388
rect 10236 -76432 10280 -76388
rect 10336 -76432 10380 -76388
rect 10436 -76432 10480 -76388
rect 10536 -76432 10580 -76388
rect 10636 -76432 10680 -76388
rect 10736 -76432 10780 -76388
rect 11236 -76432 11280 -76388
rect 11336 -76432 11380 -76388
rect 11436 -76432 11480 -76388
rect 11536 -76432 11580 -76388
rect 11636 -76432 11680 -76388
rect 11736 -76432 11780 -76388
rect 11836 -76432 11880 -76388
rect 11936 -76432 11980 -76388
rect 12036 -76432 12080 -76388
rect 12136 -76432 12180 -76388
rect 12236 -76432 12280 -76388
rect 12336 -76432 12380 -76388
rect 12436 -76432 12480 -76388
rect 12536 -76432 12580 -76388
rect 12636 -76432 12680 -76388
rect 12736 -76432 12780 -76388
rect 13236 -76432 13280 -76388
rect 13336 -76432 13380 -76388
rect 13436 -76432 13480 -76388
rect 13536 -76432 13580 -76388
rect 13636 -76432 13680 -76388
rect 13736 -76432 13780 -76388
rect 13836 -76432 13880 -76388
rect 13936 -76432 13980 -76388
rect 14036 -76432 14080 -76388
rect 14136 -76432 14180 -76388
rect 14236 -76432 14280 -76388
rect 14336 -76432 14380 -76388
rect 14436 -76432 14480 -76388
rect 14536 -76432 14580 -76388
rect 14636 -76432 14680 -76388
rect 14736 -76432 14780 -76388
rect 15236 -76432 15280 -76388
rect 15336 -76432 15380 -76388
rect 15436 -76432 15480 -76388
rect 15536 -76432 15580 -76388
rect 15636 -76432 15680 -76388
rect 15736 -76432 15780 -76388
rect 15836 -76432 15880 -76388
rect 15936 -76432 15980 -76388
rect 16036 -76432 16080 -76388
rect 16136 -76432 16180 -76388
rect 16236 -76432 16280 -76388
rect 16336 -76432 16380 -76388
rect 16436 -76432 16480 -76388
rect 16536 -76432 16580 -76388
rect 16636 -76432 16680 -76388
rect 16736 -76432 16780 -76388
rect 9236 -76532 9280 -76488
rect 9336 -76532 9380 -76488
rect 9436 -76532 9480 -76488
rect 9536 -76532 9580 -76488
rect 9636 -76532 9680 -76488
rect 9736 -76532 9780 -76488
rect 9836 -76532 9880 -76488
rect 9936 -76532 9980 -76488
rect 10036 -76532 10080 -76488
rect 10136 -76532 10180 -76488
rect 10236 -76532 10280 -76488
rect 10336 -76532 10380 -76488
rect 10436 -76532 10480 -76488
rect 10536 -76532 10580 -76488
rect 10636 -76532 10680 -76488
rect 10736 -76532 10780 -76488
rect 11236 -76532 11280 -76488
rect 11336 -76532 11380 -76488
rect 11436 -76532 11480 -76488
rect 11536 -76532 11580 -76488
rect 11636 -76532 11680 -76488
rect 11736 -76532 11780 -76488
rect 11836 -76532 11880 -76488
rect 11936 -76532 11980 -76488
rect 12036 -76532 12080 -76488
rect 12136 -76532 12180 -76488
rect 12236 -76532 12280 -76488
rect 12336 -76532 12380 -76488
rect 12436 -76532 12480 -76488
rect 12536 -76532 12580 -76488
rect 12636 -76532 12680 -76488
rect 12736 -76532 12780 -76488
rect 13236 -76532 13280 -76488
rect 13336 -76532 13380 -76488
rect 13436 -76532 13480 -76488
rect 13536 -76532 13580 -76488
rect 13636 -76532 13680 -76488
rect 13736 -76532 13780 -76488
rect 13836 -76532 13880 -76488
rect 13936 -76532 13980 -76488
rect 14036 -76532 14080 -76488
rect 14136 -76532 14180 -76488
rect 14236 -76532 14280 -76488
rect 14336 -76532 14380 -76488
rect 14436 -76532 14480 -76488
rect 14536 -76532 14580 -76488
rect 14636 -76532 14680 -76488
rect 14736 -76532 14780 -76488
rect 15236 -76532 15280 -76488
rect 15336 -76532 15380 -76488
rect 15436 -76532 15480 -76488
rect 15536 -76532 15580 -76488
rect 15636 -76532 15680 -76488
rect 15736 -76532 15780 -76488
rect 15836 -76532 15880 -76488
rect 15936 -76532 15980 -76488
rect 16036 -76532 16080 -76488
rect 16136 -76532 16180 -76488
rect 16236 -76532 16280 -76488
rect 16336 -76532 16380 -76488
rect 16436 -76532 16480 -76488
rect 16536 -76532 16580 -76488
rect 16636 -76532 16680 -76488
rect 16736 -76532 16780 -76488
rect 9236 -76632 9280 -76588
rect 9336 -76632 9380 -76588
rect 9436 -76632 9480 -76588
rect 9536 -76632 9580 -76588
rect 9636 -76632 9680 -76588
rect 9736 -76632 9780 -76588
rect 9836 -76632 9880 -76588
rect 9936 -76632 9980 -76588
rect 10036 -76632 10080 -76588
rect 10136 -76632 10180 -76588
rect 10236 -76632 10280 -76588
rect 10336 -76632 10380 -76588
rect 10436 -76632 10480 -76588
rect 10536 -76632 10580 -76588
rect 10636 -76632 10680 -76588
rect 10736 -76632 10780 -76588
rect 11236 -76632 11280 -76588
rect 11336 -76632 11380 -76588
rect 11436 -76632 11480 -76588
rect 11536 -76632 11580 -76588
rect 11636 -76632 11680 -76588
rect 11736 -76632 11780 -76588
rect 11836 -76632 11880 -76588
rect 11936 -76632 11980 -76588
rect 12036 -76632 12080 -76588
rect 12136 -76632 12180 -76588
rect 12236 -76632 12280 -76588
rect 12336 -76632 12380 -76588
rect 12436 -76632 12480 -76588
rect 12536 -76632 12580 -76588
rect 12636 -76632 12680 -76588
rect 12736 -76632 12780 -76588
rect 13236 -76632 13280 -76588
rect 13336 -76632 13380 -76588
rect 13436 -76632 13480 -76588
rect 13536 -76632 13580 -76588
rect 13636 -76632 13680 -76588
rect 13736 -76632 13780 -76588
rect 13836 -76632 13880 -76588
rect 13936 -76632 13980 -76588
rect 14036 -76632 14080 -76588
rect 14136 -76632 14180 -76588
rect 14236 -76632 14280 -76588
rect 14336 -76632 14380 -76588
rect 14436 -76632 14480 -76588
rect 14536 -76632 14580 -76588
rect 14636 -76632 14680 -76588
rect 14736 -76632 14780 -76588
rect 15236 -76632 15280 -76588
rect 15336 -76632 15380 -76588
rect 15436 -76632 15480 -76588
rect 15536 -76632 15580 -76588
rect 15636 -76632 15680 -76588
rect 15736 -76632 15780 -76588
rect 15836 -76632 15880 -76588
rect 15936 -76632 15980 -76588
rect 16036 -76632 16080 -76588
rect 16136 -76632 16180 -76588
rect 16236 -76632 16280 -76588
rect 16336 -76632 16380 -76588
rect 16436 -76632 16480 -76588
rect 16536 -76632 16580 -76588
rect 16636 -76632 16680 -76588
rect 16736 -76632 16780 -76588
rect 9236 -76732 9280 -76688
rect 9336 -76732 9380 -76688
rect 9436 -76732 9480 -76688
rect 9536 -76732 9580 -76688
rect 9636 -76732 9680 -76688
rect 9736 -76732 9780 -76688
rect 9836 -76732 9880 -76688
rect 9936 -76732 9980 -76688
rect 10036 -76732 10080 -76688
rect 10136 -76732 10180 -76688
rect 10236 -76732 10280 -76688
rect 10336 -76732 10380 -76688
rect 10436 -76732 10480 -76688
rect 10536 -76732 10580 -76688
rect 10636 -76732 10680 -76688
rect 10736 -76732 10780 -76688
rect 11236 -76732 11280 -76688
rect 11336 -76732 11380 -76688
rect 11436 -76732 11480 -76688
rect 11536 -76732 11580 -76688
rect 11636 -76732 11680 -76688
rect 11736 -76732 11780 -76688
rect 11836 -76732 11880 -76688
rect 11936 -76732 11980 -76688
rect 12036 -76732 12080 -76688
rect 12136 -76732 12180 -76688
rect 12236 -76732 12280 -76688
rect 12336 -76732 12380 -76688
rect 12436 -76732 12480 -76688
rect 12536 -76732 12580 -76688
rect 12636 -76732 12680 -76688
rect 12736 -76732 12780 -76688
rect 13236 -76732 13280 -76688
rect 13336 -76732 13380 -76688
rect 13436 -76732 13480 -76688
rect 13536 -76732 13580 -76688
rect 13636 -76732 13680 -76688
rect 13736 -76732 13780 -76688
rect 13836 -76732 13880 -76688
rect 13936 -76732 13980 -76688
rect 14036 -76732 14080 -76688
rect 14136 -76732 14180 -76688
rect 14236 -76732 14280 -76688
rect 14336 -76732 14380 -76688
rect 14436 -76732 14480 -76688
rect 14536 -76732 14580 -76688
rect 14636 -76732 14680 -76688
rect 14736 -76732 14780 -76688
rect 15236 -76732 15280 -76688
rect 15336 -76732 15380 -76688
rect 15436 -76732 15480 -76688
rect 15536 -76732 15580 -76688
rect 15636 -76732 15680 -76688
rect 15736 -76732 15780 -76688
rect 15836 -76732 15880 -76688
rect 15936 -76732 15980 -76688
rect 16036 -76732 16080 -76688
rect 16136 -76732 16180 -76688
rect 16236 -76732 16280 -76688
rect 16336 -76732 16380 -76688
rect 16436 -76732 16480 -76688
rect 16536 -76732 16580 -76688
rect 16636 -76732 16680 -76688
rect 16736 -76732 16780 -76688
rect -82968 -80503 -82924 -80459
rect -82868 -80503 -82824 -80459
rect -82768 -80503 -82724 -80459
rect -82668 -80503 -82624 -80459
rect -82568 -80503 -82524 -80459
rect -82468 -80503 -82424 -80459
rect -82368 -80503 -82324 -80459
rect -82268 -80503 -82224 -80459
rect -82168 -80503 -82124 -80459
rect -82068 -80503 -82024 -80459
rect -81968 -80503 -81924 -80459
rect -81868 -80503 -81824 -80459
rect -81768 -80503 -81724 -80459
rect -81668 -80503 -81624 -80459
rect -81568 -80503 -81524 -80459
rect -81468 -80503 -81424 -80459
rect -80968 -80503 -80924 -80459
rect -80868 -80503 -80824 -80459
rect -80768 -80503 -80724 -80459
rect -80668 -80503 -80624 -80459
rect -80568 -80503 -80524 -80459
rect -80468 -80503 -80424 -80459
rect -80368 -80503 -80324 -80459
rect -80268 -80503 -80224 -80459
rect -80168 -80503 -80124 -80459
rect -80068 -80503 -80024 -80459
rect -79968 -80503 -79924 -80459
rect -79868 -80503 -79824 -80459
rect -79768 -80503 -79724 -80459
rect -79668 -80503 -79624 -80459
rect -79568 -80503 -79524 -80459
rect -79468 -80503 -79424 -80459
rect -78968 -80503 -78924 -80459
rect -78868 -80503 -78824 -80459
rect -78768 -80503 -78724 -80459
rect -78668 -80503 -78624 -80459
rect -78568 -80503 -78524 -80459
rect -78468 -80503 -78424 -80459
rect -78368 -80503 -78324 -80459
rect -78268 -80503 -78224 -80459
rect -78168 -80503 -78124 -80459
rect -78068 -80503 -78024 -80459
rect -77968 -80503 -77924 -80459
rect -77868 -80503 -77824 -80459
rect -77768 -80503 -77724 -80459
rect -77668 -80503 -77624 -80459
rect -77568 -80503 -77524 -80459
rect -77468 -80503 -77424 -80459
rect -76968 -80503 -76924 -80459
rect -76868 -80503 -76824 -80459
rect -76768 -80503 -76724 -80459
rect -76668 -80503 -76624 -80459
rect -76568 -80503 -76524 -80459
rect -76468 -80503 -76424 -80459
rect -76368 -80503 -76324 -80459
rect -76268 -80503 -76224 -80459
rect -76168 -80503 -76124 -80459
rect -76068 -80503 -76024 -80459
rect -75968 -80503 -75924 -80459
rect -75868 -80503 -75824 -80459
rect -75768 -80503 -75724 -80459
rect -75668 -80503 -75624 -80459
rect -75568 -80503 -75524 -80459
rect -75468 -80503 -75424 -80459
rect -50017 -80505 -49973 -80461
rect -49917 -80505 -49873 -80461
rect -49817 -80505 -49773 -80461
rect -49717 -80505 -49673 -80461
rect -49617 -80505 -49573 -80461
rect -49517 -80505 -49473 -80461
rect -49417 -80505 -49373 -80461
rect -49317 -80505 -49273 -80461
rect -49217 -80505 -49173 -80461
rect -49117 -80505 -49073 -80461
rect -49017 -80505 -48973 -80461
rect -48917 -80505 -48873 -80461
rect -48817 -80505 -48773 -80461
rect -48717 -80505 -48673 -80461
rect -48617 -80505 -48573 -80461
rect -48517 -80505 -48473 -80461
rect -48017 -80505 -47973 -80461
rect -47917 -80505 -47873 -80461
rect -47817 -80505 -47773 -80461
rect -47717 -80505 -47673 -80461
rect -47617 -80505 -47573 -80461
rect -47517 -80505 -47473 -80461
rect -47417 -80505 -47373 -80461
rect -47317 -80505 -47273 -80461
rect -47217 -80505 -47173 -80461
rect -47117 -80505 -47073 -80461
rect -47017 -80505 -46973 -80461
rect -46917 -80505 -46873 -80461
rect -46817 -80505 -46773 -80461
rect -46717 -80505 -46673 -80461
rect -46617 -80505 -46573 -80461
rect -46517 -80505 -46473 -80461
rect -46017 -80505 -45973 -80461
rect -45917 -80505 -45873 -80461
rect -45817 -80505 -45773 -80461
rect -45717 -80505 -45673 -80461
rect -45617 -80505 -45573 -80461
rect -45517 -80505 -45473 -80461
rect -45417 -80505 -45373 -80461
rect -45317 -80505 -45273 -80461
rect -45217 -80505 -45173 -80461
rect -45117 -80505 -45073 -80461
rect -45017 -80505 -44973 -80461
rect -44917 -80505 -44873 -80461
rect -44817 -80505 -44773 -80461
rect -44717 -80505 -44673 -80461
rect -44617 -80505 -44573 -80461
rect -44517 -80505 -44473 -80461
rect -44017 -80505 -43973 -80461
rect -43917 -80505 -43873 -80461
rect -43817 -80505 -43773 -80461
rect -43717 -80505 -43673 -80461
rect -43617 -80505 -43573 -80461
rect -43517 -80505 -43473 -80461
rect -43417 -80505 -43373 -80461
rect -43317 -80505 -43273 -80461
rect -43217 -80505 -43173 -80461
rect -43117 -80505 -43073 -80461
rect -43017 -80505 -42973 -80461
rect -42917 -80505 -42873 -80461
rect -42817 -80505 -42773 -80461
rect -42717 -80505 -42673 -80461
rect -42617 -80505 -42573 -80461
rect -42517 -80505 -42473 -80461
rect 80737 -80499 80781 -80455
rect 80837 -80499 80881 -80455
rect 80937 -80499 80981 -80455
rect 81037 -80499 81081 -80455
rect 81137 -80499 81181 -80455
rect 81237 -80499 81281 -80455
rect 81337 -80499 81381 -80455
rect 81437 -80499 81481 -80455
rect 81537 -80499 81581 -80455
rect 81637 -80499 81681 -80455
rect 81737 -80499 81781 -80455
rect 81837 -80499 81881 -80455
rect 81937 -80499 81981 -80455
rect 82037 -80499 82081 -80455
rect 82137 -80499 82181 -80455
rect 82237 -80499 82281 -80455
rect 82737 -80499 82781 -80455
rect 82837 -80499 82881 -80455
rect 82937 -80499 82981 -80455
rect 83037 -80499 83081 -80455
rect 83137 -80499 83181 -80455
rect 83237 -80499 83281 -80455
rect 83337 -80499 83381 -80455
rect 83437 -80499 83481 -80455
rect 83537 -80499 83581 -80455
rect 83637 -80499 83681 -80455
rect 83737 -80499 83781 -80455
rect 83837 -80499 83881 -80455
rect 83937 -80499 83981 -80455
rect 84037 -80499 84081 -80455
rect 84137 -80499 84181 -80455
rect 84237 -80499 84281 -80455
rect 84737 -80499 84781 -80455
rect 84837 -80499 84881 -80455
rect 84937 -80499 84981 -80455
rect 85037 -80499 85081 -80455
rect 85137 -80499 85181 -80455
rect 85237 -80499 85281 -80455
rect 85337 -80499 85381 -80455
rect 85437 -80499 85481 -80455
rect 85537 -80499 85581 -80455
rect 85637 -80499 85681 -80455
rect 85737 -80499 85781 -80455
rect 85837 -80499 85881 -80455
rect 85937 -80499 85981 -80455
rect 86037 -80499 86081 -80455
rect 86137 -80499 86181 -80455
rect 86237 -80499 86281 -80455
rect 86737 -80499 86781 -80455
rect 86837 -80499 86881 -80455
rect 86937 -80499 86981 -80455
rect 87037 -80499 87081 -80455
rect 87137 -80499 87181 -80455
rect 87237 -80499 87281 -80455
rect 87337 -80499 87381 -80455
rect 87437 -80499 87481 -80455
rect 87537 -80499 87581 -80455
rect 87637 -80499 87681 -80455
rect 87737 -80499 87781 -80455
rect 87837 -80499 87881 -80455
rect 87937 -80499 87981 -80455
rect 88037 -80499 88081 -80455
rect 88137 -80499 88181 -80455
rect 88237 -80499 88281 -80455
rect -82968 -80603 -82924 -80559
rect -82868 -80603 -82824 -80559
rect -82768 -80603 -82724 -80559
rect -82668 -80603 -82624 -80559
rect -82568 -80603 -82524 -80559
rect -82468 -80603 -82424 -80559
rect -82368 -80603 -82324 -80559
rect -82268 -80603 -82224 -80559
rect -82168 -80603 -82124 -80559
rect -82068 -80603 -82024 -80559
rect -81968 -80603 -81924 -80559
rect -81868 -80603 -81824 -80559
rect -81768 -80603 -81724 -80559
rect -81668 -80603 -81624 -80559
rect -81568 -80603 -81524 -80559
rect -81468 -80603 -81424 -80559
rect -80968 -80603 -80924 -80559
rect -80868 -80603 -80824 -80559
rect -80768 -80603 -80724 -80559
rect -80668 -80603 -80624 -80559
rect -80568 -80603 -80524 -80559
rect -80468 -80603 -80424 -80559
rect -80368 -80603 -80324 -80559
rect -80268 -80603 -80224 -80559
rect -80168 -80603 -80124 -80559
rect -80068 -80603 -80024 -80559
rect -79968 -80603 -79924 -80559
rect -79868 -80603 -79824 -80559
rect -79768 -80603 -79724 -80559
rect -79668 -80603 -79624 -80559
rect -79568 -80603 -79524 -80559
rect -79468 -80603 -79424 -80559
rect -78968 -80603 -78924 -80559
rect -78868 -80603 -78824 -80559
rect -78768 -80603 -78724 -80559
rect -78668 -80603 -78624 -80559
rect -78568 -80603 -78524 -80559
rect -78468 -80603 -78424 -80559
rect -78368 -80603 -78324 -80559
rect -78268 -80603 -78224 -80559
rect -78168 -80603 -78124 -80559
rect -78068 -80603 -78024 -80559
rect -77968 -80603 -77924 -80559
rect -77868 -80603 -77824 -80559
rect -77768 -80603 -77724 -80559
rect -77668 -80603 -77624 -80559
rect -77568 -80603 -77524 -80559
rect -77468 -80603 -77424 -80559
rect -76968 -80603 -76924 -80559
rect -76868 -80603 -76824 -80559
rect -76768 -80603 -76724 -80559
rect -76668 -80603 -76624 -80559
rect -76568 -80603 -76524 -80559
rect -76468 -80603 -76424 -80559
rect -76368 -80603 -76324 -80559
rect -76268 -80603 -76224 -80559
rect -76168 -80603 -76124 -80559
rect -76068 -80603 -76024 -80559
rect -75968 -80603 -75924 -80559
rect -75868 -80603 -75824 -80559
rect -75768 -80603 -75724 -80559
rect -75668 -80603 -75624 -80559
rect -75568 -80603 -75524 -80559
rect -75468 -80603 -75424 -80559
rect -50017 -80605 -49973 -80561
rect -49917 -80605 -49873 -80561
rect -49817 -80605 -49773 -80561
rect -49717 -80605 -49673 -80561
rect -49617 -80605 -49573 -80561
rect -49517 -80605 -49473 -80561
rect -49417 -80605 -49373 -80561
rect -49317 -80605 -49273 -80561
rect -49217 -80605 -49173 -80561
rect -49117 -80605 -49073 -80561
rect -49017 -80605 -48973 -80561
rect -48917 -80605 -48873 -80561
rect -48817 -80605 -48773 -80561
rect -48717 -80605 -48673 -80561
rect -48617 -80605 -48573 -80561
rect -48517 -80605 -48473 -80561
rect -48017 -80605 -47973 -80561
rect -47917 -80605 -47873 -80561
rect -47817 -80605 -47773 -80561
rect -47717 -80605 -47673 -80561
rect -47617 -80605 -47573 -80561
rect -47517 -80605 -47473 -80561
rect -47417 -80605 -47373 -80561
rect -47317 -80605 -47273 -80561
rect -47217 -80605 -47173 -80561
rect -47117 -80605 -47073 -80561
rect -47017 -80605 -46973 -80561
rect -46917 -80605 -46873 -80561
rect -46817 -80605 -46773 -80561
rect -46717 -80605 -46673 -80561
rect -46617 -80605 -46573 -80561
rect -46517 -80605 -46473 -80561
rect -46017 -80605 -45973 -80561
rect -45917 -80605 -45873 -80561
rect -45817 -80605 -45773 -80561
rect -45717 -80605 -45673 -80561
rect -45617 -80605 -45573 -80561
rect -45517 -80605 -45473 -80561
rect -45417 -80605 -45373 -80561
rect -45317 -80605 -45273 -80561
rect -45217 -80605 -45173 -80561
rect -45117 -80605 -45073 -80561
rect -45017 -80605 -44973 -80561
rect -44917 -80605 -44873 -80561
rect -44817 -80605 -44773 -80561
rect -44717 -80605 -44673 -80561
rect -44617 -80605 -44573 -80561
rect -44517 -80605 -44473 -80561
rect -44017 -80605 -43973 -80561
rect -43917 -80605 -43873 -80561
rect -43817 -80605 -43773 -80561
rect -43717 -80605 -43673 -80561
rect -43617 -80605 -43573 -80561
rect -43517 -80605 -43473 -80561
rect -43417 -80605 -43373 -80561
rect -43317 -80605 -43273 -80561
rect -43217 -80605 -43173 -80561
rect -43117 -80605 -43073 -80561
rect -43017 -80605 -42973 -80561
rect -42917 -80605 -42873 -80561
rect -42817 -80605 -42773 -80561
rect -42717 -80605 -42673 -80561
rect -42617 -80605 -42573 -80561
rect -42517 -80605 -42473 -80561
rect 80737 -80599 80781 -80555
rect 80837 -80599 80881 -80555
rect 80937 -80599 80981 -80555
rect 81037 -80599 81081 -80555
rect 81137 -80599 81181 -80555
rect 81237 -80599 81281 -80555
rect 81337 -80599 81381 -80555
rect 81437 -80599 81481 -80555
rect 81537 -80599 81581 -80555
rect 81637 -80599 81681 -80555
rect 81737 -80599 81781 -80555
rect 81837 -80599 81881 -80555
rect 81937 -80599 81981 -80555
rect 82037 -80599 82081 -80555
rect 82137 -80599 82181 -80555
rect 82237 -80599 82281 -80555
rect 82737 -80599 82781 -80555
rect 82837 -80599 82881 -80555
rect 82937 -80599 82981 -80555
rect 83037 -80599 83081 -80555
rect 83137 -80599 83181 -80555
rect 83237 -80599 83281 -80555
rect 83337 -80599 83381 -80555
rect 83437 -80599 83481 -80555
rect 83537 -80599 83581 -80555
rect 83637 -80599 83681 -80555
rect 83737 -80599 83781 -80555
rect 83837 -80599 83881 -80555
rect 83937 -80599 83981 -80555
rect 84037 -80599 84081 -80555
rect 84137 -80599 84181 -80555
rect 84237 -80599 84281 -80555
rect 84737 -80599 84781 -80555
rect 84837 -80599 84881 -80555
rect 84937 -80599 84981 -80555
rect 85037 -80599 85081 -80555
rect 85137 -80599 85181 -80555
rect 85237 -80599 85281 -80555
rect 85337 -80599 85381 -80555
rect 85437 -80599 85481 -80555
rect 85537 -80599 85581 -80555
rect 85637 -80599 85681 -80555
rect 85737 -80599 85781 -80555
rect 85837 -80599 85881 -80555
rect 85937 -80599 85981 -80555
rect 86037 -80599 86081 -80555
rect 86137 -80599 86181 -80555
rect 86237 -80599 86281 -80555
rect 86737 -80599 86781 -80555
rect 86837 -80599 86881 -80555
rect 86937 -80599 86981 -80555
rect 87037 -80599 87081 -80555
rect 87137 -80599 87181 -80555
rect 87237 -80599 87281 -80555
rect 87337 -80599 87381 -80555
rect 87437 -80599 87481 -80555
rect 87537 -80599 87581 -80555
rect 87637 -80599 87681 -80555
rect 87737 -80599 87781 -80555
rect 87837 -80599 87881 -80555
rect 87937 -80599 87981 -80555
rect 88037 -80599 88081 -80555
rect 88137 -80599 88181 -80555
rect 88237 -80599 88281 -80555
rect -82968 -80703 -82924 -80659
rect -82868 -80703 -82824 -80659
rect -82768 -80703 -82724 -80659
rect -82668 -80703 -82624 -80659
rect -82568 -80703 -82524 -80659
rect -82468 -80703 -82424 -80659
rect -82368 -80703 -82324 -80659
rect -82268 -80703 -82224 -80659
rect -82168 -80703 -82124 -80659
rect -82068 -80703 -82024 -80659
rect -81968 -80703 -81924 -80659
rect -81868 -80703 -81824 -80659
rect -81768 -80703 -81724 -80659
rect -81668 -80703 -81624 -80659
rect -81568 -80703 -81524 -80659
rect -81468 -80703 -81424 -80659
rect -80968 -80703 -80924 -80659
rect -80868 -80703 -80824 -80659
rect -80768 -80703 -80724 -80659
rect -80668 -80703 -80624 -80659
rect -80568 -80703 -80524 -80659
rect -80468 -80703 -80424 -80659
rect -80368 -80703 -80324 -80659
rect -80268 -80703 -80224 -80659
rect -80168 -80703 -80124 -80659
rect -80068 -80703 -80024 -80659
rect -79968 -80703 -79924 -80659
rect -79868 -80703 -79824 -80659
rect -79768 -80703 -79724 -80659
rect -79668 -80703 -79624 -80659
rect -79568 -80703 -79524 -80659
rect -79468 -80703 -79424 -80659
rect -78968 -80703 -78924 -80659
rect -78868 -80703 -78824 -80659
rect -78768 -80703 -78724 -80659
rect -78668 -80703 -78624 -80659
rect -78568 -80703 -78524 -80659
rect -78468 -80703 -78424 -80659
rect -78368 -80703 -78324 -80659
rect -78268 -80703 -78224 -80659
rect -78168 -80703 -78124 -80659
rect -78068 -80703 -78024 -80659
rect -77968 -80703 -77924 -80659
rect -77868 -80703 -77824 -80659
rect -77768 -80703 -77724 -80659
rect -77668 -80703 -77624 -80659
rect -77568 -80703 -77524 -80659
rect -77468 -80703 -77424 -80659
rect -76968 -80703 -76924 -80659
rect -76868 -80703 -76824 -80659
rect -76768 -80703 -76724 -80659
rect -76668 -80703 -76624 -80659
rect -76568 -80703 -76524 -80659
rect -76468 -80703 -76424 -80659
rect -76368 -80703 -76324 -80659
rect -76268 -80703 -76224 -80659
rect -76168 -80703 -76124 -80659
rect -76068 -80703 -76024 -80659
rect -75968 -80703 -75924 -80659
rect -75868 -80703 -75824 -80659
rect -75768 -80703 -75724 -80659
rect -75668 -80703 -75624 -80659
rect -75568 -80703 -75524 -80659
rect -75468 -80703 -75424 -80659
rect -50017 -80705 -49973 -80661
rect -49917 -80705 -49873 -80661
rect -49817 -80705 -49773 -80661
rect -49717 -80705 -49673 -80661
rect -49617 -80705 -49573 -80661
rect -49517 -80705 -49473 -80661
rect -49417 -80705 -49373 -80661
rect -49317 -80705 -49273 -80661
rect -49217 -80705 -49173 -80661
rect -49117 -80705 -49073 -80661
rect -49017 -80705 -48973 -80661
rect -48917 -80705 -48873 -80661
rect -48817 -80705 -48773 -80661
rect -48717 -80705 -48673 -80661
rect -48617 -80705 -48573 -80661
rect -48517 -80705 -48473 -80661
rect -48017 -80705 -47973 -80661
rect -47917 -80705 -47873 -80661
rect -47817 -80705 -47773 -80661
rect -47717 -80705 -47673 -80661
rect -47617 -80705 -47573 -80661
rect -47517 -80705 -47473 -80661
rect -47417 -80705 -47373 -80661
rect -47317 -80705 -47273 -80661
rect -47217 -80705 -47173 -80661
rect -47117 -80705 -47073 -80661
rect -47017 -80705 -46973 -80661
rect -46917 -80705 -46873 -80661
rect -46817 -80705 -46773 -80661
rect -46717 -80705 -46673 -80661
rect -46617 -80705 -46573 -80661
rect -46517 -80705 -46473 -80661
rect -46017 -80705 -45973 -80661
rect -45917 -80705 -45873 -80661
rect -45817 -80705 -45773 -80661
rect -45717 -80705 -45673 -80661
rect -45617 -80705 -45573 -80661
rect -45517 -80705 -45473 -80661
rect -45417 -80705 -45373 -80661
rect -45317 -80705 -45273 -80661
rect -45217 -80705 -45173 -80661
rect -45117 -80705 -45073 -80661
rect -45017 -80705 -44973 -80661
rect -44917 -80705 -44873 -80661
rect -44817 -80705 -44773 -80661
rect -44717 -80705 -44673 -80661
rect -44617 -80705 -44573 -80661
rect -44517 -80705 -44473 -80661
rect -44017 -80705 -43973 -80661
rect -43917 -80705 -43873 -80661
rect -43817 -80705 -43773 -80661
rect -43717 -80705 -43673 -80661
rect -43617 -80705 -43573 -80661
rect -43517 -80705 -43473 -80661
rect -43417 -80705 -43373 -80661
rect -43317 -80705 -43273 -80661
rect -43217 -80705 -43173 -80661
rect -43117 -80705 -43073 -80661
rect -43017 -80705 -42973 -80661
rect -42917 -80705 -42873 -80661
rect -42817 -80705 -42773 -80661
rect -42717 -80705 -42673 -80661
rect -42617 -80705 -42573 -80661
rect -42517 -80705 -42473 -80661
rect 80737 -80699 80781 -80655
rect 80837 -80699 80881 -80655
rect 80937 -80699 80981 -80655
rect 81037 -80699 81081 -80655
rect 81137 -80699 81181 -80655
rect 81237 -80699 81281 -80655
rect 81337 -80699 81381 -80655
rect 81437 -80699 81481 -80655
rect 81537 -80699 81581 -80655
rect 81637 -80699 81681 -80655
rect 81737 -80699 81781 -80655
rect 81837 -80699 81881 -80655
rect 81937 -80699 81981 -80655
rect 82037 -80699 82081 -80655
rect 82137 -80699 82181 -80655
rect 82237 -80699 82281 -80655
rect 82737 -80699 82781 -80655
rect 82837 -80699 82881 -80655
rect 82937 -80699 82981 -80655
rect 83037 -80699 83081 -80655
rect 83137 -80699 83181 -80655
rect 83237 -80699 83281 -80655
rect 83337 -80699 83381 -80655
rect 83437 -80699 83481 -80655
rect 83537 -80699 83581 -80655
rect 83637 -80699 83681 -80655
rect 83737 -80699 83781 -80655
rect 83837 -80699 83881 -80655
rect 83937 -80699 83981 -80655
rect 84037 -80699 84081 -80655
rect 84137 -80699 84181 -80655
rect 84237 -80699 84281 -80655
rect 84737 -80699 84781 -80655
rect 84837 -80699 84881 -80655
rect 84937 -80699 84981 -80655
rect 85037 -80699 85081 -80655
rect 85137 -80699 85181 -80655
rect 85237 -80699 85281 -80655
rect 85337 -80699 85381 -80655
rect 85437 -80699 85481 -80655
rect 85537 -80699 85581 -80655
rect 85637 -80699 85681 -80655
rect 85737 -80699 85781 -80655
rect 85837 -80699 85881 -80655
rect 85937 -80699 85981 -80655
rect 86037 -80699 86081 -80655
rect 86137 -80699 86181 -80655
rect 86237 -80699 86281 -80655
rect 86737 -80699 86781 -80655
rect 86837 -80699 86881 -80655
rect 86937 -80699 86981 -80655
rect 87037 -80699 87081 -80655
rect 87137 -80699 87181 -80655
rect 87237 -80699 87281 -80655
rect 87337 -80699 87381 -80655
rect 87437 -80699 87481 -80655
rect 87537 -80699 87581 -80655
rect 87637 -80699 87681 -80655
rect 87737 -80699 87781 -80655
rect 87837 -80699 87881 -80655
rect 87937 -80699 87981 -80655
rect 88037 -80699 88081 -80655
rect 88137 -80699 88181 -80655
rect 88237 -80699 88281 -80655
rect -82968 -80803 -82924 -80759
rect -82868 -80803 -82824 -80759
rect -82768 -80803 -82724 -80759
rect -82668 -80803 -82624 -80759
rect -82568 -80803 -82524 -80759
rect -82468 -80803 -82424 -80759
rect -82368 -80803 -82324 -80759
rect -82268 -80803 -82224 -80759
rect -82168 -80803 -82124 -80759
rect -82068 -80803 -82024 -80759
rect -81968 -80803 -81924 -80759
rect -81868 -80803 -81824 -80759
rect -81768 -80803 -81724 -80759
rect -81668 -80803 -81624 -80759
rect -81568 -80803 -81524 -80759
rect -81468 -80803 -81424 -80759
rect -80968 -80803 -80924 -80759
rect -80868 -80803 -80824 -80759
rect -80768 -80803 -80724 -80759
rect -80668 -80803 -80624 -80759
rect -80568 -80803 -80524 -80759
rect -80468 -80803 -80424 -80759
rect -80368 -80803 -80324 -80759
rect -80268 -80803 -80224 -80759
rect -80168 -80803 -80124 -80759
rect -80068 -80803 -80024 -80759
rect -79968 -80803 -79924 -80759
rect -79868 -80803 -79824 -80759
rect -79768 -80803 -79724 -80759
rect -79668 -80803 -79624 -80759
rect -79568 -80803 -79524 -80759
rect -79468 -80803 -79424 -80759
rect -78968 -80803 -78924 -80759
rect -78868 -80803 -78824 -80759
rect -78768 -80803 -78724 -80759
rect -78668 -80803 -78624 -80759
rect -78568 -80803 -78524 -80759
rect -78468 -80803 -78424 -80759
rect -78368 -80803 -78324 -80759
rect -78268 -80803 -78224 -80759
rect -78168 -80803 -78124 -80759
rect -78068 -80803 -78024 -80759
rect -77968 -80803 -77924 -80759
rect -77868 -80803 -77824 -80759
rect -77768 -80803 -77724 -80759
rect -77668 -80803 -77624 -80759
rect -77568 -80803 -77524 -80759
rect -77468 -80803 -77424 -80759
rect -76968 -80803 -76924 -80759
rect -76868 -80803 -76824 -80759
rect -76768 -80803 -76724 -80759
rect -76668 -80803 -76624 -80759
rect -76568 -80803 -76524 -80759
rect -76468 -80803 -76424 -80759
rect -76368 -80803 -76324 -80759
rect -76268 -80803 -76224 -80759
rect -76168 -80803 -76124 -80759
rect -76068 -80803 -76024 -80759
rect -75968 -80803 -75924 -80759
rect -75868 -80803 -75824 -80759
rect -75768 -80803 -75724 -80759
rect -75668 -80803 -75624 -80759
rect -75568 -80803 -75524 -80759
rect -75468 -80803 -75424 -80759
rect -50017 -80805 -49973 -80761
rect -49917 -80805 -49873 -80761
rect -49817 -80805 -49773 -80761
rect -49717 -80805 -49673 -80761
rect -49617 -80805 -49573 -80761
rect -49517 -80805 -49473 -80761
rect -49417 -80805 -49373 -80761
rect -49317 -80805 -49273 -80761
rect -49217 -80805 -49173 -80761
rect -49117 -80805 -49073 -80761
rect -49017 -80805 -48973 -80761
rect -48917 -80805 -48873 -80761
rect -48817 -80805 -48773 -80761
rect -48717 -80805 -48673 -80761
rect -48617 -80805 -48573 -80761
rect -48517 -80805 -48473 -80761
rect -48017 -80805 -47973 -80761
rect -47917 -80805 -47873 -80761
rect -47817 -80805 -47773 -80761
rect -47717 -80805 -47673 -80761
rect -47617 -80805 -47573 -80761
rect -47517 -80805 -47473 -80761
rect -47417 -80805 -47373 -80761
rect -47317 -80805 -47273 -80761
rect -47217 -80805 -47173 -80761
rect -47117 -80805 -47073 -80761
rect -47017 -80805 -46973 -80761
rect -46917 -80805 -46873 -80761
rect -46817 -80805 -46773 -80761
rect -46717 -80805 -46673 -80761
rect -46617 -80805 -46573 -80761
rect -46517 -80805 -46473 -80761
rect -46017 -80805 -45973 -80761
rect -45917 -80805 -45873 -80761
rect -45817 -80805 -45773 -80761
rect -45717 -80805 -45673 -80761
rect -45617 -80805 -45573 -80761
rect -45517 -80805 -45473 -80761
rect -45417 -80805 -45373 -80761
rect -45317 -80805 -45273 -80761
rect -45217 -80805 -45173 -80761
rect -45117 -80805 -45073 -80761
rect -45017 -80805 -44973 -80761
rect -44917 -80805 -44873 -80761
rect -44817 -80805 -44773 -80761
rect -44717 -80805 -44673 -80761
rect -44617 -80805 -44573 -80761
rect -44517 -80805 -44473 -80761
rect -44017 -80805 -43973 -80761
rect -43917 -80805 -43873 -80761
rect -43817 -80805 -43773 -80761
rect -43717 -80805 -43673 -80761
rect -43617 -80805 -43573 -80761
rect -43517 -80805 -43473 -80761
rect -43417 -80805 -43373 -80761
rect -43317 -80805 -43273 -80761
rect -43217 -80805 -43173 -80761
rect -43117 -80805 -43073 -80761
rect -43017 -80805 -42973 -80761
rect -42917 -80805 -42873 -80761
rect -42817 -80805 -42773 -80761
rect -42717 -80805 -42673 -80761
rect -42617 -80805 -42573 -80761
rect -42517 -80805 -42473 -80761
rect 80737 -80799 80781 -80755
rect 80837 -80799 80881 -80755
rect 80937 -80799 80981 -80755
rect 81037 -80799 81081 -80755
rect 81137 -80799 81181 -80755
rect 81237 -80799 81281 -80755
rect 81337 -80799 81381 -80755
rect 81437 -80799 81481 -80755
rect 81537 -80799 81581 -80755
rect 81637 -80799 81681 -80755
rect 81737 -80799 81781 -80755
rect 81837 -80799 81881 -80755
rect 81937 -80799 81981 -80755
rect 82037 -80799 82081 -80755
rect 82137 -80799 82181 -80755
rect 82237 -80799 82281 -80755
rect 82737 -80799 82781 -80755
rect 82837 -80799 82881 -80755
rect 82937 -80799 82981 -80755
rect 83037 -80799 83081 -80755
rect 83137 -80799 83181 -80755
rect 83237 -80799 83281 -80755
rect 83337 -80799 83381 -80755
rect 83437 -80799 83481 -80755
rect 83537 -80799 83581 -80755
rect 83637 -80799 83681 -80755
rect 83737 -80799 83781 -80755
rect 83837 -80799 83881 -80755
rect 83937 -80799 83981 -80755
rect 84037 -80799 84081 -80755
rect 84137 -80799 84181 -80755
rect 84237 -80799 84281 -80755
rect 84737 -80799 84781 -80755
rect 84837 -80799 84881 -80755
rect 84937 -80799 84981 -80755
rect 85037 -80799 85081 -80755
rect 85137 -80799 85181 -80755
rect 85237 -80799 85281 -80755
rect 85337 -80799 85381 -80755
rect 85437 -80799 85481 -80755
rect 85537 -80799 85581 -80755
rect 85637 -80799 85681 -80755
rect 85737 -80799 85781 -80755
rect 85837 -80799 85881 -80755
rect 85937 -80799 85981 -80755
rect 86037 -80799 86081 -80755
rect 86137 -80799 86181 -80755
rect 86237 -80799 86281 -80755
rect 86737 -80799 86781 -80755
rect 86837 -80799 86881 -80755
rect 86937 -80799 86981 -80755
rect 87037 -80799 87081 -80755
rect 87137 -80799 87181 -80755
rect 87237 -80799 87281 -80755
rect 87337 -80799 87381 -80755
rect 87437 -80799 87481 -80755
rect 87537 -80799 87581 -80755
rect 87637 -80799 87681 -80755
rect 87737 -80799 87781 -80755
rect 87837 -80799 87881 -80755
rect 87937 -80799 87981 -80755
rect 88037 -80799 88081 -80755
rect 88137 -80799 88181 -80755
rect 88237 -80799 88281 -80755
rect -82968 -80903 -82924 -80859
rect -82868 -80903 -82824 -80859
rect -82768 -80903 -82724 -80859
rect -82668 -80903 -82624 -80859
rect -82568 -80903 -82524 -80859
rect -82468 -80903 -82424 -80859
rect -82368 -80903 -82324 -80859
rect -82268 -80903 -82224 -80859
rect -82168 -80903 -82124 -80859
rect -82068 -80903 -82024 -80859
rect -81968 -80903 -81924 -80859
rect -81868 -80903 -81824 -80859
rect -81768 -80903 -81724 -80859
rect -81668 -80903 -81624 -80859
rect -81568 -80903 -81524 -80859
rect -81468 -80903 -81424 -80859
rect -80968 -80903 -80924 -80859
rect -80868 -80903 -80824 -80859
rect -80768 -80903 -80724 -80859
rect -80668 -80903 -80624 -80859
rect -80568 -80903 -80524 -80859
rect -80468 -80903 -80424 -80859
rect -80368 -80903 -80324 -80859
rect -80268 -80903 -80224 -80859
rect -80168 -80903 -80124 -80859
rect -80068 -80903 -80024 -80859
rect -79968 -80903 -79924 -80859
rect -79868 -80903 -79824 -80859
rect -79768 -80903 -79724 -80859
rect -79668 -80903 -79624 -80859
rect -79568 -80903 -79524 -80859
rect -79468 -80903 -79424 -80859
rect -78968 -80903 -78924 -80859
rect -78868 -80903 -78824 -80859
rect -78768 -80903 -78724 -80859
rect -78668 -80903 -78624 -80859
rect -78568 -80903 -78524 -80859
rect -78468 -80903 -78424 -80859
rect -78368 -80903 -78324 -80859
rect -78268 -80903 -78224 -80859
rect -78168 -80903 -78124 -80859
rect -78068 -80903 -78024 -80859
rect -77968 -80903 -77924 -80859
rect -77868 -80903 -77824 -80859
rect -77768 -80903 -77724 -80859
rect -77668 -80903 -77624 -80859
rect -77568 -80903 -77524 -80859
rect -77468 -80903 -77424 -80859
rect -76968 -80903 -76924 -80859
rect -76868 -80903 -76824 -80859
rect -76768 -80903 -76724 -80859
rect -76668 -80903 -76624 -80859
rect -76568 -80903 -76524 -80859
rect -76468 -80903 -76424 -80859
rect -76368 -80903 -76324 -80859
rect -76268 -80903 -76224 -80859
rect -76168 -80903 -76124 -80859
rect -76068 -80903 -76024 -80859
rect -75968 -80903 -75924 -80859
rect -75868 -80903 -75824 -80859
rect -75768 -80903 -75724 -80859
rect -75668 -80903 -75624 -80859
rect -75568 -80903 -75524 -80859
rect -75468 -80903 -75424 -80859
rect -50017 -80905 -49973 -80861
rect -49917 -80905 -49873 -80861
rect -49817 -80905 -49773 -80861
rect -49717 -80905 -49673 -80861
rect -49617 -80905 -49573 -80861
rect -49517 -80905 -49473 -80861
rect -49417 -80905 -49373 -80861
rect -49317 -80905 -49273 -80861
rect -49217 -80905 -49173 -80861
rect -49117 -80905 -49073 -80861
rect -49017 -80905 -48973 -80861
rect -48917 -80905 -48873 -80861
rect -48817 -80905 -48773 -80861
rect -48717 -80905 -48673 -80861
rect -48617 -80905 -48573 -80861
rect -48517 -80905 -48473 -80861
rect -48017 -80905 -47973 -80861
rect -47917 -80905 -47873 -80861
rect -47817 -80905 -47773 -80861
rect -47717 -80905 -47673 -80861
rect -47617 -80905 -47573 -80861
rect -47517 -80905 -47473 -80861
rect -47417 -80905 -47373 -80861
rect -47317 -80905 -47273 -80861
rect -47217 -80905 -47173 -80861
rect -47117 -80905 -47073 -80861
rect -47017 -80905 -46973 -80861
rect -46917 -80905 -46873 -80861
rect -46817 -80905 -46773 -80861
rect -46717 -80905 -46673 -80861
rect -46617 -80905 -46573 -80861
rect -46517 -80905 -46473 -80861
rect -46017 -80905 -45973 -80861
rect -45917 -80905 -45873 -80861
rect -45817 -80905 -45773 -80861
rect -45717 -80905 -45673 -80861
rect -45617 -80905 -45573 -80861
rect -45517 -80905 -45473 -80861
rect -45417 -80905 -45373 -80861
rect -45317 -80905 -45273 -80861
rect -45217 -80905 -45173 -80861
rect -45117 -80905 -45073 -80861
rect -45017 -80905 -44973 -80861
rect -44917 -80905 -44873 -80861
rect -44817 -80905 -44773 -80861
rect -44717 -80905 -44673 -80861
rect -44617 -80905 -44573 -80861
rect -44517 -80905 -44473 -80861
rect -44017 -80905 -43973 -80861
rect -43917 -80905 -43873 -80861
rect -43817 -80905 -43773 -80861
rect -43717 -80905 -43673 -80861
rect -43617 -80905 -43573 -80861
rect -43517 -80905 -43473 -80861
rect -43417 -80905 -43373 -80861
rect -43317 -80905 -43273 -80861
rect -43217 -80905 -43173 -80861
rect -43117 -80905 -43073 -80861
rect -43017 -80905 -42973 -80861
rect -42917 -80905 -42873 -80861
rect -42817 -80905 -42773 -80861
rect -42717 -80905 -42673 -80861
rect -42617 -80905 -42573 -80861
rect -42517 -80905 -42473 -80861
rect 80737 -80899 80781 -80855
rect 80837 -80899 80881 -80855
rect 80937 -80899 80981 -80855
rect 81037 -80899 81081 -80855
rect 81137 -80899 81181 -80855
rect 81237 -80899 81281 -80855
rect 81337 -80899 81381 -80855
rect 81437 -80899 81481 -80855
rect 81537 -80899 81581 -80855
rect 81637 -80899 81681 -80855
rect 81737 -80899 81781 -80855
rect 81837 -80899 81881 -80855
rect 81937 -80899 81981 -80855
rect 82037 -80899 82081 -80855
rect 82137 -80899 82181 -80855
rect 82237 -80899 82281 -80855
rect 82737 -80899 82781 -80855
rect 82837 -80899 82881 -80855
rect 82937 -80899 82981 -80855
rect 83037 -80899 83081 -80855
rect 83137 -80899 83181 -80855
rect 83237 -80899 83281 -80855
rect 83337 -80899 83381 -80855
rect 83437 -80899 83481 -80855
rect 83537 -80899 83581 -80855
rect 83637 -80899 83681 -80855
rect 83737 -80899 83781 -80855
rect 83837 -80899 83881 -80855
rect 83937 -80899 83981 -80855
rect 84037 -80899 84081 -80855
rect 84137 -80899 84181 -80855
rect 84237 -80899 84281 -80855
rect 84737 -80899 84781 -80855
rect 84837 -80899 84881 -80855
rect 84937 -80899 84981 -80855
rect 85037 -80899 85081 -80855
rect 85137 -80899 85181 -80855
rect 85237 -80899 85281 -80855
rect 85337 -80899 85381 -80855
rect 85437 -80899 85481 -80855
rect 85537 -80899 85581 -80855
rect 85637 -80899 85681 -80855
rect 85737 -80899 85781 -80855
rect 85837 -80899 85881 -80855
rect 85937 -80899 85981 -80855
rect 86037 -80899 86081 -80855
rect 86137 -80899 86181 -80855
rect 86237 -80899 86281 -80855
rect 86737 -80899 86781 -80855
rect 86837 -80899 86881 -80855
rect 86937 -80899 86981 -80855
rect 87037 -80899 87081 -80855
rect 87137 -80899 87181 -80855
rect 87237 -80899 87281 -80855
rect 87337 -80899 87381 -80855
rect 87437 -80899 87481 -80855
rect 87537 -80899 87581 -80855
rect 87637 -80899 87681 -80855
rect 87737 -80899 87781 -80855
rect 87837 -80899 87881 -80855
rect 87937 -80899 87981 -80855
rect 88037 -80899 88081 -80855
rect 88137 -80899 88181 -80855
rect 88237 -80899 88281 -80855
rect -82968 -81003 -82924 -80959
rect -82868 -81003 -82824 -80959
rect -82768 -81003 -82724 -80959
rect -82668 -81003 -82624 -80959
rect -82568 -81003 -82524 -80959
rect -82468 -81003 -82424 -80959
rect -82368 -81003 -82324 -80959
rect -82268 -81003 -82224 -80959
rect -82168 -81003 -82124 -80959
rect -82068 -81003 -82024 -80959
rect -81968 -81003 -81924 -80959
rect -81868 -81003 -81824 -80959
rect -81768 -81003 -81724 -80959
rect -81668 -81003 -81624 -80959
rect -81568 -81003 -81524 -80959
rect -81468 -81003 -81424 -80959
rect -80968 -81003 -80924 -80959
rect -80868 -81003 -80824 -80959
rect -80768 -81003 -80724 -80959
rect -80668 -81003 -80624 -80959
rect -80568 -81003 -80524 -80959
rect -80468 -81003 -80424 -80959
rect -80368 -81003 -80324 -80959
rect -80268 -81003 -80224 -80959
rect -80168 -81003 -80124 -80959
rect -80068 -81003 -80024 -80959
rect -79968 -81003 -79924 -80959
rect -79868 -81003 -79824 -80959
rect -79768 -81003 -79724 -80959
rect -79668 -81003 -79624 -80959
rect -79568 -81003 -79524 -80959
rect -79468 -81003 -79424 -80959
rect -78968 -81003 -78924 -80959
rect -78868 -81003 -78824 -80959
rect -78768 -81003 -78724 -80959
rect -78668 -81003 -78624 -80959
rect -78568 -81003 -78524 -80959
rect -78468 -81003 -78424 -80959
rect -78368 -81003 -78324 -80959
rect -78268 -81003 -78224 -80959
rect -78168 -81003 -78124 -80959
rect -78068 -81003 -78024 -80959
rect -77968 -81003 -77924 -80959
rect -77868 -81003 -77824 -80959
rect -77768 -81003 -77724 -80959
rect -77668 -81003 -77624 -80959
rect -77568 -81003 -77524 -80959
rect -77468 -81003 -77424 -80959
rect -76968 -81003 -76924 -80959
rect -76868 -81003 -76824 -80959
rect -76768 -81003 -76724 -80959
rect -76668 -81003 -76624 -80959
rect -76568 -81003 -76524 -80959
rect -76468 -81003 -76424 -80959
rect -76368 -81003 -76324 -80959
rect -76268 -81003 -76224 -80959
rect -76168 -81003 -76124 -80959
rect -76068 -81003 -76024 -80959
rect -75968 -81003 -75924 -80959
rect -75868 -81003 -75824 -80959
rect -75768 -81003 -75724 -80959
rect -75668 -81003 -75624 -80959
rect -75568 -81003 -75524 -80959
rect -75468 -81003 -75424 -80959
rect -50017 -81005 -49973 -80961
rect -49917 -81005 -49873 -80961
rect -49817 -81005 -49773 -80961
rect -49717 -81005 -49673 -80961
rect -49617 -81005 -49573 -80961
rect -49517 -81005 -49473 -80961
rect -49417 -81005 -49373 -80961
rect -49317 -81005 -49273 -80961
rect -49217 -81005 -49173 -80961
rect -49117 -81005 -49073 -80961
rect -49017 -81005 -48973 -80961
rect -48917 -81005 -48873 -80961
rect -48817 -81005 -48773 -80961
rect -48717 -81005 -48673 -80961
rect -48617 -81005 -48573 -80961
rect -48517 -81005 -48473 -80961
rect -48017 -81005 -47973 -80961
rect -47917 -81005 -47873 -80961
rect -47817 -81005 -47773 -80961
rect -47717 -81005 -47673 -80961
rect -47617 -81005 -47573 -80961
rect -47517 -81005 -47473 -80961
rect -47417 -81005 -47373 -80961
rect -47317 -81005 -47273 -80961
rect -47217 -81005 -47173 -80961
rect -47117 -81005 -47073 -80961
rect -47017 -81005 -46973 -80961
rect -46917 -81005 -46873 -80961
rect -46817 -81005 -46773 -80961
rect -46717 -81005 -46673 -80961
rect -46617 -81005 -46573 -80961
rect -46517 -81005 -46473 -80961
rect -46017 -81005 -45973 -80961
rect -45917 -81005 -45873 -80961
rect -45817 -81005 -45773 -80961
rect -45717 -81005 -45673 -80961
rect -45617 -81005 -45573 -80961
rect -45517 -81005 -45473 -80961
rect -45417 -81005 -45373 -80961
rect -45317 -81005 -45273 -80961
rect -45217 -81005 -45173 -80961
rect -45117 -81005 -45073 -80961
rect -45017 -81005 -44973 -80961
rect -44917 -81005 -44873 -80961
rect -44817 -81005 -44773 -80961
rect -44717 -81005 -44673 -80961
rect -44617 -81005 -44573 -80961
rect -44517 -81005 -44473 -80961
rect -44017 -81005 -43973 -80961
rect -43917 -81005 -43873 -80961
rect -43817 -81005 -43773 -80961
rect -43717 -81005 -43673 -80961
rect -43617 -81005 -43573 -80961
rect -43517 -81005 -43473 -80961
rect -43417 -81005 -43373 -80961
rect -43317 -81005 -43273 -80961
rect -43217 -81005 -43173 -80961
rect -43117 -81005 -43073 -80961
rect -43017 -81005 -42973 -80961
rect -42917 -81005 -42873 -80961
rect -42817 -81005 -42773 -80961
rect -42717 -81005 -42673 -80961
rect -42617 -81005 -42573 -80961
rect -42517 -81005 -42473 -80961
rect 80737 -80999 80781 -80955
rect 80837 -80999 80881 -80955
rect 80937 -80999 80981 -80955
rect 81037 -80999 81081 -80955
rect 81137 -80999 81181 -80955
rect 81237 -80999 81281 -80955
rect 81337 -80999 81381 -80955
rect 81437 -80999 81481 -80955
rect 81537 -80999 81581 -80955
rect 81637 -80999 81681 -80955
rect 81737 -80999 81781 -80955
rect 81837 -80999 81881 -80955
rect 81937 -80999 81981 -80955
rect 82037 -80999 82081 -80955
rect 82137 -80999 82181 -80955
rect 82237 -80999 82281 -80955
rect 82737 -80999 82781 -80955
rect 82837 -80999 82881 -80955
rect 82937 -80999 82981 -80955
rect 83037 -80999 83081 -80955
rect 83137 -80999 83181 -80955
rect 83237 -80999 83281 -80955
rect 83337 -80999 83381 -80955
rect 83437 -80999 83481 -80955
rect 83537 -80999 83581 -80955
rect 83637 -80999 83681 -80955
rect 83737 -80999 83781 -80955
rect 83837 -80999 83881 -80955
rect 83937 -80999 83981 -80955
rect 84037 -80999 84081 -80955
rect 84137 -80999 84181 -80955
rect 84237 -80999 84281 -80955
rect 84737 -80999 84781 -80955
rect 84837 -80999 84881 -80955
rect 84937 -80999 84981 -80955
rect 85037 -80999 85081 -80955
rect 85137 -80999 85181 -80955
rect 85237 -80999 85281 -80955
rect 85337 -80999 85381 -80955
rect 85437 -80999 85481 -80955
rect 85537 -80999 85581 -80955
rect 85637 -80999 85681 -80955
rect 85737 -80999 85781 -80955
rect 85837 -80999 85881 -80955
rect 85937 -80999 85981 -80955
rect 86037 -80999 86081 -80955
rect 86137 -80999 86181 -80955
rect 86237 -80999 86281 -80955
rect 86737 -80999 86781 -80955
rect 86837 -80999 86881 -80955
rect 86937 -80999 86981 -80955
rect 87037 -80999 87081 -80955
rect 87137 -80999 87181 -80955
rect 87237 -80999 87281 -80955
rect 87337 -80999 87381 -80955
rect 87437 -80999 87481 -80955
rect 87537 -80999 87581 -80955
rect 87637 -80999 87681 -80955
rect 87737 -80999 87781 -80955
rect 87837 -80999 87881 -80955
rect 87937 -80999 87981 -80955
rect 88037 -80999 88081 -80955
rect 88137 -80999 88181 -80955
rect 88237 -80999 88281 -80955
rect -82968 -81103 -82924 -81059
rect -82868 -81103 -82824 -81059
rect -82768 -81103 -82724 -81059
rect -82668 -81103 -82624 -81059
rect -82568 -81103 -82524 -81059
rect -82468 -81103 -82424 -81059
rect -82368 -81103 -82324 -81059
rect -82268 -81103 -82224 -81059
rect -82168 -81103 -82124 -81059
rect -82068 -81103 -82024 -81059
rect -81968 -81103 -81924 -81059
rect -81868 -81103 -81824 -81059
rect -81768 -81103 -81724 -81059
rect -81668 -81103 -81624 -81059
rect -81568 -81103 -81524 -81059
rect -81468 -81103 -81424 -81059
rect -80968 -81103 -80924 -81059
rect -80868 -81103 -80824 -81059
rect -80768 -81103 -80724 -81059
rect -80668 -81103 -80624 -81059
rect -80568 -81103 -80524 -81059
rect -80468 -81103 -80424 -81059
rect -80368 -81103 -80324 -81059
rect -80268 -81103 -80224 -81059
rect -80168 -81103 -80124 -81059
rect -80068 -81103 -80024 -81059
rect -79968 -81103 -79924 -81059
rect -79868 -81103 -79824 -81059
rect -79768 -81103 -79724 -81059
rect -79668 -81103 -79624 -81059
rect -79568 -81103 -79524 -81059
rect -79468 -81103 -79424 -81059
rect -78968 -81103 -78924 -81059
rect -78868 -81103 -78824 -81059
rect -78768 -81103 -78724 -81059
rect -78668 -81103 -78624 -81059
rect -78568 -81103 -78524 -81059
rect -78468 -81103 -78424 -81059
rect -78368 -81103 -78324 -81059
rect -78268 -81103 -78224 -81059
rect -78168 -81103 -78124 -81059
rect -78068 -81103 -78024 -81059
rect -77968 -81103 -77924 -81059
rect -77868 -81103 -77824 -81059
rect -77768 -81103 -77724 -81059
rect -77668 -81103 -77624 -81059
rect -77568 -81103 -77524 -81059
rect -77468 -81103 -77424 -81059
rect -76968 -81103 -76924 -81059
rect -76868 -81103 -76824 -81059
rect -76768 -81103 -76724 -81059
rect -76668 -81103 -76624 -81059
rect -76568 -81103 -76524 -81059
rect -76468 -81103 -76424 -81059
rect -76368 -81103 -76324 -81059
rect -76268 -81103 -76224 -81059
rect -76168 -81103 -76124 -81059
rect -76068 -81103 -76024 -81059
rect -75968 -81103 -75924 -81059
rect -75868 -81103 -75824 -81059
rect -75768 -81103 -75724 -81059
rect -75668 -81103 -75624 -81059
rect -75568 -81103 -75524 -81059
rect -75468 -81103 -75424 -81059
rect -50017 -81105 -49973 -81061
rect -49917 -81105 -49873 -81061
rect -49817 -81105 -49773 -81061
rect -49717 -81105 -49673 -81061
rect -49617 -81105 -49573 -81061
rect -49517 -81105 -49473 -81061
rect -49417 -81105 -49373 -81061
rect -49317 -81105 -49273 -81061
rect -49217 -81105 -49173 -81061
rect -49117 -81105 -49073 -81061
rect -49017 -81105 -48973 -81061
rect -48917 -81105 -48873 -81061
rect -48817 -81105 -48773 -81061
rect -48717 -81105 -48673 -81061
rect -48617 -81105 -48573 -81061
rect -48517 -81105 -48473 -81061
rect -48017 -81105 -47973 -81061
rect -47917 -81105 -47873 -81061
rect -47817 -81105 -47773 -81061
rect -47717 -81105 -47673 -81061
rect -47617 -81105 -47573 -81061
rect -47517 -81105 -47473 -81061
rect -47417 -81105 -47373 -81061
rect -47317 -81105 -47273 -81061
rect -47217 -81105 -47173 -81061
rect -47117 -81105 -47073 -81061
rect -47017 -81105 -46973 -81061
rect -46917 -81105 -46873 -81061
rect -46817 -81105 -46773 -81061
rect -46717 -81105 -46673 -81061
rect -46617 -81105 -46573 -81061
rect -46517 -81105 -46473 -81061
rect -46017 -81105 -45973 -81061
rect -45917 -81105 -45873 -81061
rect -45817 -81105 -45773 -81061
rect -45717 -81105 -45673 -81061
rect -45617 -81105 -45573 -81061
rect -45517 -81105 -45473 -81061
rect -45417 -81105 -45373 -81061
rect -45317 -81105 -45273 -81061
rect -45217 -81105 -45173 -81061
rect -45117 -81105 -45073 -81061
rect -45017 -81105 -44973 -81061
rect -44917 -81105 -44873 -81061
rect -44817 -81105 -44773 -81061
rect -44717 -81105 -44673 -81061
rect -44617 -81105 -44573 -81061
rect -44517 -81105 -44473 -81061
rect -44017 -81105 -43973 -81061
rect -43917 -81105 -43873 -81061
rect -43817 -81105 -43773 -81061
rect -43717 -81105 -43673 -81061
rect -43617 -81105 -43573 -81061
rect -43517 -81105 -43473 -81061
rect -43417 -81105 -43373 -81061
rect -43317 -81105 -43273 -81061
rect -43217 -81105 -43173 -81061
rect -43117 -81105 -43073 -81061
rect -43017 -81105 -42973 -81061
rect -42917 -81105 -42873 -81061
rect -42817 -81105 -42773 -81061
rect -42717 -81105 -42673 -81061
rect -42617 -81105 -42573 -81061
rect -42517 -81105 -42473 -81061
rect 80737 -81099 80781 -81055
rect 80837 -81099 80881 -81055
rect 80937 -81099 80981 -81055
rect 81037 -81099 81081 -81055
rect 81137 -81099 81181 -81055
rect 81237 -81099 81281 -81055
rect 81337 -81099 81381 -81055
rect 81437 -81099 81481 -81055
rect 81537 -81099 81581 -81055
rect 81637 -81099 81681 -81055
rect 81737 -81099 81781 -81055
rect 81837 -81099 81881 -81055
rect 81937 -81099 81981 -81055
rect 82037 -81099 82081 -81055
rect 82137 -81099 82181 -81055
rect 82237 -81099 82281 -81055
rect 82737 -81099 82781 -81055
rect 82837 -81099 82881 -81055
rect 82937 -81099 82981 -81055
rect 83037 -81099 83081 -81055
rect 83137 -81099 83181 -81055
rect 83237 -81099 83281 -81055
rect 83337 -81099 83381 -81055
rect 83437 -81099 83481 -81055
rect 83537 -81099 83581 -81055
rect 83637 -81099 83681 -81055
rect 83737 -81099 83781 -81055
rect 83837 -81099 83881 -81055
rect 83937 -81099 83981 -81055
rect 84037 -81099 84081 -81055
rect 84137 -81099 84181 -81055
rect 84237 -81099 84281 -81055
rect 84737 -81099 84781 -81055
rect 84837 -81099 84881 -81055
rect 84937 -81099 84981 -81055
rect 85037 -81099 85081 -81055
rect 85137 -81099 85181 -81055
rect 85237 -81099 85281 -81055
rect 85337 -81099 85381 -81055
rect 85437 -81099 85481 -81055
rect 85537 -81099 85581 -81055
rect 85637 -81099 85681 -81055
rect 85737 -81099 85781 -81055
rect 85837 -81099 85881 -81055
rect 85937 -81099 85981 -81055
rect 86037 -81099 86081 -81055
rect 86137 -81099 86181 -81055
rect 86237 -81099 86281 -81055
rect 86737 -81099 86781 -81055
rect 86837 -81099 86881 -81055
rect 86937 -81099 86981 -81055
rect 87037 -81099 87081 -81055
rect 87137 -81099 87181 -81055
rect 87237 -81099 87281 -81055
rect 87337 -81099 87381 -81055
rect 87437 -81099 87481 -81055
rect 87537 -81099 87581 -81055
rect 87637 -81099 87681 -81055
rect 87737 -81099 87781 -81055
rect 87837 -81099 87881 -81055
rect 87937 -81099 87981 -81055
rect 88037 -81099 88081 -81055
rect 88137 -81099 88181 -81055
rect 88237 -81099 88281 -81055
rect -82968 -81203 -82924 -81159
rect -82868 -81203 -82824 -81159
rect -82768 -81203 -82724 -81159
rect -82668 -81203 -82624 -81159
rect -82568 -81203 -82524 -81159
rect -82468 -81203 -82424 -81159
rect -82368 -81203 -82324 -81159
rect -82268 -81203 -82224 -81159
rect -82168 -81203 -82124 -81159
rect -82068 -81203 -82024 -81159
rect -81968 -81203 -81924 -81159
rect -81868 -81203 -81824 -81159
rect -81768 -81203 -81724 -81159
rect -81668 -81203 -81624 -81159
rect -81568 -81203 -81524 -81159
rect -81468 -81203 -81424 -81159
rect -80968 -81203 -80924 -81159
rect -80868 -81203 -80824 -81159
rect -80768 -81203 -80724 -81159
rect -80668 -81203 -80624 -81159
rect -80568 -81203 -80524 -81159
rect -80468 -81203 -80424 -81159
rect -80368 -81203 -80324 -81159
rect -80268 -81203 -80224 -81159
rect -80168 -81203 -80124 -81159
rect -80068 -81203 -80024 -81159
rect -79968 -81203 -79924 -81159
rect -79868 -81203 -79824 -81159
rect -79768 -81203 -79724 -81159
rect -79668 -81203 -79624 -81159
rect -79568 -81203 -79524 -81159
rect -79468 -81203 -79424 -81159
rect -78968 -81203 -78924 -81159
rect -78868 -81203 -78824 -81159
rect -78768 -81203 -78724 -81159
rect -78668 -81203 -78624 -81159
rect -78568 -81203 -78524 -81159
rect -78468 -81203 -78424 -81159
rect -78368 -81203 -78324 -81159
rect -78268 -81203 -78224 -81159
rect -78168 -81203 -78124 -81159
rect -78068 -81203 -78024 -81159
rect -77968 -81203 -77924 -81159
rect -77868 -81203 -77824 -81159
rect -77768 -81203 -77724 -81159
rect -77668 -81203 -77624 -81159
rect -77568 -81203 -77524 -81159
rect -77468 -81203 -77424 -81159
rect -76968 -81203 -76924 -81159
rect -76868 -81203 -76824 -81159
rect -76768 -81203 -76724 -81159
rect -76668 -81203 -76624 -81159
rect -76568 -81203 -76524 -81159
rect -76468 -81203 -76424 -81159
rect -76368 -81203 -76324 -81159
rect -76268 -81203 -76224 -81159
rect -76168 -81203 -76124 -81159
rect -76068 -81203 -76024 -81159
rect -75968 -81203 -75924 -81159
rect -75868 -81203 -75824 -81159
rect -75768 -81203 -75724 -81159
rect -75668 -81203 -75624 -81159
rect -75568 -81203 -75524 -81159
rect -75468 -81203 -75424 -81159
rect -50017 -81205 -49973 -81161
rect -49917 -81205 -49873 -81161
rect -49817 -81205 -49773 -81161
rect -49717 -81205 -49673 -81161
rect -49617 -81205 -49573 -81161
rect -49517 -81205 -49473 -81161
rect -49417 -81205 -49373 -81161
rect -49317 -81205 -49273 -81161
rect -49217 -81205 -49173 -81161
rect -49117 -81205 -49073 -81161
rect -49017 -81205 -48973 -81161
rect -48917 -81205 -48873 -81161
rect -48817 -81205 -48773 -81161
rect -48717 -81205 -48673 -81161
rect -48617 -81205 -48573 -81161
rect -48517 -81205 -48473 -81161
rect -48017 -81205 -47973 -81161
rect -47917 -81205 -47873 -81161
rect -47817 -81205 -47773 -81161
rect -47717 -81205 -47673 -81161
rect -47617 -81205 -47573 -81161
rect -47517 -81205 -47473 -81161
rect -47417 -81205 -47373 -81161
rect -47317 -81205 -47273 -81161
rect -47217 -81205 -47173 -81161
rect -47117 -81205 -47073 -81161
rect -47017 -81205 -46973 -81161
rect -46917 -81205 -46873 -81161
rect -46817 -81205 -46773 -81161
rect -46717 -81205 -46673 -81161
rect -46617 -81205 -46573 -81161
rect -46517 -81205 -46473 -81161
rect -46017 -81205 -45973 -81161
rect -45917 -81205 -45873 -81161
rect -45817 -81205 -45773 -81161
rect -45717 -81205 -45673 -81161
rect -45617 -81205 -45573 -81161
rect -45517 -81205 -45473 -81161
rect -45417 -81205 -45373 -81161
rect -45317 -81205 -45273 -81161
rect -45217 -81205 -45173 -81161
rect -45117 -81205 -45073 -81161
rect -45017 -81205 -44973 -81161
rect -44917 -81205 -44873 -81161
rect -44817 -81205 -44773 -81161
rect -44717 -81205 -44673 -81161
rect -44617 -81205 -44573 -81161
rect -44517 -81205 -44473 -81161
rect -44017 -81205 -43973 -81161
rect -43917 -81205 -43873 -81161
rect -43817 -81205 -43773 -81161
rect -43717 -81205 -43673 -81161
rect -43617 -81205 -43573 -81161
rect -43517 -81205 -43473 -81161
rect -43417 -81205 -43373 -81161
rect -43317 -81205 -43273 -81161
rect -43217 -81205 -43173 -81161
rect -43117 -81205 -43073 -81161
rect -43017 -81205 -42973 -81161
rect -42917 -81205 -42873 -81161
rect -42817 -81205 -42773 -81161
rect -42717 -81205 -42673 -81161
rect -42617 -81205 -42573 -81161
rect -42517 -81205 -42473 -81161
rect 80737 -81199 80781 -81155
rect 80837 -81199 80881 -81155
rect 80937 -81199 80981 -81155
rect 81037 -81199 81081 -81155
rect 81137 -81199 81181 -81155
rect 81237 -81199 81281 -81155
rect 81337 -81199 81381 -81155
rect 81437 -81199 81481 -81155
rect 81537 -81199 81581 -81155
rect 81637 -81199 81681 -81155
rect 81737 -81199 81781 -81155
rect 81837 -81199 81881 -81155
rect 81937 -81199 81981 -81155
rect 82037 -81199 82081 -81155
rect 82137 -81199 82181 -81155
rect 82237 -81199 82281 -81155
rect 82737 -81199 82781 -81155
rect 82837 -81199 82881 -81155
rect 82937 -81199 82981 -81155
rect 83037 -81199 83081 -81155
rect 83137 -81199 83181 -81155
rect 83237 -81199 83281 -81155
rect 83337 -81199 83381 -81155
rect 83437 -81199 83481 -81155
rect 83537 -81199 83581 -81155
rect 83637 -81199 83681 -81155
rect 83737 -81199 83781 -81155
rect 83837 -81199 83881 -81155
rect 83937 -81199 83981 -81155
rect 84037 -81199 84081 -81155
rect 84137 -81199 84181 -81155
rect 84237 -81199 84281 -81155
rect 84737 -81199 84781 -81155
rect 84837 -81199 84881 -81155
rect 84937 -81199 84981 -81155
rect 85037 -81199 85081 -81155
rect 85137 -81199 85181 -81155
rect 85237 -81199 85281 -81155
rect 85337 -81199 85381 -81155
rect 85437 -81199 85481 -81155
rect 85537 -81199 85581 -81155
rect 85637 -81199 85681 -81155
rect 85737 -81199 85781 -81155
rect 85837 -81199 85881 -81155
rect 85937 -81199 85981 -81155
rect 86037 -81199 86081 -81155
rect 86137 -81199 86181 -81155
rect 86237 -81199 86281 -81155
rect 86737 -81199 86781 -81155
rect 86837 -81199 86881 -81155
rect 86937 -81199 86981 -81155
rect 87037 -81199 87081 -81155
rect 87137 -81199 87181 -81155
rect 87237 -81199 87281 -81155
rect 87337 -81199 87381 -81155
rect 87437 -81199 87481 -81155
rect 87537 -81199 87581 -81155
rect 87637 -81199 87681 -81155
rect 87737 -81199 87781 -81155
rect 87837 -81199 87881 -81155
rect 87937 -81199 87981 -81155
rect 88037 -81199 88081 -81155
rect 88137 -81199 88181 -81155
rect 88237 -81199 88281 -81155
rect -82968 -81303 -82924 -81259
rect -82868 -81303 -82824 -81259
rect -82768 -81303 -82724 -81259
rect -82668 -81303 -82624 -81259
rect -82568 -81303 -82524 -81259
rect -82468 -81303 -82424 -81259
rect -82368 -81303 -82324 -81259
rect -82268 -81303 -82224 -81259
rect -82168 -81303 -82124 -81259
rect -82068 -81303 -82024 -81259
rect -81968 -81303 -81924 -81259
rect -81868 -81303 -81824 -81259
rect -81768 -81303 -81724 -81259
rect -81668 -81303 -81624 -81259
rect -81568 -81303 -81524 -81259
rect -81468 -81303 -81424 -81259
rect -80968 -81303 -80924 -81259
rect -80868 -81303 -80824 -81259
rect -80768 -81303 -80724 -81259
rect -80668 -81303 -80624 -81259
rect -80568 -81303 -80524 -81259
rect -80468 -81303 -80424 -81259
rect -80368 -81303 -80324 -81259
rect -80268 -81303 -80224 -81259
rect -80168 -81303 -80124 -81259
rect -80068 -81303 -80024 -81259
rect -79968 -81303 -79924 -81259
rect -79868 -81303 -79824 -81259
rect -79768 -81303 -79724 -81259
rect -79668 -81303 -79624 -81259
rect -79568 -81303 -79524 -81259
rect -79468 -81303 -79424 -81259
rect -78968 -81303 -78924 -81259
rect -78868 -81303 -78824 -81259
rect -78768 -81303 -78724 -81259
rect -78668 -81303 -78624 -81259
rect -78568 -81303 -78524 -81259
rect -78468 -81303 -78424 -81259
rect -78368 -81303 -78324 -81259
rect -78268 -81303 -78224 -81259
rect -78168 -81303 -78124 -81259
rect -78068 -81303 -78024 -81259
rect -77968 -81303 -77924 -81259
rect -77868 -81303 -77824 -81259
rect -77768 -81303 -77724 -81259
rect -77668 -81303 -77624 -81259
rect -77568 -81303 -77524 -81259
rect -77468 -81303 -77424 -81259
rect -76968 -81303 -76924 -81259
rect -76868 -81303 -76824 -81259
rect -76768 -81303 -76724 -81259
rect -76668 -81303 -76624 -81259
rect -76568 -81303 -76524 -81259
rect -76468 -81303 -76424 -81259
rect -76368 -81303 -76324 -81259
rect -76268 -81303 -76224 -81259
rect -76168 -81303 -76124 -81259
rect -76068 -81303 -76024 -81259
rect -75968 -81303 -75924 -81259
rect -75868 -81303 -75824 -81259
rect -75768 -81303 -75724 -81259
rect -75668 -81303 -75624 -81259
rect -75568 -81303 -75524 -81259
rect -75468 -81303 -75424 -81259
rect -50017 -81305 -49973 -81261
rect -49917 -81305 -49873 -81261
rect -49817 -81305 -49773 -81261
rect -49717 -81305 -49673 -81261
rect -49617 -81305 -49573 -81261
rect -49517 -81305 -49473 -81261
rect -49417 -81305 -49373 -81261
rect -49317 -81305 -49273 -81261
rect -49217 -81305 -49173 -81261
rect -49117 -81305 -49073 -81261
rect -49017 -81305 -48973 -81261
rect -48917 -81305 -48873 -81261
rect -48817 -81305 -48773 -81261
rect -48717 -81305 -48673 -81261
rect -48617 -81305 -48573 -81261
rect -48517 -81305 -48473 -81261
rect -48017 -81305 -47973 -81261
rect -47917 -81305 -47873 -81261
rect -47817 -81305 -47773 -81261
rect -47717 -81305 -47673 -81261
rect -47617 -81305 -47573 -81261
rect -47517 -81305 -47473 -81261
rect -47417 -81305 -47373 -81261
rect -47317 -81305 -47273 -81261
rect -47217 -81305 -47173 -81261
rect -47117 -81305 -47073 -81261
rect -47017 -81305 -46973 -81261
rect -46917 -81305 -46873 -81261
rect -46817 -81305 -46773 -81261
rect -46717 -81305 -46673 -81261
rect -46617 -81305 -46573 -81261
rect -46517 -81305 -46473 -81261
rect -46017 -81305 -45973 -81261
rect -45917 -81305 -45873 -81261
rect -45817 -81305 -45773 -81261
rect -45717 -81305 -45673 -81261
rect -45617 -81305 -45573 -81261
rect -45517 -81305 -45473 -81261
rect -45417 -81305 -45373 -81261
rect -45317 -81305 -45273 -81261
rect -45217 -81305 -45173 -81261
rect -45117 -81305 -45073 -81261
rect -45017 -81305 -44973 -81261
rect -44917 -81305 -44873 -81261
rect -44817 -81305 -44773 -81261
rect -44717 -81305 -44673 -81261
rect -44617 -81305 -44573 -81261
rect -44517 -81305 -44473 -81261
rect -44017 -81305 -43973 -81261
rect -43917 -81305 -43873 -81261
rect -43817 -81305 -43773 -81261
rect -43717 -81305 -43673 -81261
rect -43617 -81305 -43573 -81261
rect -43517 -81305 -43473 -81261
rect -43417 -81305 -43373 -81261
rect -43317 -81305 -43273 -81261
rect -43217 -81305 -43173 -81261
rect -43117 -81305 -43073 -81261
rect -43017 -81305 -42973 -81261
rect -42917 -81305 -42873 -81261
rect -42817 -81305 -42773 -81261
rect -42717 -81305 -42673 -81261
rect -42617 -81305 -42573 -81261
rect -42517 -81305 -42473 -81261
rect 80737 -81299 80781 -81255
rect 80837 -81299 80881 -81255
rect 80937 -81299 80981 -81255
rect 81037 -81299 81081 -81255
rect 81137 -81299 81181 -81255
rect 81237 -81299 81281 -81255
rect 81337 -81299 81381 -81255
rect 81437 -81299 81481 -81255
rect 81537 -81299 81581 -81255
rect 81637 -81299 81681 -81255
rect 81737 -81299 81781 -81255
rect 81837 -81299 81881 -81255
rect 81937 -81299 81981 -81255
rect 82037 -81299 82081 -81255
rect 82137 -81299 82181 -81255
rect 82237 -81299 82281 -81255
rect 82737 -81299 82781 -81255
rect 82837 -81299 82881 -81255
rect 82937 -81299 82981 -81255
rect 83037 -81299 83081 -81255
rect 83137 -81299 83181 -81255
rect 83237 -81299 83281 -81255
rect 83337 -81299 83381 -81255
rect 83437 -81299 83481 -81255
rect 83537 -81299 83581 -81255
rect 83637 -81299 83681 -81255
rect 83737 -81299 83781 -81255
rect 83837 -81299 83881 -81255
rect 83937 -81299 83981 -81255
rect 84037 -81299 84081 -81255
rect 84137 -81299 84181 -81255
rect 84237 -81299 84281 -81255
rect 84737 -81299 84781 -81255
rect 84837 -81299 84881 -81255
rect 84937 -81299 84981 -81255
rect 85037 -81299 85081 -81255
rect 85137 -81299 85181 -81255
rect 85237 -81299 85281 -81255
rect 85337 -81299 85381 -81255
rect 85437 -81299 85481 -81255
rect 85537 -81299 85581 -81255
rect 85637 -81299 85681 -81255
rect 85737 -81299 85781 -81255
rect 85837 -81299 85881 -81255
rect 85937 -81299 85981 -81255
rect 86037 -81299 86081 -81255
rect 86137 -81299 86181 -81255
rect 86237 -81299 86281 -81255
rect 86737 -81299 86781 -81255
rect 86837 -81299 86881 -81255
rect 86937 -81299 86981 -81255
rect 87037 -81299 87081 -81255
rect 87137 -81299 87181 -81255
rect 87237 -81299 87281 -81255
rect 87337 -81299 87381 -81255
rect 87437 -81299 87481 -81255
rect 87537 -81299 87581 -81255
rect 87637 -81299 87681 -81255
rect 87737 -81299 87781 -81255
rect 87837 -81299 87881 -81255
rect 87937 -81299 87981 -81255
rect 88037 -81299 88081 -81255
rect 88137 -81299 88181 -81255
rect 88237 -81299 88281 -81255
rect -82968 -81403 -82924 -81359
rect -82868 -81403 -82824 -81359
rect -82768 -81403 -82724 -81359
rect -82668 -81403 -82624 -81359
rect -82568 -81403 -82524 -81359
rect -82468 -81403 -82424 -81359
rect -82368 -81403 -82324 -81359
rect -82268 -81403 -82224 -81359
rect -82168 -81403 -82124 -81359
rect -82068 -81403 -82024 -81359
rect -81968 -81403 -81924 -81359
rect -81868 -81403 -81824 -81359
rect -81768 -81403 -81724 -81359
rect -81668 -81403 -81624 -81359
rect -81568 -81403 -81524 -81359
rect -81468 -81403 -81424 -81359
rect -80968 -81403 -80924 -81359
rect -80868 -81403 -80824 -81359
rect -80768 -81403 -80724 -81359
rect -80668 -81403 -80624 -81359
rect -80568 -81403 -80524 -81359
rect -80468 -81403 -80424 -81359
rect -80368 -81403 -80324 -81359
rect -80268 -81403 -80224 -81359
rect -80168 -81403 -80124 -81359
rect -80068 -81403 -80024 -81359
rect -79968 -81403 -79924 -81359
rect -79868 -81403 -79824 -81359
rect -79768 -81403 -79724 -81359
rect -79668 -81403 -79624 -81359
rect -79568 -81403 -79524 -81359
rect -79468 -81403 -79424 -81359
rect -78968 -81403 -78924 -81359
rect -78868 -81403 -78824 -81359
rect -78768 -81403 -78724 -81359
rect -78668 -81403 -78624 -81359
rect -78568 -81403 -78524 -81359
rect -78468 -81403 -78424 -81359
rect -78368 -81403 -78324 -81359
rect -78268 -81403 -78224 -81359
rect -78168 -81403 -78124 -81359
rect -78068 -81403 -78024 -81359
rect -77968 -81403 -77924 -81359
rect -77868 -81403 -77824 -81359
rect -77768 -81403 -77724 -81359
rect -77668 -81403 -77624 -81359
rect -77568 -81403 -77524 -81359
rect -77468 -81403 -77424 -81359
rect -76968 -81403 -76924 -81359
rect -76868 -81403 -76824 -81359
rect -76768 -81403 -76724 -81359
rect -76668 -81403 -76624 -81359
rect -76568 -81403 -76524 -81359
rect -76468 -81403 -76424 -81359
rect -76368 -81403 -76324 -81359
rect -76268 -81403 -76224 -81359
rect -76168 -81403 -76124 -81359
rect -76068 -81403 -76024 -81359
rect -75968 -81403 -75924 -81359
rect -75868 -81403 -75824 -81359
rect -75768 -81403 -75724 -81359
rect -75668 -81403 -75624 -81359
rect -75568 -81403 -75524 -81359
rect -75468 -81403 -75424 -81359
rect -50017 -81405 -49973 -81361
rect -49917 -81405 -49873 -81361
rect -49817 -81405 -49773 -81361
rect -49717 -81405 -49673 -81361
rect -49617 -81405 -49573 -81361
rect -49517 -81405 -49473 -81361
rect -49417 -81405 -49373 -81361
rect -49317 -81405 -49273 -81361
rect -49217 -81405 -49173 -81361
rect -49117 -81405 -49073 -81361
rect -49017 -81405 -48973 -81361
rect -48917 -81405 -48873 -81361
rect -48817 -81405 -48773 -81361
rect -48717 -81405 -48673 -81361
rect -48617 -81405 -48573 -81361
rect -48517 -81405 -48473 -81361
rect -48017 -81405 -47973 -81361
rect -47917 -81405 -47873 -81361
rect -47817 -81405 -47773 -81361
rect -47717 -81405 -47673 -81361
rect -47617 -81405 -47573 -81361
rect -47517 -81405 -47473 -81361
rect -47417 -81405 -47373 -81361
rect -47317 -81405 -47273 -81361
rect -47217 -81405 -47173 -81361
rect -47117 -81405 -47073 -81361
rect -47017 -81405 -46973 -81361
rect -46917 -81405 -46873 -81361
rect -46817 -81405 -46773 -81361
rect -46717 -81405 -46673 -81361
rect -46617 -81405 -46573 -81361
rect -46517 -81405 -46473 -81361
rect -46017 -81405 -45973 -81361
rect -45917 -81405 -45873 -81361
rect -45817 -81405 -45773 -81361
rect -45717 -81405 -45673 -81361
rect -45617 -81405 -45573 -81361
rect -45517 -81405 -45473 -81361
rect -45417 -81405 -45373 -81361
rect -45317 -81405 -45273 -81361
rect -45217 -81405 -45173 -81361
rect -45117 -81405 -45073 -81361
rect -45017 -81405 -44973 -81361
rect -44917 -81405 -44873 -81361
rect -44817 -81405 -44773 -81361
rect -44717 -81405 -44673 -81361
rect -44617 -81405 -44573 -81361
rect -44517 -81405 -44473 -81361
rect -44017 -81405 -43973 -81361
rect -43917 -81405 -43873 -81361
rect -43817 -81405 -43773 -81361
rect -43717 -81405 -43673 -81361
rect -43617 -81405 -43573 -81361
rect -43517 -81405 -43473 -81361
rect -43417 -81405 -43373 -81361
rect -43317 -81405 -43273 -81361
rect -43217 -81405 -43173 -81361
rect -43117 -81405 -43073 -81361
rect -43017 -81405 -42973 -81361
rect -42917 -81405 -42873 -81361
rect -42817 -81405 -42773 -81361
rect -42717 -81405 -42673 -81361
rect -42617 -81405 -42573 -81361
rect -42517 -81405 -42473 -81361
rect 80737 -81399 80781 -81355
rect 80837 -81399 80881 -81355
rect 80937 -81399 80981 -81355
rect 81037 -81399 81081 -81355
rect 81137 -81399 81181 -81355
rect 81237 -81399 81281 -81355
rect 81337 -81399 81381 -81355
rect 81437 -81399 81481 -81355
rect 81537 -81399 81581 -81355
rect 81637 -81399 81681 -81355
rect 81737 -81399 81781 -81355
rect 81837 -81399 81881 -81355
rect 81937 -81399 81981 -81355
rect 82037 -81399 82081 -81355
rect 82137 -81399 82181 -81355
rect 82237 -81399 82281 -81355
rect 82737 -81399 82781 -81355
rect 82837 -81399 82881 -81355
rect 82937 -81399 82981 -81355
rect 83037 -81399 83081 -81355
rect 83137 -81399 83181 -81355
rect 83237 -81399 83281 -81355
rect 83337 -81399 83381 -81355
rect 83437 -81399 83481 -81355
rect 83537 -81399 83581 -81355
rect 83637 -81399 83681 -81355
rect 83737 -81399 83781 -81355
rect 83837 -81399 83881 -81355
rect 83937 -81399 83981 -81355
rect 84037 -81399 84081 -81355
rect 84137 -81399 84181 -81355
rect 84237 -81399 84281 -81355
rect 84737 -81399 84781 -81355
rect 84837 -81399 84881 -81355
rect 84937 -81399 84981 -81355
rect 85037 -81399 85081 -81355
rect 85137 -81399 85181 -81355
rect 85237 -81399 85281 -81355
rect 85337 -81399 85381 -81355
rect 85437 -81399 85481 -81355
rect 85537 -81399 85581 -81355
rect 85637 -81399 85681 -81355
rect 85737 -81399 85781 -81355
rect 85837 -81399 85881 -81355
rect 85937 -81399 85981 -81355
rect 86037 -81399 86081 -81355
rect 86137 -81399 86181 -81355
rect 86237 -81399 86281 -81355
rect 86737 -81399 86781 -81355
rect 86837 -81399 86881 -81355
rect 86937 -81399 86981 -81355
rect 87037 -81399 87081 -81355
rect 87137 -81399 87181 -81355
rect 87237 -81399 87281 -81355
rect 87337 -81399 87381 -81355
rect 87437 -81399 87481 -81355
rect 87537 -81399 87581 -81355
rect 87637 -81399 87681 -81355
rect 87737 -81399 87781 -81355
rect 87837 -81399 87881 -81355
rect 87937 -81399 87981 -81355
rect 88037 -81399 88081 -81355
rect 88137 -81399 88181 -81355
rect 88237 -81399 88281 -81355
rect -82968 -81503 -82924 -81459
rect -82868 -81503 -82824 -81459
rect -82768 -81503 -82724 -81459
rect -82668 -81503 -82624 -81459
rect -82568 -81503 -82524 -81459
rect -82468 -81503 -82424 -81459
rect -82368 -81503 -82324 -81459
rect -82268 -81503 -82224 -81459
rect -82168 -81503 -82124 -81459
rect -82068 -81503 -82024 -81459
rect -81968 -81503 -81924 -81459
rect -81868 -81503 -81824 -81459
rect -81768 -81503 -81724 -81459
rect -81668 -81503 -81624 -81459
rect -81568 -81503 -81524 -81459
rect -81468 -81503 -81424 -81459
rect -80968 -81503 -80924 -81459
rect -80868 -81503 -80824 -81459
rect -80768 -81503 -80724 -81459
rect -80668 -81503 -80624 -81459
rect -80568 -81503 -80524 -81459
rect -80468 -81503 -80424 -81459
rect -80368 -81503 -80324 -81459
rect -80268 -81503 -80224 -81459
rect -80168 -81503 -80124 -81459
rect -80068 -81503 -80024 -81459
rect -79968 -81503 -79924 -81459
rect -79868 -81503 -79824 -81459
rect -79768 -81503 -79724 -81459
rect -79668 -81503 -79624 -81459
rect -79568 -81503 -79524 -81459
rect -79468 -81503 -79424 -81459
rect -78968 -81503 -78924 -81459
rect -78868 -81503 -78824 -81459
rect -78768 -81503 -78724 -81459
rect -78668 -81503 -78624 -81459
rect -78568 -81503 -78524 -81459
rect -78468 -81503 -78424 -81459
rect -78368 -81503 -78324 -81459
rect -78268 -81503 -78224 -81459
rect -78168 -81503 -78124 -81459
rect -78068 -81503 -78024 -81459
rect -77968 -81503 -77924 -81459
rect -77868 -81503 -77824 -81459
rect -77768 -81503 -77724 -81459
rect -77668 -81503 -77624 -81459
rect -77568 -81503 -77524 -81459
rect -77468 -81503 -77424 -81459
rect -76968 -81503 -76924 -81459
rect -76868 -81503 -76824 -81459
rect -76768 -81503 -76724 -81459
rect -76668 -81503 -76624 -81459
rect -76568 -81503 -76524 -81459
rect -76468 -81503 -76424 -81459
rect -76368 -81503 -76324 -81459
rect -76268 -81503 -76224 -81459
rect -76168 -81503 -76124 -81459
rect -76068 -81503 -76024 -81459
rect -75968 -81503 -75924 -81459
rect -75868 -81503 -75824 -81459
rect -75768 -81503 -75724 -81459
rect -75668 -81503 -75624 -81459
rect -75568 -81503 -75524 -81459
rect -75468 -81503 -75424 -81459
rect -50017 -81505 -49973 -81461
rect -49917 -81505 -49873 -81461
rect -49817 -81505 -49773 -81461
rect -49717 -81505 -49673 -81461
rect -49617 -81505 -49573 -81461
rect -49517 -81505 -49473 -81461
rect -49417 -81505 -49373 -81461
rect -49317 -81505 -49273 -81461
rect -49217 -81505 -49173 -81461
rect -49117 -81505 -49073 -81461
rect -49017 -81505 -48973 -81461
rect -48917 -81505 -48873 -81461
rect -48817 -81505 -48773 -81461
rect -48717 -81505 -48673 -81461
rect -48617 -81505 -48573 -81461
rect -48517 -81505 -48473 -81461
rect -48017 -81505 -47973 -81461
rect -47917 -81505 -47873 -81461
rect -47817 -81505 -47773 -81461
rect -47717 -81505 -47673 -81461
rect -47617 -81505 -47573 -81461
rect -47517 -81505 -47473 -81461
rect -47417 -81505 -47373 -81461
rect -47317 -81505 -47273 -81461
rect -47217 -81505 -47173 -81461
rect -47117 -81505 -47073 -81461
rect -47017 -81505 -46973 -81461
rect -46917 -81505 -46873 -81461
rect -46817 -81505 -46773 -81461
rect -46717 -81505 -46673 -81461
rect -46617 -81505 -46573 -81461
rect -46517 -81505 -46473 -81461
rect -46017 -81505 -45973 -81461
rect -45917 -81505 -45873 -81461
rect -45817 -81505 -45773 -81461
rect -45717 -81505 -45673 -81461
rect -45617 -81505 -45573 -81461
rect -45517 -81505 -45473 -81461
rect -45417 -81505 -45373 -81461
rect -45317 -81505 -45273 -81461
rect -45217 -81505 -45173 -81461
rect -45117 -81505 -45073 -81461
rect -45017 -81505 -44973 -81461
rect -44917 -81505 -44873 -81461
rect -44817 -81505 -44773 -81461
rect -44717 -81505 -44673 -81461
rect -44617 -81505 -44573 -81461
rect -44517 -81505 -44473 -81461
rect -44017 -81505 -43973 -81461
rect -43917 -81505 -43873 -81461
rect -43817 -81505 -43773 -81461
rect -43717 -81505 -43673 -81461
rect -43617 -81505 -43573 -81461
rect -43517 -81505 -43473 -81461
rect -43417 -81505 -43373 -81461
rect -43317 -81505 -43273 -81461
rect -43217 -81505 -43173 -81461
rect -43117 -81505 -43073 -81461
rect -43017 -81505 -42973 -81461
rect -42917 -81505 -42873 -81461
rect -42817 -81505 -42773 -81461
rect -42717 -81505 -42673 -81461
rect -42617 -81505 -42573 -81461
rect -42517 -81505 -42473 -81461
rect 80737 -81499 80781 -81455
rect 80837 -81499 80881 -81455
rect 80937 -81499 80981 -81455
rect 81037 -81499 81081 -81455
rect 81137 -81499 81181 -81455
rect 81237 -81499 81281 -81455
rect 81337 -81499 81381 -81455
rect 81437 -81499 81481 -81455
rect 81537 -81499 81581 -81455
rect 81637 -81499 81681 -81455
rect 81737 -81499 81781 -81455
rect 81837 -81499 81881 -81455
rect 81937 -81499 81981 -81455
rect 82037 -81499 82081 -81455
rect 82137 -81499 82181 -81455
rect 82237 -81499 82281 -81455
rect 82737 -81499 82781 -81455
rect 82837 -81499 82881 -81455
rect 82937 -81499 82981 -81455
rect 83037 -81499 83081 -81455
rect 83137 -81499 83181 -81455
rect 83237 -81499 83281 -81455
rect 83337 -81499 83381 -81455
rect 83437 -81499 83481 -81455
rect 83537 -81499 83581 -81455
rect 83637 -81499 83681 -81455
rect 83737 -81499 83781 -81455
rect 83837 -81499 83881 -81455
rect 83937 -81499 83981 -81455
rect 84037 -81499 84081 -81455
rect 84137 -81499 84181 -81455
rect 84237 -81499 84281 -81455
rect 84737 -81499 84781 -81455
rect 84837 -81499 84881 -81455
rect 84937 -81499 84981 -81455
rect 85037 -81499 85081 -81455
rect 85137 -81499 85181 -81455
rect 85237 -81499 85281 -81455
rect 85337 -81499 85381 -81455
rect 85437 -81499 85481 -81455
rect 85537 -81499 85581 -81455
rect 85637 -81499 85681 -81455
rect 85737 -81499 85781 -81455
rect 85837 -81499 85881 -81455
rect 85937 -81499 85981 -81455
rect 86037 -81499 86081 -81455
rect 86137 -81499 86181 -81455
rect 86237 -81499 86281 -81455
rect 86737 -81499 86781 -81455
rect 86837 -81499 86881 -81455
rect 86937 -81499 86981 -81455
rect 87037 -81499 87081 -81455
rect 87137 -81499 87181 -81455
rect 87237 -81499 87281 -81455
rect 87337 -81499 87381 -81455
rect 87437 -81499 87481 -81455
rect 87537 -81499 87581 -81455
rect 87637 -81499 87681 -81455
rect 87737 -81499 87781 -81455
rect 87837 -81499 87881 -81455
rect 87937 -81499 87981 -81455
rect 88037 -81499 88081 -81455
rect 88137 -81499 88181 -81455
rect 88237 -81499 88281 -81455
rect -82968 -81603 -82924 -81559
rect -82868 -81603 -82824 -81559
rect -82768 -81603 -82724 -81559
rect -82668 -81603 -82624 -81559
rect -82568 -81603 -82524 -81559
rect -82468 -81603 -82424 -81559
rect -82368 -81603 -82324 -81559
rect -82268 -81603 -82224 -81559
rect -82168 -81603 -82124 -81559
rect -82068 -81603 -82024 -81559
rect -81968 -81603 -81924 -81559
rect -81868 -81603 -81824 -81559
rect -81768 -81603 -81724 -81559
rect -81668 -81603 -81624 -81559
rect -81568 -81603 -81524 -81559
rect -81468 -81603 -81424 -81559
rect -80968 -81603 -80924 -81559
rect -80868 -81603 -80824 -81559
rect -80768 -81603 -80724 -81559
rect -80668 -81603 -80624 -81559
rect -80568 -81603 -80524 -81559
rect -80468 -81603 -80424 -81559
rect -80368 -81603 -80324 -81559
rect -80268 -81603 -80224 -81559
rect -80168 -81603 -80124 -81559
rect -80068 -81603 -80024 -81559
rect -79968 -81603 -79924 -81559
rect -79868 -81603 -79824 -81559
rect -79768 -81603 -79724 -81559
rect -79668 -81603 -79624 -81559
rect -79568 -81603 -79524 -81559
rect -79468 -81603 -79424 -81559
rect -78968 -81603 -78924 -81559
rect -78868 -81603 -78824 -81559
rect -78768 -81603 -78724 -81559
rect -78668 -81603 -78624 -81559
rect -78568 -81603 -78524 -81559
rect -78468 -81603 -78424 -81559
rect -78368 -81603 -78324 -81559
rect -78268 -81603 -78224 -81559
rect -78168 -81603 -78124 -81559
rect -78068 -81603 -78024 -81559
rect -77968 -81603 -77924 -81559
rect -77868 -81603 -77824 -81559
rect -77768 -81603 -77724 -81559
rect -77668 -81603 -77624 -81559
rect -77568 -81603 -77524 -81559
rect -77468 -81603 -77424 -81559
rect -76968 -81603 -76924 -81559
rect -76868 -81603 -76824 -81559
rect -76768 -81603 -76724 -81559
rect -76668 -81603 -76624 -81559
rect -76568 -81603 -76524 -81559
rect -76468 -81603 -76424 -81559
rect -76368 -81603 -76324 -81559
rect -76268 -81603 -76224 -81559
rect -76168 -81603 -76124 -81559
rect -76068 -81603 -76024 -81559
rect -75968 -81603 -75924 -81559
rect -75868 -81603 -75824 -81559
rect -75768 -81603 -75724 -81559
rect -75668 -81603 -75624 -81559
rect -75568 -81603 -75524 -81559
rect -75468 -81603 -75424 -81559
rect -50017 -81605 -49973 -81561
rect -49917 -81605 -49873 -81561
rect -49817 -81605 -49773 -81561
rect -49717 -81605 -49673 -81561
rect -49617 -81605 -49573 -81561
rect -49517 -81605 -49473 -81561
rect -49417 -81605 -49373 -81561
rect -49317 -81605 -49273 -81561
rect -49217 -81605 -49173 -81561
rect -49117 -81605 -49073 -81561
rect -49017 -81605 -48973 -81561
rect -48917 -81605 -48873 -81561
rect -48817 -81605 -48773 -81561
rect -48717 -81605 -48673 -81561
rect -48617 -81605 -48573 -81561
rect -48517 -81605 -48473 -81561
rect -48017 -81605 -47973 -81561
rect -47917 -81605 -47873 -81561
rect -47817 -81605 -47773 -81561
rect -47717 -81605 -47673 -81561
rect -47617 -81605 -47573 -81561
rect -47517 -81605 -47473 -81561
rect -47417 -81605 -47373 -81561
rect -47317 -81605 -47273 -81561
rect -47217 -81605 -47173 -81561
rect -47117 -81605 -47073 -81561
rect -47017 -81605 -46973 -81561
rect -46917 -81605 -46873 -81561
rect -46817 -81605 -46773 -81561
rect -46717 -81605 -46673 -81561
rect -46617 -81605 -46573 -81561
rect -46517 -81605 -46473 -81561
rect -46017 -81605 -45973 -81561
rect -45917 -81605 -45873 -81561
rect -45817 -81605 -45773 -81561
rect -45717 -81605 -45673 -81561
rect -45617 -81605 -45573 -81561
rect -45517 -81605 -45473 -81561
rect -45417 -81605 -45373 -81561
rect -45317 -81605 -45273 -81561
rect -45217 -81605 -45173 -81561
rect -45117 -81605 -45073 -81561
rect -45017 -81605 -44973 -81561
rect -44917 -81605 -44873 -81561
rect -44817 -81605 -44773 -81561
rect -44717 -81605 -44673 -81561
rect -44617 -81605 -44573 -81561
rect -44517 -81605 -44473 -81561
rect -44017 -81605 -43973 -81561
rect -43917 -81605 -43873 -81561
rect -43817 -81605 -43773 -81561
rect -43717 -81605 -43673 -81561
rect -43617 -81605 -43573 -81561
rect -43517 -81605 -43473 -81561
rect -43417 -81605 -43373 -81561
rect -43317 -81605 -43273 -81561
rect -43217 -81605 -43173 -81561
rect -43117 -81605 -43073 -81561
rect -43017 -81605 -42973 -81561
rect -42917 -81605 -42873 -81561
rect -42817 -81605 -42773 -81561
rect -42717 -81605 -42673 -81561
rect -42617 -81605 -42573 -81561
rect -42517 -81605 -42473 -81561
rect 80737 -81599 80781 -81555
rect 80837 -81599 80881 -81555
rect 80937 -81599 80981 -81555
rect 81037 -81599 81081 -81555
rect 81137 -81599 81181 -81555
rect 81237 -81599 81281 -81555
rect 81337 -81599 81381 -81555
rect 81437 -81599 81481 -81555
rect 81537 -81599 81581 -81555
rect 81637 -81599 81681 -81555
rect 81737 -81599 81781 -81555
rect 81837 -81599 81881 -81555
rect 81937 -81599 81981 -81555
rect 82037 -81599 82081 -81555
rect 82137 -81599 82181 -81555
rect 82237 -81599 82281 -81555
rect 82737 -81599 82781 -81555
rect 82837 -81599 82881 -81555
rect 82937 -81599 82981 -81555
rect 83037 -81599 83081 -81555
rect 83137 -81599 83181 -81555
rect 83237 -81599 83281 -81555
rect 83337 -81599 83381 -81555
rect 83437 -81599 83481 -81555
rect 83537 -81599 83581 -81555
rect 83637 -81599 83681 -81555
rect 83737 -81599 83781 -81555
rect 83837 -81599 83881 -81555
rect 83937 -81599 83981 -81555
rect 84037 -81599 84081 -81555
rect 84137 -81599 84181 -81555
rect 84237 -81599 84281 -81555
rect 84737 -81599 84781 -81555
rect 84837 -81599 84881 -81555
rect 84937 -81599 84981 -81555
rect 85037 -81599 85081 -81555
rect 85137 -81599 85181 -81555
rect 85237 -81599 85281 -81555
rect 85337 -81599 85381 -81555
rect 85437 -81599 85481 -81555
rect 85537 -81599 85581 -81555
rect 85637 -81599 85681 -81555
rect 85737 -81599 85781 -81555
rect 85837 -81599 85881 -81555
rect 85937 -81599 85981 -81555
rect 86037 -81599 86081 -81555
rect 86137 -81599 86181 -81555
rect 86237 -81599 86281 -81555
rect 86737 -81599 86781 -81555
rect 86837 -81599 86881 -81555
rect 86937 -81599 86981 -81555
rect 87037 -81599 87081 -81555
rect 87137 -81599 87181 -81555
rect 87237 -81599 87281 -81555
rect 87337 -81599 87381 -81555
rect 87437 -81599 87481 -81555
rect 87537 -81599 87581 -81555
rect 87637 -81599 87681 -81555
rect 87737 -81599 87781 -81555
rect 87837 -81599 87881 -81555
rect 87937 -81599 87981 -81555
rect 88037 -81599 88081 -81555
rect 88137 -81599 88181 -81555
rect 88237 -81599 88281 -81555
rect -82968 -81703 -82924 -81659
rect -82868 -81703 -82824 -81659
rect -82768 -81703 -82724 -81659
rect -82668 -81703 -82624 -81659
rect -82568 -81703 -82524 -81659
rect -82468 -81703 -82424 -81659
rect -82368 -81703 -82324 -81659
rect -82268 -81703 -82224 -81659
rect -82168 -81703 -82124 -81659
rect -82068 -81703 -82024 -81659
rect -81968 -81703 -81924 -81659
rect -81868 -81703 -81824 -81659
rect -81768 -81703 -81724 -81659
rect -81668 -81703 -81624 -81659
rect -81568 -81703 -81524 -81659
rect -81468 -81703 -81424 -81659
rect -80968 -81703 -80924 -81659
rect -80868 -81703 -80824 -81659
rect -80768 -81703 -80724 -81659
rect -80668 -81703 -80624 -81659
rect -80568 -81703 -80524 -81659
rect -80468 -81703 -80424 -81659
rect -80368 -81703 -80324 -81659
rect -80268 -81703 -80224 -81659
rect -80168 -81703 -80124 -81659
rect -80068 -81703 -80024 -81659
rect -79968 -81703 -79924 -81659
rect -79868 -81703 -79824 -81659
rect -79768 -81703 -79724 -81659
rect -79668 -81703 -79624 -81659
rect -79568 -81703 -79524 -81659
rect -79468 -81703 -79424 -81659
rect -78968 -81703 -78924 -81659
rect -78868 -81703 -78824 -81659
rect -78768 -81703 -78724 -81659
rect -78668 -81703 -78624 -81659
rect -78568 -81703 -78524 -81659
rect -78468 -81703 -78424 -81659
rect -78368 -81703 -78324 -81659
rect -78268 -81703 -78224 -81659
rect -78168 -81703 -78124 -81659
rect -78068 -81703 -78024 -81659
rect -77968 -81703 -77924 -81659
rect -77868 -81703 -77824 -81659
rect -77768 -81703 -77724 -81659
rect -77668 -81703 -77624 -81659
rect -77568 -81703 -77524 -81659
rect -77468 -81703 -77424 -81659
rect -76968 -81703 -76924 -81659
rect -76868 -81703 -76824 -81659
rect -76768 -81703 -76724 -81659
rect -76668 -81703 -76624 -81659
rect -76568 -81703 -76524 -81659
rect -76468 -81703 -76424 -81659
rect -76368 -81703 -76324 -81659
rect -76268 -81703 -76224 -81659
rect -76168 -81703 -76124 -81659
rect -76068 -81703 -76024 -81659
rect -75968 -81703 -75924 -81659
rect -75868 -81703 -75824 -81659
rect -75768 -81703 -75724 -81659
rect -75668 -81703 -75624 -81659
rect -75568 -81703 -75524 -81659
rect -75468 -81703 -75424 -81659
rect -50017 -81705 -49973 -81661
rect -49917 -81705 -49873 -81661
rect -49817 -81705 -49773 -81661
rect -49717 -81705 -49673 -81661
rect -49617 -81705 -49573 -81661
rect -49517 -81705 -49473 -81661
rect -49417 -81705 -49373 -81661
rect -49317 -81705 -49273 -81661
rect -49217 -81705 -49173 -81661
rect -49117 -81705 -49073 -81661
rect -49017 -81705 -48973 -81661
rect -48917 -81705 -48873 -81661
rect -48817 -81705 -48773 -81661
rect -48717 -81705 -48673 -81661
rect -48617 -81705 -48573 -81661
rect -48517 -81705 -48473 -81661
rect -48017 -81705 -47973 -81661
rect -47917 -81705 -47873 -81661
rect -47817 -81705 -47773 -81661
rect -47717 -81705 -47673 -81661
rect -47617 -81705 -47573 -81661
rect -47517 -81705 -47473 -81661
rect -47417 -81705 -47373 -81661
rect -47317 -81705 -47273 -81661
rect -47217 -81705 -47173 -81661
rect -47117 -81705 -47073 -81661
rect -47017 -81705 -46973 -81661
rect -46917 -81705 -46873 -81661
rect -46817 -81705 -46773 -81661
rect -46717 -81705 -46673 -81661
rect -46617 -81705 -46573 -81661
rect -46517 -81705 -46473 -81661
rect -46017 -81705 -45973 -81661
rect -45917 -81705 -45873 -81661
rect -45817 -81705 -45773 -81661
rect -45717 -81705 -45673 -81661
rect -45617 -81705 -45573 -81661
rect -45517 -81705 -45473 -81661
rect -45417 -81705 -45373 -81661
rect -45317 -81705 -45273 -81661
rect -45217 -81705 -45173 -81661
rect -45117 -81705 -45073 -81661
rect -45017 -81705 -44973 -81661
rect -44917 -81705 -44873 -81661
rect -44817 -81705 -44773 -81661
rect -44717 -81705 -44673 -81661
rect -44617 -81705 -44573 -81661
rect -44517 -81705 -44473 -81661
rect -44017 -81705 -43973 -81661
rect -43917 -81705 -43873 -81661
rect -43817 -81705 -43773 -81661
rect -43717 -81705 -43673 -81661
rect -43617 -81705 -43573 -81661
rect -43517 -81705 -43473 -81661
rect -43417 -81705 -43373 -81661
rect -43317 -81705 -43273 -81661
rect -43217 -81705 -43173 -81661
rect -43117 -81705 -43073 -81661
rect -43017 -81705 -42973 -81661
rect -42917 -81705 -42873 -81661
rect -42817 -81705 -42773 -81661
rect -42717 -81705 -42673 -81661
rect -42617 -81705 -42573 -81661
rect -42517 -81705 -42473 -81661
rect 80737 -81699 80781 -81655
rect 80837 -81699 80881 -81655
rect 80937 -81699 80981 -81655
rect 81037 -81699 81081 -81655
rect 81137 -81699 81181 -81655
rect 81237 -81699 81281 -81655
rect 81337 -81699 81381 -81655
rect 81437 -81699 81481 -81655
rect 81537 -81699 81581 -81655
rect 81637 -81699 81681 -81655
rect 81737 -81699 81781 -81655
rect 81837 -81699 81881 -81655
rect 81937 -81699 81981 -81655
rect 82037 -81699 82081 -81655
rect 82137 -81699 82181 -81655
rect 82237 -81699 82281 -81655
rect 82737 -81699 82781 -81655
rect 82837 -81699 82881 -81655
rect 82937 -81699 82981 -81655
rect 83037 -81699 83081 -81655
rect 83137 -81699 83181 -81655
rect 83237 -81699 83281 -81655
rect 83337 -81699 83381 -81655
rect 83437 -81699 83481 -81655
rect 83537 -81699 83581 -81655
rect 83637 -81699 83681 -81655
rect 83737 -81699 83781 -81655
rect 83837 -81699 83881 -81655
rect 83937 -81699 83981 -81655
rect 84037 -81699 84081 -81655
rect 84137 -81699 84181 -81655
rect 84237 -81699 84281 -81655
rect 84737 -81699 84781 -81655
rect 84837 -81699 84881 -81655
rect 84937 -81699 84981 -81655
rect 85037 -81699 85081 -81655
rect 85137 -81699 85181 -81655
rect 85237 -81699 85281 -81655
rect 85337 -81699 85381 -81655
rect 85437 -81699 85481 -81655
rect 85537 -81699 85581 -81655
rect 85637 -81699 85681 -81655
rect 85737 -81699 85781 -81655
rect 85837 -81699 85881 -81655
rect 85937 -81699 85981 -81655
rect 86037 -81699 86081 -81655
rect 86137 -81699 86181 -81655
rect 86237 -81699 86281 -81655
rect 86737 -81699 86781 -81655
rect 86837 -81699 86881 -81655
rect 86937 -81699 86981 -81655
rect 87037 -81699 87081 -81655
rect 87137 -81699 87181 -81655
rect 87237 -81699 87281 -81655
rect 87337 -81699 87381 -81655
rect 87437 -81699 87481 -81655
rect 87537 -81699 87581 -81655
rect 87637 -81699 87681 -81655
rect 87737 -81699 87781 -81655
rect 87837 -81699 87881 -81655
rect 87937 -81699 87981 -81655
rect 88037 -81699 88081 -81655
rect 88137 -81699 88181 -81655
rect 88237 -81699 88281 -81655
rect -82968 -81803 -82924 -81759
rect -82868 -81803 -82824 -81759
rect -82768 -81803 -82724 -81759
rect -82668 -81803 -82624 -81759
rect -82568 -81803 -82524 -81759
rect -82468 -81803 -82424 -81759
rect -82368 -81803 -82324 -81759
rect -82268 -81803 -82224 -81759
rect -82168 -81803 -82124 -81759
rect -82068 -81803 -82024 -81759
rect -81968 -81803 -81924 -81759
rect -81868 -81803 -81824 -81759
rect -81768 -81803 -81724 -81759
rect -81668 -81803 -81624 -81759
rect -81568 -81803 -81524 -81759
rect -81468 -81803 -81424 -81759
rect -80968 -81803 -80924 -81759
rect -80868 -81803 -80824 -81759
rect -80768 -81803 -80724 -81759
rect -80668 -81803 -80624 -81759
rect -80568 -81803 -80524 -81759
rect -80468 -81803 -80424 -81759
rect -80368 -81803 -80324 -81759
rect -80268 -81803 -80224 -81759
rect -80168 -81803 -80124 -81759
rect -80068 -81803 -80024 -81759
rect -79968 -81803 -79924 -81759
rect -79868 -81803 -79824 -81759
rect -79768 -81803 -79724 -81759
rect -79668 -81803 -79624 -81759
rect -79568 -81803 -79524 -81759
rect -79468 -81803 -79424 -81759
rect -78968 -81803 -78924 -81759
rect -78868 -81803 -78824 -81759
rect -78768 -81803 -78724 -81759
rect -78668 -81803 -78624 -81759
rect -78568 -81803 -78524 -81759
rect -78468 -81803 -78424 -81759
rect -78368 -81803 -78324 -81759
rect -78268 -81803 -78224 -81759
rect -78168 -81803 -78124 -81759
rect -78068 -81803 -78024 -81759
rect -77968 -81803 -77924 -81759
rect -77868 -81803 -77824 -81759
rect -77768 -81803 -77724 -81759
rect -77668 -81803 -77624 -81759
rect -77568 -81803 -77524 -81759
rect -77468 -81803 -77424 -81759
rect -76968 -81803 -76924 -81759
rect -76868 -81803 -76824 -81759
rect -76768 -81803 -76724 -81759
rect -76668 -81803 -76624 -81759
rect -76568 -81803 -76524 -81759
rect -76468 -81803 -76424 -81759
rect -76368 -81803 -76324 -81759
rect -76268 -81803 -76224 -81759
rect -76168 -81803 -76124 -81759
rect -76068 -81803 -76024 -81759
rect -75968 -81803 -75924 -81759
rect -75868 -81803 -75824 -81759
rect -75768 -81803 -75724 -81759
rect -75668 -81803 -75624 -81759
rect -75568 -81803 -75524 -81759
rect -75468 -81803 -75424 -81759
rect -50017 -81805 -49973 -81761
rect -49917 -81805 -49873 -81761
rect -49817 -81805 -49773 -81761
rect -49717 -81805 -49673 -81761
rect -49617 -81805 -49573 -81761
rect -49517 -81805 -49473 -81761
rect -49417 -81805 -49373 -81761
rect -49317 -81805 -49273 -81761
rect -49217 -81805 -49173 -81761
rect -49117 -81805 -49073 -81761
rect -49017 -81805 -48973 -81761
rect -48917 -81805 -48873 -81761
rect -48817 -81805 -48773 -81761
rect -48717 -81805 -48673 -81761
rect -48617 -81805 -48573 -81761
rect -48517 -81805 -48473 -81761
rect -48017 -81805 -47973 -81761
rect -47917 -81805 -47873 -81761
rect -47817 -81805 -47773 -81761
rect -47717 -81805 -47673 -81761
rect -47617 -81805 -47573 -81761
rect -47517 -81805 -47473 -81761
rect -47417 -81805 -47373 -81761
rect -47317 -81805 -47273 -81761
rect -47217 -81805 -47173 -81761
rect -47117 -81805 -47073 -81761
rect -47017 -81805 -46973 -81761
rect -46917 -81805 -46873 -81761
rect -46817 -81805 -46773 -81761
rect -46717 -81805 -46673 -81761
rect -46617 -81805 -46573 -81761
rect -46517 -81805 -46473 -81761
rect -46017 -81805 -45973 -81761
rect -45917 -81805 -45873 -81761
rect -45817 -81805 -45773 -81761
rect -45717 -81805 -45673 -81761
rect -45617 -81805 -45573 -81761
rect -45517 -81805 -45473 -81761
rect -45417 -81805 -45373 -81761
rect -45317 -81805 -45273 -81761
rect -45217 -81805 -45173 -81761
rect -45117 -81805 -45073 -81761
rect -45017 -81805 -44973 -81761
rect -44917 -81805 -44873 -81761
rect -44817 -81805 -44773 -81761
rect -44717 -81805 -44673 -81761
rect -44617 -81805 -44573 -81761
rect -44517 -81805 -44473 -81761
rect -44017 -81805 -43973 -81761
rect -43917 -81805 -43873 -81761
rect -43817 -81805 -43773 -81761
rect -43717 -81805 -43673 -81761
rect -43617 -81805 -43573 -81761
rect -43517 -81805 -43473 -81761
rect -43417 -81805 -43373 -81761
rect -43317 -81805 -43273 -81761
rect -43217 -81805 -43173 -81761
rect -43117 -81805 -43073 -81761
rect -43017 -81805 -42973 -81761
rect -42917 -81805 -42873 -81761
rect -42817 -81805 -42773 -81761
rect -42717 -81805 -42673 -81761
rect -42617 -81805 -42573 -81761
rect -42517 -81805 -42473 -81761
rect 80737 -81799 80781 -81755
rect 80837 -81799 80881 -81755
rect 80937 -81799 80981 -81755
rect 81037 -81799 81081 -81755
rect 81137 -81799 81181 -81755
rect 81237 -81799 81281 -81755
rect 81337 -81799 81381 -81755
rect 81437 -81799 81481 -81755
rect 81537 -81799 81581 -81755
rect 81637 -81799 81681 -81755
rect 81737 -81799 81781 -81755
rect 81837 -81799 81881 -81755
rect 81937 -81799 81981 -81755
rect 82037 -81799 82081 -81755
rect 82137 -81799 82181 -81755
rect 82237 -81799 82281 -81755
rect 82737 -81799 82781 -81755
rect 82837 -81799 82881 -81755
rect 82937 -81799 82981 -81755
rect 83037 -81799 83081 -81755
rect 83137 -81799 83181 -81755
rect 83237 -81799 83281 -81755
rect 83337 -81799 83381 -81755
rect 83437 -81799 83481 -81755
rect 83537 -81799 83581 -81755
rect 83637 -81799 83681 -81755
rect 83737 -81799 83781 -81755
rect 83837 -81799 83881 -81755
rect 83937 -81799 83981 -81755
rect 84037 -81799 84081 -81755
rect 84137 -81799 84181 -81755
rect 84237 -81799 84281 -81755
rect 84737 -81799 84781 -81755
rect 84837 -81799 84881 -81755
rect 84937 -81799 84981 -81755
rect 85037 -81799 85081 -81755
rect 85137 -81799 85181 -81755
rect 85237 -81799 85281 -81755
rect 85337 -81799 85381 -81755
rect 85437 -81799 85481 -81755
rect 85537 -81799 85581 -81755
rect 85637 -81799 85681 -81755
rect 85737 -81799 85781 -81755
rect 85837 -81799 85881 -81755
rect 85937 -81799 85981 -81755
rect 86037 -81799 86081 -81755
rect 86137 -81799 86181 -81755
rect 86237 -81799 86281 -81755
rect 86737 -81799 86781 -81755
rect 86837 -81799 86881 -81755
rect 86937 -81799 86981 -81755
rect 87037 -81799 87081 -81755
rect 87137 -81799 87181 -81755
rect 87237 -81799 87281 -81755
rect 87337 -81799 87381 -81755
rect 87437 -81799 87481 -81755
rect 87537 -81799 87581 -81755
rect 87637 -81799 87681 -81755
rect 87737 -81799 87781 -81755
rect 87837 -81799 87881 -81755
rect 87937 -81799 87981 -81755
rect 88037 -81799 88081 -81755
rect 88137 -81799 88181 -81755
rect 88237 -81799 88281 -81755
rect -82968 -81903 -82924 -81859
rect -82868 -81903 -82824 -81859
rect -82768 -81903 -82724 -81859
rect -82668 -81903 -82624 -81859
rect -82568 -81903 -82524 -81859
rect -82468 -81903 -82424 -81859
rect -82368 -81903 -82324 -81859
rect -82268 -81903 -82224 -81859
rect -82168 -81903 -82124 -81859
rect -82068 -81903 -82024 -81859
rect -81968 -81903 -81924 -81859
rect -81868 -81903 -81824 -81859
rect -81768 -81903 -81724 -81859
rect -81668 -81903 -81624 -81859
rect -81568 -81903 -81524 -81859
rect -81468 -81903 -81424 -81859
rect -80968 -81903 -80924 -81859
rect -80868 -81903 -80824 -81859
rect -80768 -81903 -80724 -81859
rect -80668 -81903 -80624 -81859
rect -80568 -81903 -80524 -81859
rect -80468 -81903 -80424 -81859
rect -80368 -81903 -80324 -81859
rect -80268 -81903 -80224 -81859
rect -80168 -81903 -80124 -81859
rect -80068 -81903 -80024 -81859
rect -79968 -81903 -79924 -81859
rect -79868 -81903 -79824 -81859
rect -79768 -81903 -79724 -81859
rect -79668 -81903 -79624 -81859
rect -79568 -81903 -79524 -81859
rect -79468 -81903 -79424 -81859
rect -78968 -81903 -78924 -81859
rect -78868 -81903 -78824 -81859
rect -78768 -81903 -78724 -81859
rect -78668 -81903 -78624 -81859
rect -78568 -81903 -78524 -81859
rect -78468 -81903 -78424 -81859
rect -78368 -81903 -78324 -81859
rect -78268 -81903 -78224 -81859
rect -78168 -81903 -78124 -81859
rect -78068 -81903 -78024 -81859
rect -77968 -81903 -77924 -81859
rect -77868 -81903 -77824 -81859
rect -77768 -81903 -77724 -81859
rect -77668 -81903 -77624 -81859
rect -77568 -81903 -77524 -81859
rect -77468 -81903 -77424 -81859
rect -76968 -81903 -76924 -81859
rect -76868 -81903 -76824 -81859
rect -76768 -81903 -76724 -81859
rect -76668 -81903 -76624 -81859
rect -76568 -81903 -76524 -81859
rect -76468 -81903 -76424 -81859
rect -76368 -81903 -76324 -81859
rect -76268 -81903 -76224 -81859
rect -76168 -81903 -76124 -81859
rect -76068 -81903 -76024 -81859
rect -75968 -81903 -75924 -81859
rect -75868 -81903 -75824 -81859
rect -75768 -81903 -75724 -81859
rect -75668 -81903 -75624 -81859
rect -75568 -81903 -75524 -81859
rect -75468 -81903 -75424 -81859
rect -50017 -81905 -49973 -81861
rect -49917 -81905 -49873 -81861
rect -49817 -81905 -49773 -81861
rect -49717 -81905 -49673 -81861
rect -49617 -81905 -49573 -81861
rect -49517 -81905 -49473 -81861
rect -49417 -81905 -49373 -81861
rect -49317 -81905 -49273 -81861
rect -49217 -81905 -49173 -81861
rect -49117 -81905 -49073 -81861
rect -49017 -81905 -48973 -81861
rect -48917 -81905 -48873 -81861
rect -48817 -81905 -48773 -81861
rect -48717 -81905 -48673 -81861
rect -48617 -81905 -48573 -81861
rect -48517 -81905 -48473 -81861
rect -48017 -81905 -47973 -81861
rect -47917 -81905 -47873 -81861
rect -47817 -81905 -47773 -81861
rect -47717 -81905 -47673 -81861
rect -47617 -81905 -47573 -81861
rect -47517 -81905 -47473 -81861
rect -47417 -81905 -47373 -81861
rect -47317 -81905 -47273 -81861
rect -47217 -81905 -47173 -81861
rect -47117 -81905 -47073 -81861
rect -47017 -81905 -46973 -81861
rect -46917 -81905 -46873 -81861
rect -46817 -81905 -46773 -81861
rect -46717 -81905 -46673 -81861
rect -46617 -81905 -46573 -81861
rect -46517 -81905 -46473 -81861
rect -46017 -81905 -45973 -81861
rect -45917 -81905 -45873 -81861
rect -45817 -81905 -45773 -81861
rect -45717 -81905 -45673 -81861
rect -45617 -81905 -45573 -81861
rect -45517 -81905 -45473 -81861
rect -45417 -81905 -45373 -81861
rect -45317 -81905 -45273 -81861
rect -45217 -81905 -45173 -81861
rect -45117 -81905 -45073 -81861
rect -45017 -81905 -44973 -81861
rect -44917 -81905 -44873 -81861
rect -44817 -81905 -44773 -81861
rect -44717 -81905 -44673 -81861
rect -44617 -81905 -44573 -81861
rect -44517 -81905 -44473 -81861
rect -44017 -81905 -43973 -81861
rect -43917 -81905 -43873 -81861
rect -43817 -81905 -43773 -81861
rect -43717 -81905 -43673 -81861
rect -43617 -81905 -43573 -81861
rect -43517 -81905 -43473 -81861
rect -43417 -81905 -43373 -81861
rect -43317 -81905 -43273 -81861
rect -43217 -81905 -43173 -81861
rect -43117 -81905 -43073 -81861
rect -43017 -81905 -42973 -81861
rect -42917 -81905 -42873 -81861
rect -42817 -81905 -42773 -81861
rect -42717 -81905 -42673 -81861
rect -42617 -81905 -42573 -81861
rect -42517 -81905 -42473 -81861
rect 80737 -81899 80781 -81855
rect 80837 -81899 80881 -81855
rect 80937 -81899 80981 -81855
rect 81037 -81899 81081 -81855
rect 81137 -81899 81181 -81855
rect 81237 -81899 81281 -81855
rect 81337 -81899 81381 -81855
rect 81437 -81899 81481 -81855
rect 81537 -81899 81581 -81855
rect 81637 -81899 81681 -81855
rect 81737 -81899 81781 -81855
rect 81837 -81899 81881 -81855
rect 81937 -81899 81981 -81855
rect 82037 -81899 82081 -81855
rect 82137 -81899 82181 -81855
rect 82237 -81899 82281 -81855
rect 82737 -81899 82781 -81855
rect 82837 -81899 82881 -81855
rect 82937 -81899 82981 -81855
rect 83037 -81899 83081 -81855
rect 83137 -81899 83181 -81855
rect 83237 -81899 83281 -81855
rect 83337 -81899 83381 -81855
rect 83437 -81899 83481 -81855
rect 83537 -81899 83581 -81855
rect 83637 -81899 83681 -81855
rect 83737 -81899 83781 -81855
rect 83837 -81899 83881 -81855
rect 83937 -81899 83981 -81855
rect 84037 -81899 84081 -81855
rect 84137 -81899 84181 -81855
rect 84237 -81899 84281 -81855
rect 84737 -81899 84781 -81855
rect 84837 -81899 84881 -81855
rect 84937 -81899 84981 -81855
rect 85037 -81899 85081 -81855
rect 85137 -81899 85181 -81855
rect 85237 -81899 85281 -81855
rect 85337 -81899 85381 -81855
rect 85437 -81899 85481 -81855
rect 85537 -81899 85581 -81855
rect 85637 -81899 85681 -81855
rect 85737 -81899 85781 -81855
rect 85837 -81899 85881 -81855
rect 85937 -81899 85981 -81855
rect 86037 -81899 86081 -81855
rect 86137 -81899 86181 -81855
rect 86237 -81899 86281 -81855
rect 86737 -81899 86781 -81855
rect 86837 -81899 86881 -81855
rect 86937 -81899 86981 -81855
rect 87037 -81899 87081 -81855
rect 87137 -81899 87181 -81855
rect 87237 -81899 87281 -81855
rect 87337 -81899 87381 -81855
rect 87437 -81899 87481 -81855
rect 87537 -81899 87581 -81855
rect 87637 -81899 87681 -81855
rect 87737 -81899 87781 -81855
rect 87837 -81899 87881 -81855
rect 87937 -81899 87981 -81855
rect 88037 -81899 88081 -81855
rect 88137 -81899 88181 -81855
rect 88237 -81899 88281 -81855
rect -82968 -82003 -82924 -81959
rect -82868 -82003 -82824 -81959
rect -82768 -82003 -82724 -81959
rect -82668 -82003 -82624 -81959
rect -82568 -82003 -82524 -81959
rect -82468 -82003 -82424 -81959
rect -82368 -82003 -82324 -81959
rect -82268 -82003 -82224 -81959
rect -82168 -82003 -82124 -81959
rect -82068 -82003 -82024 -81959
rect -81968 -82003 -81924 -81959
rect -81868 -82003 -81824 -81959
rect -81768 -82003 -81724 -81959
rect -81668 -82003 -81624 -81959
rect -81568 -82003 -81524 -81959
rect -81468 -82003 -81424 -81959
rect -80968 -82003 -80924 -81959
rect -80868 -82003 -80824 -81959
rect -80768 -82003 -80724 -81959
rect -80668 -82003 -80624 -81959
rect -80568 -82003 -80524 -81959
rect -80468 -82003 -80424 -81959
rect -80368 -82003 -80324 -81959
rect -80268 -82003 -80224 -81959
rect -80168 -82003 -80124 -81959
rect -80068 -82003 -80024 -81959
rect -79968 -82003 -79924 -81959
rect -79868 -82003 -79824 -81959
rect -79768 -82003 -79724 -81959
rect -79668 -82003 -79624 -81959
rect -79568 -82003 -79524 -81959
rect -79468 -82003 -79424 -81959
rect -78968 -82003 -78924 -81959
rect -78868 -82003 -78824 -81959
rect -78768 -82003 -78724 -81959
rect -78668 -82003 -78624 -81959
rect -78568 -82003 -78524 -81959
rect -78468 -82003 -78424 -81959
rect -78368 -82003 -78324 -81959
rect -78268 -82003 -78224 -81959
rect -78168 -82003 -78124 -81959
rect -78068 -82003 -78024 -81959
rect -77968 -82003 -77924 -81959
rect -77868 -82003 -77824 -81959
rect -77768 -82003 -77724 -81959
rect -77668 -82003 -77624 -81959
rect -77568 -82003 -77524 -81959
rect -77468 -82003 -77424 -81959
rect -76968 -82003 -76924 -81959
rect -76868 -82003 -76824 -81959
rect -76768 -82003 -76724 -81959
rect -76668 -82003 -76624 -81959
rect -76568 -82003 -76524 -81959
rect -76468 -82003 -76424 -81959
rect -76368 -82003 -76324 -81959
rect -76268 -82003 -76224 -81959
rect -76168 -82003 -76124 -81959
rect -76068 -82003 -76024 -81959
rect -75968 -82003 -75924 -81959
rect -75868 -82003 -75824 -81959
rect -75768 -82003 -75724 -81959
rect -75668 -82003 -75624 -81959
rect -75568 -82003 -75524 -81959
rect -75468 -82003 -75424 -81959
rect -50017 -82005 -49973 -81961
rect -49917 -82005 -49873 -81961
rect -49817 -82005 -49773 -81961
rect -49717 -82005 -49673 -81961
rect -49617 -82005 -49573 -81961
rect -49517 -82005 -49473 -81961
rect -49417 -82005 -49373 -81961
rect -49317 -82005 -49273 -81961
rect -49217 -82005 -49173 -81961
rect -49117 -82005 -49073 -81961
rect -49017 -82005 -48973 -81961
rect -48917 -82005 -48873 -81961
rect -48817 -82005 -48773 -81961
rect -48717 -82005 -48673 -81961
rect -48617 -82005 -48573 -81961
rect -48517 -82005 -48473 -81961
rect -48017 -82005 -47973 -81961
rect -47917 -82005 -47873 -81961
rect -47817 -82005 -47773 -81961
rect -47717 -82005 -47673 -81961
rect -47617 -82005 -47573 -81961
rect -47517 -82005 -47473 -81961
rect -47417 -82005 -47373 -81961
rect -47317 -82005 -47273 -81961
rect -47217 -82005 -47173 -81961
rect -47117 -82005 -47073 -81961
rect -47017 -82005 -46973 -81961
rect -46917 -82005 -46873 -81961
rect -46817 -82005 -46773 -81961
rect -46717 -82005 -46673 -81961
rect -46617 -82005 -46573 -81961
rect -46517 -82005 -46473 -81961
rect -46017 -82005 -45973 -81961
rect -45917 -82005 -45873 -81961
rect -45817 -82005 -45773 -81961
rect -45717 -82005 -45673 -81961
rect -45617 -82005 -45573 -81961
rect -45517 -82005 -45473 -81961
rect -45417 -82005 -45373 -81961
rect -45317 -82005 -45273 -81961
rect -45217 -82005 -45173 -81961
rect -45117 -82005 -45073 -81961
rect -45017 -82005 -44973 -81961
rect -44917 -82005 -44873 -81961
rect -44817 -82005 -44773 -81961
rect -44717 -82005 -44673 -81961
rect -44617 -82005 -44573 -81961
rect -44517 -82005 -44473 -81961
rect -44017 -82005 -43973 -81961
rect -43917 -82005 -43873 -81961
rect -43817 -82005 -43773 -81961
rect -43717 -82005 -43673 -81961
rect -43617 -82005 -43573 -81961
rect -43517 -82005 -43473 -81961
rect -43417 -82005 -43373 -81961
rect -43317 -82005 -43273 -81961
rect -43217 -82005 -43173 -81961
rect -43117 -82005 -43073 -81961
rect -43017 -82005 -42973 -81961
rect -42917 -82005 -42873 -81961
rect -42817 -82005 -42773 -81961
rect -42717 -82005 -42673 -81961
rect -42617 -82005 -42573 -81961
rect -42517 -82005 -42473 -81961
rect 80737 -81999 80781 -81955
rect 80837 -81999 80881 -81955
rect 80937 -81999 80981 -81955
rect 81037 -81999 81081 -81955
rect 81137 -81999 81181 -81955
rect 81237 -81999 81281 -81955
rect 81337 -81999 81381 -81955
rect 81437 -81999 81481 -81955
rect 81537 -81999 81581 -81955
rect 81637 -81999 81681 -81955
rect 81737 -81999 81781 -81955
rect 81837 -81999 81881 -81955
rect 81937 -81999 81981 -81955
rect 82037 -81999 82081 -81955
rect 82137 -81999 82181 -81955
rect 82237 -81999 82281 -81955
rect 82737 -81999 82781 -81955
rect 82837 -81999 82881 -81955
rect 82937 -81999 82981 -81955
rect 83037 -81999 83081 -81955
rect 83137 -81999 83181 -81955
rect 83237 -81999 83281 -81955
rect 83337 -81999 83381 -81955
rect 83437 -81999 83481 -81955
rect 83537 -81999 83581 -81955
rect 83637 -81999 83681 -81955
rect 83737 -81999 83781 -81955
rect 83837 -81999 83881 -81955
rect 83937 -81999 83981 -81955
rect 84037 -81999 84081 -81955
rect 84137 -81999 84181 -81955
rect 84237 -81999 84281 -81955
rect 84737 -81999 84781 -81955
rect 84837 -81999 84881 -81955
rect 84937 -81999 84981 -81955
rect 85037 -81999 85081 -81955
rect 85137 -81999 85181 -81955
rect 85237 -81999 85281 -81955
rect 85337 -81999 85381 -81955
rect 85437 -81999 85481 -81955
rect 85537 -81999 85581 -81955
rect 85637 -81999 85681 -81955
rect 85737 -81999 85781 -81955
rect 85837 -81999 85881 -81955
rect 85937 -81999 85981 -81955
rect 86037 -81999 86081 -81955
rect 86137 -81999 86181 -81955
rect 86237 -81999 86281 -81955
rect 86737 -81999 86781 -81955
rect 86837 -81999 86881 -81955
rect 86937 -81999 86981 -81955
rect 87037 -81999 87081 -81955
rect 87137 -81999 87181 -81955
rect 87237 -81999 87281 -81955
rect 87337 -81999 87381 -81955
rect 87437 -81999 87481 -81955
rect 87537 -81999 87581 -81955
rect 87637 -81999 87681 -81955
rect 87737 -81999 87781 -81955
rect 87837 -81999 87881 -81955
rect 87937 -81999 87981 -81955
rect 88037 -81999 88081 -81955
rect 88137 -81999 88181 -81955
rect 88237 -81999 88281 -81955
rect -50075 -106237 -50031 -106193
rect -49975 -106237 -49931 -106193
rect -49875 -106237 -49831 -106193
rect -49775 -106237 -49731 -106193
rect -49675 -106237 -49631 -106193
rect -49575 -106237 -49531 -106193
rect -49475 -106237 -49431 -106193
rect -49375 -106237 -49331 -106193
rect -49275 -106237 -49231 -106193
rect -49175 -106237 -49131 -106193
rect -49075 -106237 -49031 -106193
rect -48975 -106237 -48931 -106193
rect -48875 -106237 -48831 -106193
rect -48775 -106237 -48731 -106193
rect -48675 -106237 -48631 -106193
rect -48575 -106237 -48531 -106193
rect -48075 -106237 -48031 -106193
rect -47975 -106237 -47931 -106193
rect -47875 -106237 -47831 -106193
rect -47775 -106237 -47731 -106193
rect -47675 -106237 -47631 -106193
rect -47575 -106237 -47531 -106193
rect -47475 -106237 -47431 -106193
rect -47375 -106237 -47331 -106193
rect -47275 -106237 -47231 -106193
rect -47175 -106237 -47131 -106193
rect -47075 -106237 -47031 -106193
rect -46975 -106237 -46931 -106193
rect -46875 -106237 -46831 -106193
rect -46775 -106237 -46731 -106193
rect -46675 -106237 -46631 -106193
rect -46575 -106237 -46531 -106193
rect -46075 -106237 -46031 -106193
rect -45975 -106237 -45931 -106193
rect -45875 -106237 -45831 -106193
rect -45775 -106237 -45731 -106193
rect -45675 -106237 -45631 -106193
rect -45575 -106237 -45531 -106193
rect -45475 -106237 -45431 -106193
rect -45375 -106237 -45331 -106193
rect -45275 -106237 -45231 -106193
rect -45175 -106237 -45131 -106193
rect -45075 -106237 -45031 -106193
rect -44975 -106237 -44931 -106193
rect -44875 -106237 -44831 -106193
rect -44775 -106237 -44731 -106193
rect -44675 -106237 -44631 -106193
rect -44575 -106237 -44531 -106193
rect -44075 -106237 -44031 -106193
rect -43975 -106237 -43931 -106193
rect -43875 -106237 -43831 -106193
rect -43775 -106237 -43731 -106193
rect -43675 -106237 -43631 -106193
rect -43575 -106237 -43531 -106193
rect -43475 -106237 -43431 -106193
rect -43375 -106237 -43331 -106193
rect -43275 -106237 -43231 -106193
rect -43175 -106237 -43131 -106193
rect -43075 -106237 -43031 -106193
rect -42975 -106237 -42931 -106193
rect -42875 -106237 -42831 -106193
rect -42775 -106237 -42731 -106193
rect -42675 -106237 -42631 -106193
rect -42575 -106237 -42531 -106193
rect -50075 -106337 -50031 -106293
rect -49975 -106337 -49931 -106293
rect -49875 -106337 -49831 -106293
rect -49775 -106337 -49731 -106293
rect -49675 -106337 -49631 -106293
rect -49575 -106337 -49531 -106293
rect -49475 -106337 -49431 -106293
rect -49375 -106337 -49331 -106293
rect -49275 -106337 -49231 -106293
rect -49175 -106337 -49131 -106293
rect -49075 -106337 -49031 -106293
rect -48975 -106337 -48931 -106293
rect -48875 -106337 -48831 -106293
rect -48775 -106337 -48731 -106293
rect -48675 -106337 -48631 -106293
rect -48575 -106337 -48531 -106293
rect -48075 -106337 -48031 -106293
rect -47975 -106337 -47931 -106293
rect -47875 -106337 -47831 -106293
rect -47775 -106337 -47731 -106293
rect -47675 -106337 -47631 -106293
rect -47575 -106337 -47531 -106293
rect -47475 -106337 -47431 -106293
rect -47375 -106337 -47331 -106293
rect -47275 -106337 -47231 -106293
rect -47175 -106337 -47131 -106293
rect -47075 -106337 -47031 -106293
rect -46975 -106337 -46931 -106293
rect -46875 -106337 -46831 -106293
rect -46775 -106337 -46731 -106293
rect -46675 -106337 -46631 -106293
rect -46575 -106337 -46531 -106293
rect -46075 -106337 -46031 -106293
rect -45975 -106337 -45931 -106293
rect -45875 -106337 -45831 -106293
rect -45775 -106337 -45731 -106293
rect -45675 -106337 -45631 -106293
rect -45575 -106337 -45531 -106293
rect -45475 -106337 -45431 -106293
rect -45375 -106337 -45331 -106293
rect -45275 -106337 -45231 -106293
rect -45175 -106337 -45131 -106293
rect -45075 -106337 -45031 -106293
rect -44975 -106337 -44931 -106293
rect -44875 -106337 -44831 -106293
rect -44775 -106337 -44731 -106293
rect -44675 -106337 -44631 -106293
rect -44575 -106337 -44531 -106293
rect -44075 -106337 -44031 -106293
rect -43975 -106337 -43931 -106293
rect -43875 -106337 -43831 -106293
rect -43775 -106337 -43731 -106293
rect -43675 -106337 -43631 -106293
rect -43575 -106337 -43531 -106293
rect -43475 -106337 -43431 -106293
rect -43375 -106337 -43331 -106293
rect -43275 -106337 -43231 -106293
rect -43175 -106337 -43131 -106293
rect -43075 -106337 -43031 -106293
rect -42975 -106337 -42931 -106293
rect -42875 -106337 -42831 -106293
rect -42775 -106337 -42731 -106293
rect -42675 -106337 -42631 -106293
rect -42575 -106337 -42531 -106293
rect -50075 -106437 -50031 -106393
rect -49975 -106437 -49931 -106393
rect -49875 -106437 -49831 -106393
rect -49775 -106437 -49731 -106393
rect -49675 -106437 -49631 -106393
rect -49575 -106437 -49531 -106393
rect -49475 -106437 -49431 -106393
rect -49375 -106437 -49331 -106393
rect -49275 -106437 -49231 -106393
rect -49175 -106437 -49131 -106393
rect -49075 -106437 -49031 -106393
rect -48975 -106437 -48931 -106393
rect -48875 -106437 -48831 -106393
rect -48775 -106437 -48731 -106393
rect -48675 -106437 -48631 -106393
rect -48575 -106437 -48531 -106393
rect -48075 -106437 -48031 -106393
rect -47975 -106437 -47931 -106393
rect -47875 -106437 -47831 -106393
rect -47775 -106437 -47731 -106393
rect -47675 -106437 -47631 -106393
rect -47575 -106437 -47531 -106393
rect -47475 -106437 -47431 -106393
rect -47375 -106437 -47331 -106393
rect -47275 -106437 -47231 -106393
rect -47175 -106437 -47131 -106393
rect -47075 -106437 -47031 -106393
rect -46975 -106437 -46931 -106393
rect -46875 -106437 -46831 -106393
rect -46775 -106437 -46731 -106393
rect -46675 -106437 -46631 -106393
rect -46575 -106437 -46531 -106393
rect -46075 -106437 -46031 -106393
rect -45975 -106437 -45931 -106393
rect -45875 -106437 -45831 -106393
rect -45775 -106437 -45731 -106393
rect -45675 -106437 -45631 -106393
rect -45575 -106437 -45531 -106393
rect -45475 -106437 -45431 -106393
rect -45375 -106437 -45331 -106393
rect -45275 -106437 -45231 -106393
rect -45175 -106437 -45131 -106393
rect -45075 -106437 -45031 -106393
rect -44975 -106437 -44931 -106393
rect -44875 -106437 -44831 -106393
rect -44775 -106437 -44731 -106393
rect -44675 -106437 -44631 -106393
rect -44575 -106437 -44531 -106393
rect -44075 -106437 -44031 -106393
rect -43975 -106437 -43931 -106393
rect -43875 -106437 -43831 -106393
rect -43775 -106437 -43731 -106393
rect -43675 -106437 -43631 -106393
rect -43575 -106437 -43531 -106393
rect -43475 -106437 -43431 -106393
rect -43375 -106437 -43331 -106393
rect -43275 -106437 -43231 -106393
rect -43175 -106437 -43131 -106393
rect -43075 -106437 -43031 -106393
rect -42975 -106437 -42931 -106393
rect -42875 -106437 -42831 -106393
rect -42775 -106437 -42731 -106393
rect -42675 -106437 -42631 -106393
rect -42575 -106437 -42531 -106393
rect -50075 -106537 -50031 -106493
rect -49975 -106537 -49931 -106493
rect -49875 -106537 -49831 -106493
rect -49775 -106537 -49731 -106493
rect -49675 -106537 -49631 -106493
rect -49575 -106537 -49531 -106493
rect -49475 -106537 -49431 -106493
rect -49375 -106537 -49331 -106493
rect -49275 -106537 -49231 -106493
rect -49175 -106537 -49131 -106493
rect -49075 -106537 -49031 -106493
rect -48975 -106537 -48931 -106493
rect -48875 -106537 -48831 -106493
rect -48775 -106537 -48731 -106493
rect -48675 -106537 -48631 -106493
rect -48575 -106537 -48531 -106493
rect -48075 -106537 -48031 -106493
rect -47975 -106537 -47931 -106493
rect -47875 -106537 -47831 -106493
rect -47775 -106537 -47731 -106493
rect -47675 -106537 -47631 -106493
rect -47575 -106537 -47531 -106493
rect -47475 -106537 -47431 -106493
rect -47375 -106537 -47331 -106493
rect -47275 -106537 -47231 -106493
rect -47175 -106537 -47131 -106493
rect -47075 -106537 -47031 -106493
rect -46975 -106537 -46931 -106493
rect -46875 -106537 -46831 -106493
rect -46775 -106537 -46731 -106493
rect -46675 -106537 -46631 -106493
rect -46575 -106537 -46531 -106493
rect -46075 -106537 -46031 -106493
rect -45975 -106537 -45931 -106493
rect -45875 -106537 -45831 -106493
rect -45775 -106537 -45731 -106493
rect -45675 -106537 -45631 -106493
rect -45575 -106537 -45531 -106493
rect -45475 -106537 -45431 -106493
rect -45375 -106537 -45331 -106493
rect -45275 -106537 -45231 -106493
rect -45175 -106537 -45131 -106493
rect -45075 -106537 -45031 -106493
rect -44975 -106537 -44931 -106493
rect -44875 -106537 -44831 -106493
rect -44775 -106537 -44731 -106493
rect -44675 -106537 -44631 -106493
rect -44575 -106537 -44531 -106493
rect -44075 -106537 -44031 -106493
rect -43975 -106537 -43931 -106493
rect -43875 -106537 -43831 -106493
rect -43775 -106537 -43731 -106493
rect -43675 -106537 -43631 -106493
rect -43575 -106537 -43531 -106493
rect -43475 -106537 -43431 -106493
rect -43375 -106537 -43331 -106493
rect -43275 -106537 -43231 -106493
rect -43175 -106537 -43131 -106493
rect -43075 -106537 -43031 -106493
rect -42975 -106537 -42931 -106493
rect -42875 -106537 -42831 -106493
rect -42775 -106537 -42731 -106493
rect -42675 -106537 -42631 -106493
rect -42575 -106537 -42531 -106493
rect -50075 -106637 -50031 -106593
rect -49975 -106637 -49931 -106593
rect -49875 -106637 -49831 -106593
rect -49775 -106637 -49731 -106593
rect -49675 -106637 -49631 -106593
rect -49575 -106637 -49531 -106593
rect -49475 -106637 -49431 -106593
rect -49375 -106637 -49331 -106593
rect -49275 -106637 -49231 -106593
rect -49175 -106637 -49131 -106593
rect -49075 -106637 -49031 -106593
rect -48975 -106637 -48931 -106593
rect -48875 -106637 -48831 -106593
rect -48775 -106637 -48731 -106593
rect -48675 -106637 -48631 -106593
rect -48575 -106637 -48531 -106593
rect -48075 -106637 -48031 -106593
rect -47975 -106637 -47931 -106593
rect -47875 -106637 -47831 -106593
rect -47775 -106637 -47731 -106593
rect -47675 -106637 -47631 -106593
rect -47575 -106637 -47531 -106593
rect -47475 -106637 -47431 -106593
rect -47375 -106637 -47331 -106593
rect -47275 -106637 -47231 -106593
rect -47175 -106637 -47131 -106593
rect -47075 -106637 -47031 -106593
rect -46975 -106637 -46931 -106593
rect -46875 -106637 -46831 -106593
rect -46775 -106637 -46731 -106593
rect -46675 -106637 -46631 -106593
rect -46575 -106637 -46531 -106593
rect -46075 -106637 -46031 -106593
rect -45975 -106637 -45931 -106593
rect -45875 -106637 -45831 -106593
rect -45775 -106637 -45731 -106593
rect -45675 -106637 -45631 -106593
rect -45575 -106637 -45531 -106593
rect -45475 -106637 -45431 -106593
rect -45375 -106637 -45331 -106593
rect -45275 -106637 -45231 -106593
rect -45175 -106637 -45131 -106593
rect -45075 -106637 -45031 -106593
rect -44975 -106637 -44931 -106593
rect -44875 -106637 -44831 -106593
rect -44775 -106637 -44731 -106593
rect -44675 -106637 -44631 -106593
rect -44575 -106637 -44531 -106593
rect -44075 -106637 -44031 -106593
rect -43975 -106637 -43931 -106593
rect -43875 -106637 -43831 -106593
rect -43775 -106637 -43731 -106593
rect -43675 -106637 -43631 -106593
rect -43575 -106637 -43531 -106593
rect -43475 -106637 -43431 -106593
rect -43375 -106637 -43331 -106593
rect -43275 -106637 -43231 -106593
rect -43175 -106637 -43131 -106593
rect -43075 -106637 -43031 -106593
rect -42975 -106637 -42931 -106593
rect -42875 -106637 -42831 -106593
rect -42775 -106637 -42731 -106593
rect -42675 -106637 -42631 -106593
rect -42575 -106637 -42531 -106593
rect -50075 -106737 -50031 -106693
rect -49975 -106737 -49931 -106693
rect -49875 -106737 -49831 -106693
rect -49775 -106737 -49731 -106693
rect -49675 -106737 -49631 -106693
rect -49575 -106737 -49531 -106693
rect -49475 -106737 -49431 -106693
rect -49375 -106737 -49331 -106693
rect -49275 -106737 -49231 -106693
rect -49175 -106737 -49131 -106693
rect -49075 -106737 -49031 -106693
rect -48975 -106737 -48931 -106693
rect -48875 -106737 -48831 -106693
rect -48775 -106737 -48731 -106693
rect -48675 -106737 -48631 -106693
rect -48575 -106737 -48531 -106693
rect -48075 -106737 -48031 -106693
rect -47975 -106737 -47931 -106693
rect -47875 -106737 -47831 -106693
rect -47775 -106737 -47731 -106693
rect -47675 -106737 -47631 -106693
rect -47575 -106737 -47531 -106693
rect -47475 -106737 -47431 -106693
rect -47375 -106737 -47331 -106693
rect -47275 -106737 -47231 -106693
rect -47175 -106737 -47131 -106693
rect -47075 -106737 -47031 -106693
rect -46975 -106737 -46931 -106693
rect -46875 -106737 -46831 -106693
rect -46775 -106737 -46731 -106693
rect -46675 -106737 -46631 -106693
rect -46575 -106737 -46531 -106693
rect -46075 -106737 -46031 -106693
rect -45975 -106737 -45931 -106693
rect -45875 -106737 -45831 -106693
rect -45775 -106737 -45731 -106693
rect -45675 -106737 -45631 -106693
rect -45575 -106737 -45531 -106693
rect -45475 -106737 -45431 -106693
rect -45375 -106737 -45331 -106693
rect -45275 -106737 -45231 -106693
rect -45175 -106737 -45131 -106693
rect -45075 -106737 -45031 -106693
rect -44975 -106737 -44931 -106693
rect -44875 -106737 -44831 -106693
rect -44775 -106737 -44731 -106693
rect -44675 -106737 -44631 -106693
rect -44575 -106737 -44531 -106693
rect -44075 -106737 -44031 -106693
rect -43975 -106737 -43931 -106693
rect -43875 -106737 -43831 -106693
rect -43775 -106737 -43731 -106693
rect -43675 -106737 -43631 -106693
rect -43575 -106737 -43531 -106693
rect -43475 -106737 -43431 -106693
rect -43375 -106737 -43331 -106693
rect -43275 -106737 -43231 -106693
rect -43175 -106737 -43131 -106693
rect -43075 -106737 -43031 -106693
rect -42975 -106737 -42931 -106693
rect -42875 -106737 -42831 -106693
rect -42775 -106737 -42731 -106693
rect -42675 -106737 -42631 -106693
rect -42575 -106737 -42531 -106693
rect -50075 -106837 -50031 -106793
rect -49975 -106837 -49931 -106793
rect -49875 -106837 -49831 -106793
rect -49775 -106837 -49731 -106793
rect -49675 -106837 -49631 -106793
rect -49575 -106837 -49531 -106793
rect -49475 -106837 -49431 -106793
rect -49375 -106837 -49331 -106793
rect -49275 -106837 -49231 -106793
rect -49175 -106837 -49131 -106793
rect -49075 -106837 -49031 -106793
rect -48975 -106837 -48931 -106793
rect -48875 -106837 -48831 -106793
rect -48775 -106837 -48731 -106793
rect -48675 -106837 -48631 -106793
rect -48575 -106837 -48531 -106793
rect -48075 -106837 -48031 -106793
rect -47975 -106837 -47931 -106793
rect -47875 -106837 -47831 -106793
rect -47775 -106837 -47731 -106793
rect -47675 -106837 -47631 -106793
rect -47575 -106837 -47531 -106793
rect -47475 -106837 -47431 -106793
rect -47375 -106837 -47331 -106793
rect -47275 -106837 -47231 -106793
rect -47175 -106837 -47131 -106793
rect -47075 -106837 -47031 -106793
rect -46975 -106837 -46931 -106793
rect -46875 -106837 -46831 -106793
rect -46775 -106837 -46731 -106793
rect -46675 -106837 -46631 -106793
rect -46575 -106837 -46531 -106793
rect -46075 -106837 -46031 -106793
rect -45975 -106837 -45931 -106793
rect -45875 -106837 -45831 -106793
rect -45775 -106837 -45731 -106793
rect -45675 -106837 -45631 -106793
rect -45575 -106837 -45531 -106793
rect -45475 -106837 -45431 -106793
rect -45375 -106837 -45331 -106793
rect -45275 -106837 -45231 -106793
rect -45175 -106837 -45131 -106793
rect -45075 -106837 -45031 -106793
rect -44975 -106837 -44931 -106793
rect -44875 -106837 -44831 -106793
rect -44775 -106837 -44731 -106793
rect -44675 -106837 -44631 -106793
rect -44575 -106837 -44531 -106793
rect -44075 -106837 -44031 -106793
rect -43975 -106837 -43931 -106793
rect -43875 -106837 -43831 -106793
rect -43775 -106837 -43731 -106793
rect -43675 -106837 -43631 -106793
rect -43575 -106837 -43531 -106793
rect -43475 -106837 -43431 -106793
rect -43375 -106837 -43331 -106793
rect -43275 -106837 -43231 -106793
rect -43175 -106837 -43131 -106793
rect -43075 -106837 -43031 -106793
rect -42975 -106837 -42931 -106793
rect -42875 -106837 -42831 -106793
rect -42775 -106837 -42731 -106793
rect -42675 -106837 -42631 -106793
rect -42575 -106837 -42531 -106793
rect -50075 -106937 -50031 -106893
rect -49975 -106937 -49931 -106893
rect -49875 -106937 -49831 -106893
rect -49775 -106937 -49731 -106893
rect -49675 -106937 -49631 -106893
rect -49575 -106937 -49531 -106893
rect -49475 -106937 -49431 -106893
rect -49375 -106937 -49331 -106893
rect -49275 -106937 -49231 -106893
rect -49175 -106937 -49131 -106893
rect -49075 -106937 -49031 -106893
rect -48975 -106937 -48931 -106893
rect -48875 -106937 -48831 -106893
rect -48775 -106937 -48731 -106893
rect -48675 -106937 -48631 -106893
rect -48575 -106937 -48531 -106893
rect -48075 -106937 -48031 -106893
rect -47975 -106937 -47931 -106893
rect -47875 -106937 -47831 -106893
rect -47775 -106937 -47731 -106893
rect -47675 -106937 -47631 -106893
rect -47575 -106937 -47531 -106893
rect -47475 -106937 -47431 -106893
rect -47375 -106937 -47331 -106893
rect -47275 -106937 -47231 -106893
rect -47175 -106937 -47131 -106893
rect -47075 -106937 -47031 -106893
rect -46975 -106937 -46931 -106893
rect -46875 -106937 -46831 -106893
rect -46775 -106937 -46731 -106893
rect -46675 -106937 -46631 -106893
rect -46575 -106937 -46531 -106893
rect -46075 -106937 -46031 -106893
rect -45975 -106937 -45931 -106893
rect -45875 -106937 -45831 -106893
rect -45775 -106937 -45731 -106893
rect -45675 -106937 -45631 -106893
rect -45575 -106937 -45531 -106893
rect -45475 -106937 -45431 -106893
rect -45375 -106937 -45331 -106893
rect -45275 -106937 -45231 -106893
rect -45175 -106937 -45131 -106893
rect -45075 -106937 -45031 -106893
rect -44975 -106937 -44931 -106893
rect -44875 -106937 -44831 -106893
rect -44775 -106937 -44731 -106893
rect -44675 -106937 -44631 -106893
rect -44575 -106937 -44531 -106893
rect -44075 -106937 -44031 -106893
rect -43975 -106937 -43931 -106893
rect -43875 -106937 -43831 -106893
rect -43775 -106937 -43731 -106893
rect -43675 -106937 -43631 -106893
rect -43575 -106937 -43531 -106893
rect -43475 -106937 -43431 -106893
rect -43375 -106937 -43331 -106893
rect -43275 -106937 -43231 -106893
rect -43175 -106937 -43131 -106893
rect -43075 -106937 -43031 -106893
rect -42975 -106937 -42931 -106893
rect -42875 -106937 -42831 -106893
rect -42775 -106937 -42731 -106893
rect -42675 -106937 -42631 -106893
rect -42575 -106937 -42531 -106893
rect -50075 -107037 -50031 -106993
rect -49975 -107037 -49931 -106993
rect -49875 -107037 -49831 -106993
rect -49775 -107037 -49731 -106993
rect -49675 -107037 -49631 -106993
rect -49575 -107037 -49531 -106993
rect -49475 -107037 -49431 -106993
rect -49375 -107037 -49331 -106993
rect -49275 -107037 -49231 -106993
rect -49175 -107037 -49131 -106993
rect -49075 -107037 -49031 -106993
rect -48975 -107037 -48931 -106993
rect -48875 -107037 -48831 -106993
rect -48775 -107037 -48731 -106993
rect -48675 -107037 -48631 -106993
rect -48575 -107037 -48531 -106993
rect -48075 -107037 -48031 -106993
rect -47975 -107037 -47931 -106993
rect -47875 -107037 -47831 -106993
rect -47775 -107037 -47731 -106993
rect -47675 -107037 -47631 -106993
rect -47575 -107037 -47531 -106993
rect -47475 -107037 -47431 -106993
rect -47375 -107037 -47331 -106993
rect -47275 -107037 -47231 -106993
rect -47175 -107037 -47131 -106993
rect -47075 -107037 -47031 -106993
rect -46975 -107037 -46931 -106993
rect -46875 -107037 -46831 -106993
rect -46775 -107037 -46731 -106993
rect -46675 -107037 -46631 -106993
rect -46575 -107037 -46531 -106993
rect -46075 -107037 -46031 -106993
rect -45975 -107037 -45931 -106993
rect -45875 -107037 -45831 -106993
rect -45775 -107037 -45731 -106993
rect -45675 -107037 -45631 -106993
rect -45575 -107037 -45531 -106993
rect -45475 -107037 -45431 -106993
rect -45375 -107037 -45331 -106993
rect -45275 -107037 -45231 -106993
rect -45175 -107037 -45131 -106993
rect -45075 -107037 -45031 -106993
rect -44975 -107037 -44931 -106993
rect -44875 -107037 -44831 -106993
rect -44775 -107037 -44731 -106993
rect -44675 -107037 -44631 -106993
rect -44575 -107037 -44531 -106993
rect -44075 -107037 -44031 -106993
rect -43975 -107037 -43931 -106993
rect -43875 -107037 -43831 -106993
rect -43775 -107037 -43731 -106993
rect -43675 -107037 -43631 -106993
rect -43575 -107037 -43531 -106993
rect -43475 -107037 -43431 -106993
rect -43375 -107037 -43331 -106993
rect -43275 -107037 -43231 -106993
rect -43175 -107037 -43131 -106993
rect -43075 -107037 -43031 -106993
rect -42975 -107037 -42931 -106993
rect -42875 -107037 -42831 -106993
rect -42775 -107037 -42731 -106993
rect -42675 -107037 -42631 -106993
rect -42575 -107037 -42531 -106993
rect -50075 -107137 -50031 -107093
rect -49975 -107137 -49931 -107093
rect -49875 -107137 -49831 -107093
rect -49775 -107137 -49731 -107093
rect -49675 -107137 -49631 -107093
rect -49575 -107137 -49531 -107093
rect -49475 -107137 -49431 -107093
rect -49375 -107137 -49331 -107093
rect -49275 -107137 -49231 -107093
rect -49175 -107137 -49131 -107093
rect -49075 -107137 -49031 -107093
rect -48975 -107137 -48931 -107093
rect -48875 -107137 -48831 -107093
rect -48775 -107137 -48731 -107093
rect -48675 -107137 -48631 -107093
rect -48575 -107137 -48531 -107093
rect -48075 -107137 -48031 -107093
rect -47975 -107137 -47931 -107093
rect -47875 -107137 -47831 -107093
rect -47775 -107137 -47731 -107093
rect -47675 -107137 -47631 -107093
rect -47575 -107137 -47531 -107093
rect -47475 -107137 -47431 -107093
rect -47375 -107137 -47331 -107093
rect -47275 -107137 -47231 -107093
rect -47175 -107137 -47131 -107093
rect -47075 -107137 -47031 -107093
rect -46975 -107137 -46931 -107093
rect -46875 -107137 -46831 -107093
rect -46775 -107137 -46731 -107093
rect -46675 -107137 -46631 -107093
rect -46575 -107137 -46531 -107093
rect -46075 -107137 -46031 -107093
rect -45975 -107137 -45931 -107093
rect -45875 -107137 -45831 -107093
rect -45775 -107137 -45731 -107093
rect -45675 -107137 -45631 -107093
rect -45575 -107137 -45531 -107093
rect -45475 -107137 -45431 -107093
rect -45375 -107137 -45331 -107093
rect -45275 -107137 -45231 -107093
rect -45175 -107137 -45131 -107093
rect -45075 -107137 -45031 -107093
rect -44975 -107137 -44931 -107093
rect -44875 -107137 -44831 -107093
rect -44775 -107137 -44731 -107093
rect -44675 -107137 -44631 -107093
rect -44575 -107137 -44531 -107093
rect -44075 -107137 -44031 -107093
rect -43975 -107137 -43931 -107093
rect -43875 -107137 -43831 -107093
rect -43775 -107137 -43731 -107093
rect -43675 -107137 -43631 -107093
rect -43575 -107137 -43531 -107093
rect -43475 -107137 -43431 -107093
rect -43375 -107137 -43331 -107093
rect -43275 -107137 -43231 -107093
rect -43175 -107137 -43131 -107093
rect -43075 -107137 -43031 -107093
rect -42975 -107137 -42931 -107093
rect -42875 -107137 -42831 -107093
rect -42775 -107137 -42731 -107093
rect -42675 -107137 -42631 -107093
rect -42575 -107137 -42531 -107093
rect -50075 -107237 -50031 -107193
rect -49975 -107237 -49931 -107193
rect -49875 -107237 -49831 -107193
rect -49775 -107237 -49731 -107193
rect -49675 -107237 -49631 -107193
rect -49575 -107237 -49531 -107193
rect -49475 -107237 -49431 -107193
rect -49375 -107237 -49331 -107193
rect -49275 -107237 -49231 -107193
rect -49175 -107237 -49131 -107193
rect -49075 -107237 -49031 -107193
rect -48975 -107237 -48931 -107193
rect -48875 -107237 -48831 -107193
rect -48775 -107237 -48731 -107193
rect -48675 -107237 -48631 -107193
rect -48575 -107237 -48531 -107193
rect -48075 -107237 -48031 -107193
rect -47975 -107237 -47931 -107193
rect -47875 -107237 -47831 -107193
rect -47775 -107237 -47731 -107193
rect -47675 -107237 -47631 -107193
rect -47575 -107237 -47531 -107193
rect -47475 -107237 -47431 -107193
rect -47375 -107237 -47331 -107193
rect -47275 -107237 -47231 -107193
rect -47175 -107237 -47131 -107193
rect -47075 -107237 -47031 -107193
rect -46975 -107237 -46931 -107193
rect -46875 -107237 -46831 -107193
rect -46775 -107237 -46731 -107193
rect -46675 -107237 -46631 -107193
rect -46575 -107237 -46531 -107193
rect -46075 -107237 -46031 -107193
rect -45975 -107237 -45931 -107193
rect -45875 -107237 -45831 -107193
rect -45775 -107237 -45731 -107193
rect -45675 -107237 -45631 -107193
rect -45575 -107237 -45531 -107193
rect -45475 -107237 -45431 -107193
rect -45375 -107237 -45331 -107193
rect -45275 -107237 -45231 -107193
rect -45175 -107237 -45131 -107193
rect -45075 -107237 -45031 -107193
rect -44975 -107237 -44931 -107193
rect -44875 -107237 -44831 -107193
rect -44775 -107237 -44731 -107193
rect -44675 -107237 -44631 -107193
rect -44575 -107237 -44531 -107193
rect -44075 -107237 -44031 -107193
rect -43975 -107237 -43931 -107193
rect -43875 -107237 -43831 -107193
rect -43775 -107237 -43731 -107193
rect -43675 -107237 -43631 -107193
rect -43575 -107237 -43531 -107193
rect -43475 -107237 -43431 -107193
rect -43375 -107237 -43331 -107193
rect -43275 -107237 -43231 -107193
rect -43175 -107237 -43131 -107193
rect -43075 -107237 -43031 -107193
rect -42975 -107237 -42931 -107193
rect -42875 -107237 -42831 -107193
rect -42775 -107237 -42731 -107193
rect -42675 -107237 -42631 -107193
rect -42575 -107237 -42531 -107193
rect -50075 -107337 -50031 -107293
rect -49975 -107337 -49931 -107293
rect -49875 -107337 -49831 -107293
rect -49775 -107337 -49731 -107293
rect -49675 -107337 -49631 -107293
rect -49575 -107337 -49531 -107293
rect -49475 -107337 -49431 -107293
rect -49375 -107337 -49331 -107293
rect -49275 -107337 -49231 -107293
rect -49175 -107337 -49131 -107293
rect -49075 -107337 -49031 -107293
rect -48975 -107337 -48931 -107293
rect -48875 -107337 -48831 -107293
rect -48775 -107337 -48731 -107293
rect -48675 -107337 -48631 -107293
rect -48575 -107337 -48531 -107293
rect -48075 -107337 -48031 -107293
rect -47975 -107337 -47931 -107293
rect -47875 -107337 -47831 -107293
rect -47775 -107337 -47731 -107293
rect -47675 -107337 -47631 -107293
rect -47575 -107337 -47531 -107293
rect -47475 -107337 -47431 -107293
rect -47375 -107337 -47331 -107293
rect -47275 -107337 -47231 -107293
rect -47175 -107337 -47131 -107293
rect -47075 -107337 -47031 -107293
rect -46975 -107337 -46931 -107293
rect -46875 -107337 -46831 -107293
rect -46775 -107337 -46731 -107293
rect -46675 -107337 -46631 -107293
rect -46575 -107337 -46531 -107293
rect -46075 -107337 -46031 -107293
rect -45975 -107337 -45931 -107293
rect -45875 -107337 -45831 -107293
rect -45775 -107337 -45731 -107293
rect -45675 -107337 -45631 -107293
rect -45575 -107337 -45531 -107293
rect -45475 -107337 -45431 -107293
rect -45375 -107337 -45331 -107293
rect -45275 -107337 -45231 -107293
rect -45175 -107337 -45131 -107293
rect -45075 -107337 -45031 -107293
rect -44975 -107337 -44931 -107293
rect -44875 -107337 -44831 -107293
rect -44775 -107337 -44731 -107293
rect -44675 -107337 -44631 -107293
rect -44575 -107337 -44531 -107293
rect -44075 -107337 -44031 -107293
rect -43975 -107337 -43931 -107293
rect -43875 -107337 -43831 -107293
rect -43775 -107337 -43731 -107293
rect -43675 -107337 -43631 -107293
rect -43575 -107337 -43531 -107293
rect -43475 -107337 -43431 -107293
rect -43375 -107337 -43331 -107293
rect -43275 -107337 -43231 -107293
rect -43175 -107337 -43131 -107293
rect -43075 -107337 -43031 -107293
rect -42975 -107337 -42931 -107293
rect -42875 -107337 -42831 -107293
rect -42775 -107337 -42731 -107293
rect -42675 -107337 -42631 -107293
rect -42575 -107337 -42531 -107293
rect -50075 -107437 -50031 -107393
rect -49975 -107437 -49931 -107393
rect -49875 -107437 -49831 -107393
rect -49775 -107437 -49731 -107393
rect -49675 -107437 -49631 -107393
rect -49575 -107437 -49531 -107393
rect -49475 -107437 -49431 -107393
rect -49375 -107437 -49331 -107393
rect -49275 -107437 -49231 -107393
rect -49175 -107437 -49131 -107393
rect -49075 -107437 -49031 -107393
rect -48975 -107437 -48931 -107393
rect -48875 -107437 -48831 -107393
rect -48775 -107437 -48731 -107393
rect -48675 -107437 -48631 -107393
rect -48575 -107437 -48531 -107393
rect -48075 -107437 -48031 -107393
rect -47975 -107437 -47931 -107393
rect -47875 -107437 -47831 -107393
rect -47775 -107437 -47731 -107393
rect -47675 -107437 -47631 -107393
rect -47575 -107437 -47531 -107393
rect -47475 -107437 -47431 -107393
rect -47375 -107437 -47331 -107393
rect -47275 -107437 -47231 -107393
rect -47175 -107437 -47131 -107393
rect -47075 -107437 -47031 -107393
rect -46975 -107437 -46931 -107393
rect -46875 -107437 -46831 -107393
rect -46775 -107437 -46731 -107393
rect -46675 -107437 -46631 -107393
rect -46575 -107437 -46531 -107393
rect -46075 -107437 -46031 -107393
rect -45975 -107437 -45931 -107393
rect -45875 -107437 -45831 -107393
rect -45775 -107437 -45731 -107393
rect -45675 -107437 -45631 -107393
rect -45575 -107437 -45531 -107393
rect -45475 -107437 -45431 -107393
rect -45375 -107437 -45331 -107393
rect -45275 -107437 -45231 -107393
rect -45175 -107437 -45131 -107393
rect -45075 -107437 -45031 -107393
rect -44975 -107437 -44931 -107393
rect -44875 -107437 -44831 -107393
rect -44775 -107437 -44731 -107393
rect -44675 -107437 -44631 -107393
rect -44575 -107437 -44531 -107393
rect -44075 -107437 -44031 -107393
rect -43975 -107437 -43931 -107393
rect -43875 -107437 -43831 -107393
rect -43775 -107437 -43731 -107393
rect -43675 -107437 -43631 -107393
rect -43575 -107437 -43531 -107393
rect -43475 -107437 -43431 -107393
rect -43375 -107437 -43331 -107393
rect -43275 -107437 -43231 -107393
rect -43175 -107437 -43131 -107393
rect -43075 -107437 -43031 -107393
rect -42975 -107437 -42931 -107393
rect -42875 -107437 -42831 -107393
rect -42775 -107437 -42731 -107393
rect -42675 -107437 -42631 -107393
rect -42575 -107437 -42531 -107393
rect -50075 -107537 -50031 -107493
rect -49975 -107537 -49931 -107493
rect -49875 -107537 -49831 -107493
rect -49775 -107537 -49731 -107493
rect -49675 -107537 -49631 -107493
rect -49575 -107537 -49531 -107493
rect -49475 -107537 -49431 -107493
rect -49375 -107537 -49331 -107493
rect -49275 -107537 -49231 -107493
rect -49175 -107537 -49131 -107493
rect -49075 -107537 -49031 -107493
rect -48975 -107537 -48931 -107493
rect -48875 -107537 -48831 -107493
rect -48775 -107537 -48731 -107493
rect -48675 -107537 -48631 -107493
rect -48575 -107537 -48531 -107493
rect -48075 -107537 -48031 -107493
rect -47975 -107537 -47931 -107493
rect -47875 -107537 -47831 -107493
rect -47775 -107537 -47731 -107493
rect -47675 -107537 -47631 -107493
rect -47575 -107537 -47531 -107493
rect -47475 -107537 -47431 -107493
rect -47375 -107537 -47331 -107493
rect -47275 -107537 -47231 -107493
rect -47175 -107537 -47131 -107493
rect -47075 -107537 -47031 -107493
rect -46975 -107537 -46931 -107493
rect -46875 -107537 -46831 -107493
rect -46775 -107537 -46731 -107493
rect -46675 -107537 -46631 -107493
rect -46575 -107537 -46531 -107493
rect -46075 -107537 -46031 -107493
rect -45975 -107537 -45931 -107493
rect -45875 -107537 -45831 -107493
rect -45775 -107537 -45731 -107493
rect -45675 -107537 -45631 -107493
rect -45575 -107537 -45531 -107493
rect -45475 -107537 -45431 -107493
rect -45375 -107537 -45331 -107493
rect -45275 -107537 -45231 -107493
rect -45175 -107537 -45131 -107493
rect -45075 -107537 -45031 -107493
rect -44975 -107537 -44931 -107493
rect -44875 -107537 -44831 -107493
rect -44775 -107537 -44731 -107493
rect -44675 -107537 -44631 -107493
rect -44575 -107537 -44531 -107493
rect -44075 -107537 -44031 -107493
rect -43975 -107537 -43931 -107493
rect -43875 -107537 -43831 -107493
rect -43775 -107537 -43731 -107493
rect -43675 -107537 -43631 -107493
rect -43575 -107537 -43531 -107493
rect -43475 -107537 -43431 -107493
rect -43375 -107537 -43331 -107493
rect -43275 -107537 -43231 -107493
rect -43175 -107537 -43131 -107493
rect -43075 -107537 -43031 -107493
rect -42975 -107537 -42931 -107493
rect -42875 -107537 -42831 -107493
rect -42775 -107537 -42731 -107493
rect -42675 -107537 -42631 -107493
rect -42575 -107537 -42531 -107493
rect -50075 -107637 -50031 -107593
rect -49975 -107637 -49931 -107593
rect -49875 -107637 -49831 -107593
rect -49775 -107637 -49731 -107593
rect -49675 -107637 -49631 -107593
rect -49575 -107637 -49531 -107593
rect -49475 -107637 -49431 -107593
rect -49375 -107637 -49331 -107593
rect -49275 -107637 -49231 -107593
rect -49175 -107637 -49131 -107593
rect -49075 -107637 -49031 -107593
rect -48975 -107637 -48931 -107593
rect -48875 -107637 -48831 -107593
rect -48775 -107637 -48731 -107593
rect -48675 -107637 -48631 -107593
rect -48575 -107637 -48531 -107593
rect -48075 -107637 -48031 -107593
rect -47975 -107637 -47931 -107593
rect -47875 -107637 -47831 -107593
rect -47775 -107637 -47731 -107593
rect -47675 -107637 -47631 -107593
rect -47575 -107637 -47531 -107593
rect -47475 -107637 -47431 -107593
rect -47375 -107637 -47331 -107593
rect -47275 -107637 -47231 -107593
rect -47175 -107637 -47131 -107593
rect -47075 -107637 -47031 -107593
rect -46975 -107637 -46931 -107593
rect -46875 -107637 -46831 -107593
rect -46775 -107637 -46731 -107593
rect -46675 -107637 -46631 -107593
rect -46575 -107637 -46531 -107593
rect -46075 -107637 -46031 -107593
rect -45975 -107637 -45931 -107593
rect -45875 -107637 -45831 -107593
rect -45775 -107637 -45731 -107593
rect -45675 -107637 -45631 -107593
rect -45575 -107637 -45531 -107593
rect -45475 -107637 -45431 -107593
rect -45375 -107637 -45331 -107593
rect -45275 -107637 -45231 -107593
rect -45175 -107637 -45131 -107593
rect -45075 -107637 -45031 -107593
rect -44975 -107637 -44931 -107593
rect -44875 -107637 -44831 -107593
rect -44775 -107637 -44731 -107593
rect -44675 -107637 -44631 -107593
rect -44575 -107637 -44531 -107593
rect -44075 -107637 -44031 -107593
rect -43975 -107637 -43931 -107593
rect -43875 -107637 -43831 -107593
rect -43775 -107637 -43731 -107593
rect -43675 -107637 -43631 -107593
rect -43575 -107637 -43531 -107593
rect -43475 -107637 -43431 -107593
rect -43375 -107637 -43331 -107593
rect -43275 -107637 -43231 -107593
rect -43175 -107637 -43131 -107593
rect -43075 -107637 -43031 -107593
rect -42975 -107637 -42931 -107593
rect -42875 -107637 -42831 -107593
rect -42775 -107637 -42731 -107593
rect -42675 -107637 -42631 -107593
rect -42575 -107637 -42531 -107593
rect -50075 -107737 -50031 -107693
rect -49975 -107737 -49931 -107693
rect -49875 -107737 -49831 -107693
rect -49775 -107737 -49731 -107693
rect -49675 -107737 -49631 -107693
rect -49575 -107737 -49531 -107693
rect -49475 -107737 -49431 -107693
rect -49375 -107737 -49331 -107693
rect -49275 -107737 -49231 -107693
rect -49175 -107737 -49131 -107693
rect -49075 -107737 -49031 -107693
rect -48975 -107737 -48931 -107693
rect -48875 -107737 -48831 -107693
rect -48775 -107737 -48731 -107693
rect -48675 -107737 -48631 -107693
rect -48575 -107737 -48531 -107693
rect -48075 -107737 -48031 -107693
rect -47975 -107737 -47931 -107693
rect -47875 -107737 -47831 -107693
rect -47775 -107737 -47731 -107693
rect -47675 -107737 -47631 -107693
rect -47575 -107737 -47531 -107693
rect -47475 -107737 -47431 -107693
rect -47375 -107737 -47331 -107693
rect -47275 -107737 -47231 -107693
rect -47175 -107737 -47131 -107693
rect -47075 -107737 -47031 -107693
rect -46975 -107737 -46931 -107693
rect -46875 -107737 -46831 -107693
rect -46775 -107737 -46731 -107693
rect -46675 -107737 -46631 -107693
rect -46575 -107737 -46531 -107693
rect -46075 -107737 -46031 -107693
rect -45975 -107737 -45931 -107693
rect -45875 -107737 -45831 -107693
rect -45775 -107737 -45731 -107693
rect -45675 -107737 -45631 -107693
rect -45575 -107737 -45531 -107693
rect -45475 -107737 -45431 -107693
rect -45375 -107737 -45331 -107693
rect -45275 -107737 -45231 -107693
rect -45175 -107737 -45131 -107693
rect -45075 -107737 -45031 -107693
rect -44975 -107737 -44931 -107693
rect -44875 -107737 -44831 -107693
rect -44775 -107737 -44731 -107693
rect -44675 -107737 -44631 -107693
rect -44575 -107737 -44531 -107693
rect -44075 -107737 -44031 -107693
rect -43975 -107737 -43931 -107693
rect -43875 -107737 -43831 -107693
rect -43775 -107737 -43731 -107693
rect -43675 -107737 -43631 -107693
rect -43575 -107737 -43531 -107693
rect -43475 -107737 -43431 -107693
rect -43375 -107737 -43331 -107693
rect -43275 -107737 -43231 -107693
rect -43175 -107737 -43131 -107693
rect -43075 -107737 -43031 -107693
rect -42975 -107737 -42931 -107693
rect -42875 -107737 -42831 -107693
rect -42775 -107737 -42731 -107693
rect -42675 -107737 -42631 -107693
rect -42575 -107737 -42531 -107693
rect -13354 -131295 -13310 -131251
rect -13254 -131295 -13210 -131251
rect -13154 -131295 -13110 -131251
rect -13054 -131295 -13010 -131251
rect -12954 -131295 -12910 -131251
rect -12854 -131295 -12810 -131251
rect -12754 -131295 -12710 -131251
rect -12654 -131295 -12610 -131251
rect -12554 -131295 -12510 -131251
rect -12454 -131295 -12410 -131251
rect -12354 -131295 -12310 -131251
rect -12254 -131295 -12210 -131251
rect -12154 -131295 -12110 -131251
rect -12054 -131295 -12010 -131251
rect -11954 -131295 -11910 -131251
rect -11854 -131295 -11810 -131251
rect -11354 -131295 -11310 -131251
rect -11254 -131295 -11210 -131251
rect -11154 -131295 -11110 -131251
rect -11054 -131295 -11010 -131251
rect -10954 -131295 -10910 -131251
rect -10854 -131295 -10810 -131251
rect -10754 -131295 -10710 -131251
rect -10654 -131295 -10610 -131251
rect -10554 -131295 -10510 -131251
rect -10454 -131295 -10410 -131251
rect -10354 -131295 -10310 -131251
rect -10254 -131295 -10210 -131251
rect -10154 -131295 -10110 -131251
rect -10054 -131295 -10010 -131251
rect -9954 -131295 -9910 -131251
rect -9854 -131295 -9810 -131251
rect -9354 -131295 -9310 -131251
rect -9254 -131295 -9210 -131251
rect -9154 -131295 -9110 -131251
rect -9054 -131295 -9010 -131251
rect -8954 -131295 -8910 -131251
rect -8854 -131295 -8810 -131251
rect -8754 -131295 -8710 -131251
rect -8654 -131295 -8610 -131251
rect -8554 -131295 -8510 -131251
rect -8454 -131295 -8410 -131251
rect -8354 -131295 -8310 -131251
rect -8254 -131295 -8210 -131251
rect -8154 -131295 -8110 -131251
rect -8054 -131295 -8010 -131251
rect -7954 -131295 -7910 -131251
rect -7854 -131295 -7810 -131251
rect -7354 -131295 -7310 -131251
rect -7254 -131295 -7210 -131251
rect -7154 -131295 -7110 -131251
rect -7054 -131295 -7010 -131251
rect -6954 -131295 -6910 -131251
rect -6854 -131295 -6810 -131251
rect -6754 -131295 -6710 -131251
rect -6654 -131295 -6610 -131251
rect -6554 -131295 -6510 -131251
rect -6454 -131295 -6410 -131251
rect -6354 -131295 -6310 -131251
rect -6254 -131295 -6210 -131251
rect -6154 -131295 -6110 -131251
rect -6054 -131295 -6010 -131251
rect -5954 -131295 -5910 -131251
rect -5854 -131295 -5810 -131251
rect -13354 -131395 -13310 -131351
rect -13254 -131395 -13210 -131351
rect -13154 -131395 -13110 -131351
rect -13054 -131395 -13010 -131351
rect -12954 -131395 -12910 -131351
rect -12854 -131395 -12810 -131351
rect -12754 -131395 -12710 -131351
rect -12654 -131395 -12610 -131351
rect -12554 -131395 -12510 -131351
rect -12454 -131395 -12410 -131351
rect -12354 -131395 -12310 -131351
rect -12254 -131395 -12210 -131351
rect -12154 -131395 -12110 -131351
rect -12054 -131395 -12010 -131351
rect -11954 -131395 -11910 -131351
rect -11854 -131395 -11810 -131351
rect -11354 -131395 -11310 -131351
rect -11254 -131395 -11210 -131351
rect -11154 -131395 -11110 -131351
rect -11054 -131395 -11010 -131351
rect -10954 -131395 -10910 -131351
rect -10854 -131395 -10810 -131351
rect -10754 -131395 -10710 -131351
rect -10654 -131395 -10610 -131351
rect -10554 -131395 -10510 -131351
rect -10454 -131395 -10410 -131351
rect -10354 -131395 -10310 -131351
rect -10254 -131395 -10210 -131351
rect -10154 -131395 -10110 -131351
rect -10054 -131395 -10010 -131351
rect -9954 -131395 -9910 -131351
rect -9854 -131395 -9810 -131351
rect -9354 -131395 -9310 -131351
rect -9254 -131395 -9210 -131351
rect -9154 -131395 -9110 -131351
rect -9054 -131395 -9010 -131351
rect -8954 -131395 -8910 -131351
rect -8854 -131395 -8810 -131351
rect -8754 -131395 -8710 -131351
rect -8654 -131395 -8610 -131351
rect -8554 -131395 -8510 -131351
rect -8454 -131395 -8410 -131351
rect -8354 -131395 -8310 -131351
rect -8254 -131395 -8210 -131351
rect -8154 -131395 -8110 -131351
rect -8054 -131395 -8010 -131351
rect -7954 -131395 -7910 -131351
rect -7854 -131395 -7810 -131351
rect -7354 -131395 -7310 -131351
rect -7254 -131395 -7210 -131351
rect -7154 -131395 -7110 -131351
rect -7054 -131395 -7010 -131351
rect -6954 -131395 -6910 -131351
rect -6854 -131395 -6810 -131351
rect -6754 -131395 -6710 -131351
rect -6654 -131395 -6610 -131351
rect -6554 -131395 -6510 -131351
rect -6454 -131395 -6410 -131351
rect -6354 -131395 -6310 -131351
rect -6254 -131395 -6210 -131351
rect -6154 -131395 -6110 -131351
rect -6054 -131395 -6010 -131351
rect -5954 -131395 -5910 -131351
rect -5854 -131395 -5810 -131351
rect 37387 -131429 37431 -131385
rect 37487 -131429 37531 -131385
rect 37587 -131429 37631 -131385
rect 37687 -131429 37731 -131385
rect 37787 -131429 37831 -131385
rect 37887 -131429 37931 -131385
rect 37987 -131429 38031 -131385
rect 38087 -131429 38131 -131385
rect 38187 -131429 38231 -131385
rect 38287 -131429 38331 -131385
rect 38387 -131429 38431 -131385
rect 38487 -131429 38531 -131385
rect 38587 -131429 38631 -131385
rect 38687 -131429 38731 -131385
rect 38787 -131429 38831 -131385
rect 38887 -131429 38931 -131385
rect 39387 -131429 39431 -131385
rect 39487 -131429 39531 -131385
rect 39587 -131429 39631 -131385
rect 39687 -131429 39731 -131385
rect 39787 -131429 39831 -131385
rect 39887 -131429 39931 -131385
rect 39987 -131429 40031 -131385
rect 40087 -131429 40131 -131385
rect 40187 -131429 40231 -131385
rect 40287 -131429 40331 -131385
rect 40387 -131429 40431 -131385
rect 40487 -131429 40531 -131385
rect 40587 -131429 40631 -131385
rect 40687 -131429 40731 -131385
rect 40787 -131429 40831 -131385
rect 40887 -131429 40931 -131385
rect 41387 -131429 41431 -131385
rect 41487 -131429 41531 -131385
rect 41587 -131429 41631 -131385
rect 41687 -131429 41731 -131385
rect 41787 -131429 41831 -131385
rect 41887 -131429 41931 -131385
rect 41987 -131429 42031 -131385
rect 42087 -131429 42131 -131385
rect 42187 -131429 42231 -131385
rect 42287 -131429 42331 -131385
rect 42387 -131429 42431 -131385
rect 42487 -131429 42531 -131385
rect 42587 -131429 42631 -131385
rect 42687 -131429 42731 -131385
rect 42787 -131429 42831 -131385
rect 42887 -131429 42931 -131385
rect 43387 -131429 43431 -131385
rect 43487 -131429 43531 -131385
rect 43587 -131429 43631 -131385
rect 43687 -131429 43731 -131385
rect 43787 -131429 43831 -131385
rect 43887 -131429 43931 -131385
rect 43987 -131429 44031 -131385
rect 44087 -131429 44131 -131385
rect 44187 -131429 44231 -131385
rect 44287 -131429 44331 -131385
rect 44387 -131429 44431 -131385
rect 44487 -131429 44531 -131385
rect 44587 -131429 44631 -131385
rect 44687 -131429 44731 -131385
rect 44787 -131429 44831 -131385
rect 44887 -131429 44931 -131385
rect -13354 -131495 -13310 -131451
rect -13254 -131495 -13210 -131451
rect -13154 -131495 -13110 -131451
rect -13054 -131495 -13010 -131451
rect -12954 -131495 -12910 -131451
rect -12854 -131495 -12810 -131451
rect -12754 -131495 -12710 -131451
rect -12654 -131495 -12610 -131451
rect -12554 -131495 -12510 -131451
rect -12454 -131495 -12410 -131451
rect -12354 -131495 -12310 -131451
rect -12254 -131495 -12210 -131451
rect -12154 -131495 -12110 -131451
rect -12054 -131495 -12010 -131451
rect -11954 -131495 -11910 -131451
rect -11854 -131495 -11810 -131451
rect -11354 -131495 -11310 -131451
rect -11254 -131495 -11210 -131451
rect -11154 -131495 -11110 -131451
rect -11054 -131495 -11010 -131451
rect -10954 -131495 -10910 -131451
rect -10854 -131495 -10810 -131451
rect -10754 -131495 -10710 -131451
rect -10654 -131495 -10610 -131451
rect -10554 -131495 -10510 -131451
rect -10454 -131495 -10410 -131451
rect -10354 -131495 -10310 -131451
rect -10254 -131495 -10210 -131451
rect -10154 -131495 -10110 -131451
rect -10054 -131495 -10010 -131451
rect -9954 -131495 -9910 -131451
rect -9854 -131495 -9810 -131451
rect -9354 -131495 -9310 -131451
rect -9254 -131495 -9210 -131451
rect -9154 -131495 -9110 -131451
rect -9054 -131495 -9010 -131451
rect -8954 -131495 -8910 -131451
rect -8854 -131495 -8810 -131451
rect -8754 -131495 -8710 -131451
rect -8654 -131495 -8610 -131451
rect -8554 -131495 -8510 -131451
rect -8454 -131495 -8410 -131451
rect -8354 -131495 -8310 -131451
rect -8254 -131495 -8210 -131451
rect -8154 -131495 -8110 -131451
rect -8054 -131495 -8010 -131451
rect -7954 -131495 -7910 -131451
rect -7854 -131495 -7810 -131451
rect -7354 -131495 -7310 -131451
rect -7254 -131495 -7210 -131451
rect -7154 -131495 -7110 -131451
rect -7054 -131495 -7010 -131451
rect -6954 -131495 -6910 -131451
rect -6854 -131495 -6810 -131451
rect -6754 -131495 -6710 -131451
rect -6654 -131495 -6610 -131451
rect -6554 -131495 -6510 -131451
rect -6454 -131495 -6410 -131451
rect -6354 -131495 -6310 -131451
rect -6254 -131495 -6210 -131451
rect -6154 -131495 -6110 -131451
rect -6054 -131495 -6010 -131451
rect -5954 -131495 -5910 -131451
rect -5854 -131495 -5810 -131451
rect 37387 -131529 37431 -131485
rect 37487 -131529 37531 -131485
rect 37587 -131529 37631 -131485
rect 37687 -131529 37731 -131485
rect 37787 -131529 37831 -131485
rect 37887 -131529 37931 -131485
rect 37987 -131529 38031 -131485
rect 38087 -131529 38131 -131485
rect 38187 -131529 38231 -131485
rect 38287 -131529 38331 -131485
rect 38387 -131529 38431 -131485
rect 38487 -131529 38531 -131485
rect 38587 -131529 38631 -131485
rect 38687 -131529 38731 -131485
rect 38787 -131529 38831 -131485
rect 38887 -131529 38931 -131485
rect 39387 -131529 39431 -131485
rect 39487 -131529 39531 -131485
rect 39587 -131529 39631 -131485
rect 39687 -131529 39731 -131485
rect 39787 -131529 39831 -131485
rect 39887 -131529 39931 -131485
rect 39987 -131529 40031 -131485
rect 40087 -131529 40131 -131485
rect 40187 -131529 40231 -131485
rect 40287 -131529 40331 -131485
rect 40387 -131529 40431 -131485
rect 40487 -131529 40531 -131485
rect 40587 -131529 40631 -131485
rect 40687 -131529 40731 -131485
rect 40787 -131529 40831 -131485
rect 40887 -131529 40931 -131485
rect 41387 -131529 41431 -131485
rect 41487 -131529 41531 -131485
rect 41587 -131529 41631 -131485
rect 41687 -131529 41731 -131485
rect 41787 -131529 41831 -131485
rect 41887 -131529 41931 -131485
rect 41987 -131529 42031 -131485
rect 42087 -131529 42131 -131485
rect 42187 -131529 42231 -131485
rect 42287 -131529 42331 -131485
rect 42387 -131529 42431 -131485
rect 42487 -131529 42531 -131485
rect 42587 -131529 42631 -131485
rect 42687 -131529 42731 -131485
rect 42787 -131529 42831 -131485
rect 42887 -131529 42931 -131485
rect 43387 -131529 43431 -131485
rect 43487 -131529 43531 -131485
rect 43587 -131529 43631 -131485
rect 43687 -131529 43731 -131485
rect 43787 -131529 43831 -131485
rect 43887 -131529 43931 -131485
rect 43987 -131529 44031 -131485
rect 44087 -131529 44131 -131485
rect 44187 -131529 44231 -131485
rect 44287 -131529 44331 -131485
rect 44387 -131529 44431 -131485
rect 44487 -131529 44531 -131485
rect 44587 -131529 44631 -131485
rect 44687 -131529 44731 -131485
rect 44787 -131529 44831 -131485
rect 44887 -131529 44931 -131485
rect -13354 -131595 -13310 -131551
rect -13254 -131595 -13210 -131551
rect -13154 -131595 -13110 -131551
rect -13054 -131595 -13010 -131551
rect -12954 -131595 -12910 -131551
rect -12854 -131595 -12810 -131551
rect -12754 -131595 -12710 -131551
rect -12654 -131595 -12610 -131551
rect -12554 -131595 -12510 -131551
rect -12454 -131595 -12410 -131551
rect -12354 -131595 -12310 -131551
rect -12254 -131595 -12210 -131551
rect -12154 -131595 -12110 -131551
rect -12054 -131595 -12010 -131551
rect -11954 -131595 -11910 -131551
rect -11854 -131595 -11810 -131551
rect -11354 -131595 -11310 -131551
rect -11254 -131595 -11210 -131551
rect -11154 -131595 -11110 -131551
rect -11054 -131595 -11010 -131551
rect -10954 -131595 -10910 -131551
rect -10854 -131595 -10810 -131551
rect -10754 -131595 -10710 -131551
rect -10654 -131595 -10610 -131551
rect -10554 -131595 -10510 -131551
rect -10454 -131595 -10410 -131551
rect -10354 -131595 -10310 -131551
rect -10254 -131595 -10210 -131551
rect -10154 -131595 -10110 -131551
rect -10054 -131595 -10010 -131551
rect -9954 -131595 -9910 -131551
rect -9854 -131595 -9810 -131551
rect -9354 -131595 -9310 -131551
rect -9254 -131595 -9210 -131551
rect -9154 -131595 -9110 -131551
rect -9054 -131595 -9010 -131551
rect -8954 -131595 -8910 -131551
rect -8854 -131595 -8810 -131551
rect -8754 -131595 -8710 -131551
rect -8654 -131595 -8610 -131551
rect -8554 -131595 -8510 -131551
rect -8454 -131595 -8410 -131551
rect -8354 -131595 -8310 -131551
rect -8254 -131595 -8210 -131551
rect -8154 -131595 -8110 -131551
rect -8054 -131595 -8010 -131551
rect -7954 -131595 -7910 -131551
rect -7854 -131595 -7810 -131551
rect -7354 -131595 -7310 -131551
rect -7254 -131595 -7210 -131551
rect -7154 -131595 -7110 -131551
rect -7054 -131595 -7010 -131551
rect -6954 -131595 -6910 -131551
rect -6854 -131595 -6810 -131551
rect -6754 -131595 -6710 -131551
rect -6654 -131595 -6610 -131551
rect -6554 -131595 -6510 -131551
rect -6454 -131595 -6410 -131551
rect -6354 -131595 -6310 -131551
rect -6254 -131595 -6210 -131551
rect -6154 -131595 -6110 -131551
rect -6054 -131595 -6010 -131551
rect -5954 -131595 -5910 -131551
rect -5854 -131595 -5810 -131551
rect 37387 -131629 37431 -131585
rect 37487 -131629 37531 -131585
rect 37587 -131629 37631 -131585
rect 37687 -131629 37731 -131585
rect 37787 -131629 37831 -131585
rect 37887 -131629 37931 -131585
rect 37987 -131629 38031 -131585
rect 38087 -131629 38131 -131585
rect 38187 -131629 38231 -131585
rect 38287 -131629 38331 -131585
rect 38387 -131629 38431 -131585
rect 38487 -131629 38531 -131585
rect 38587 -131629 38631 -131585
rect 38687 -131629 38731 -131585
rect 38787 -131629 38831 -131585
rect 38887 -131629 38931 -131585
rect 39387 -131629 39431 -131585
rect 39487 -131629 39531 -131585
rect 39587 -131629 39631 -131585
rect 39687 -131629 39731 -131585
rect 39787 -131629 39831 -131585
rect 39887 -131629 39931 -131585
rect 39987 -131629 40031 -131585
rect 40087 -131629 40131 -131585
rect 40187 -131629 40231 -131585
rect 40287 -131629 40331 -131585
rect 40387 -131629 40431 -131585
rect 40487 -131629 40531 -131585
rect 40587 -131629 40631 -131585
rect 40687 -131629 40731 -131585
rect 40787 -131629 40831 -131585
rect 40887 -131629 40931 -131585
rect 41387 -131629 41431 -131585
rect 41487 -131629 41531 -131585
rect 41587 -131629 41631 -131585
rect 41687 -131629 41731 -131585
rect 41787 -131629 41831 -131585
rect 41887 -131629 41931 -131585
rect 41987 -131629 42031 -131585
rect 42087 -131629 42131 -131585
rect 42187 -131629 42231 -131585
rect 42287 -131629 42331 -131585
rect 42387 -131629 42431 -131585
rect 42487 -131629 42531 -131585
rect 42587 -131629 42631 -131585
rect 42687 -131629 42731 -131585
rect 42787 -131629 42831 -131585
rect 42887 -131629 42931 -131585
rect 43387 -131629 43431 -131585
rect 43487 -131629 43531 -131585
rect 43587 -131629 43631 -131585
rect 43687 -131629 43731 -131585
rect 43787 -131629 43831 -131585
rect 43887 -131629 43931 -131585
rect 43987 -131629 44031 -131585
rect 44087 -131629 44131 -131585
rect 44187 -131629 44231 -131585
rect 44287 -131629 44331 -131585
rect 44387 -131629 44431 -131585
rect 44487 -131629 44531 -131585
rect 44587 -131629 44631 -131585
rect 44687 -131629 44731 -131585
rect 44787 -131629 44831 -131585
rect 44887 -131629 44931 -131585
rect -13354 -131695 -13310 -131651
rect -13254 -131695 -13210 -131651
rect -13154 -131695 -13110 -131651
rect -13054 -131695 -13010 -131651
rect -12954 -131695 -12910 -131651
rect -12854 -131695 -12810 -131651
rect -12754 -131695 -12710 -131651
rect -12654 -131695 -12610 -131651
rect -12554 -131695 -12510 -131651
rect -12454 -131695 -12410 -131651
rect -12354 -131695 -12310 -131651
rect -12254 -131695 -12210 -131651
rect -12154 -131695 -12110 -131651
rect -12054 -131695 -12010 -131651
rect -11954 -131695 -11910 -131651
rect -11854 -131695 -11810 -131651
rect -11354 -131695 -11310 -131651
rect -11254 -131695 -11210 -131651
rect -11154 -131695 -11110 -131651
rect -11054 -131695 -11010 -131651
rect -10954 -131695 -10910 -131651
rect -10854 -131695 -10810 -131651
rect -10754 -131695 -10710 -131651
rect -10654 -131695 -10610 -131651
rect -10554 -131695 -10510 -131651
rect -10454 -131695 -10410 -131651
rect -10354 -131695 -10310 -131651
rect -10254 -131695 -10210 -131651
rect -10154 -131695 -10110 -131651
rect -10054 -131695 -10010 -131651
rect -9954 -131695 -9910 -131651
rect -9854 -131695 -9810 -131651
rect -9354 -131695 -9310 -131651
rect -9254 -131695 -9210 -131651
rect -9154 -131695 -9110 -131651
rect -9054 -131695 -9010 -131651
rect -8954 -131695 -8910 -131651
rect -8854 -131695 -8810 -131651
rect -8754 -131695 -8710 -131651
rect -8654 -131695 -8610 -131651
rect -8554 -131695 -8510 -131651
rect -8454 -131695 -8410 -131651
rect -8354 -131695 -8310 -131651
rect -8254 -131695 -8210 -131651
rect -8154 -131695 -8110 -131651
rect -8054 -131695 -8010 -131651
rect -7954 -131695 -7910 -131651
rect -7854 -131695 -7810 -131651
rect -7354 -131695 -7310 -131651
rect -7254 -131695 -7210 -131651
rect -7154 -131695 -7110 -131651
rect -7054 -131695 -7010 -131651
rect -6954 -131695 -6910 -131651
rect -6854 -131695 -6810 -131651
rect -6754 -131695 -6710 -131651
rect -6654 -131695 -6610 -131651
rect -6554 -131695 -6510 -131651
rect -6454 -131695 -6410 -131651
rect -6354 -131695 -6310 -131651
rect -6254 -131695 -6210 -131651
rect -6154 -131695 -6110 -131651
rect -6054 -131695 -6010 -131651
rect -5954 -131695 -5910 -131651
rect -5854 -131695 -5810 -131651
rect 37387 -131729 37431 -131685
rect 37487 -131729 37531 -131685
rect 37587 -131729 37631 -131685
rect 37687 -131729 37731 -131685
rect 37787 -131729 37831 -131685
rect 37887 -131729 37931 -131685
rect 37987 -131729 38031 -131685
rect 38087 -131729 38131 -131685
rect 38187 -131729 38231 -131685
rect 38287 -131729 38331 -131685
rect 38387 -131729 38431 -131685
rect 38487 -131729 38531 -131685
rect 38587 -131729 38631 -131685
rect 38687 -131729 38731 -131685
rect 38787 -131729 38831 -131685
rect 38887 -131729 38931 -131685
rect 39387 -131729 39431 -131685
rect 39487 -131729 39531 -131685
rect 39587 -131729 39631 -131685
rect 39687 -131729 39731 -131685
rect 39787 -131729 39831 -131685
rect 39887 -131729 39931 -131685
rect 39987 -131729 40031 -131685
rect 40087 -131729 40131 -131685
rect 40187 -131729 40231 -131685
rect 40287 -131729 40331 -131685
rect 40387 -131729 40431 -131685
rect 40487 -131729 40531 -131685
rect 40587 -131729 40631 -131685
rect 40687 -131729 40731 -131685
rect 40787 -131729 40831 -131685
rect 40887 -131729 40931 -131685
rect 41387 -131729 41431 -131685
rect 41487 -131729 41531 -131685
rect 41587 -131729 41631 -131685
rect 41687 -131729 41731 -131685
rect 41787 -131729 41831 -131685
rect 41887 -131729 41931 -131685
rect 41987 -131729 42031 -131685
rect 42087 -131729 42131 -131685
rect 42187 -131729 42231 -131685
rect 42287 -131729 42331 -131685
rect 42387 -131729 42431 -131685
rect 42487 -131729 42531 -131685
rect 42587 -131729 42631 -131685
rect 42687 -131729 42731 -131685
rect 42787 -131729 42831 -131685
rect 42887 -131729 42931 -131685
rect 43387 -131729 43431 -131685
rect 43487 -131729 43531 -131685
rect 43587 -131729 43631 -131685
rect 43687 -131729 43731 -131685
rect 43787 -131729 43831 -131685
rect 43887 -131729 43931 -131685
rect 43987 -131729 44031 -131685
rect 44087 -131729 44131 -131685
rect 44187 -131729 44231 -131685
rect 44287 -131729 44331 -131685
rect 44387 -131729 44431 -131685
rect 44487 -131729 44531 -131685
rect 44587 -131729 44631 -131685
rect 44687 -131729 44731 -131685
rect 44787 -131729 44831 -131685
rect 44887 -131729 44931 -131685
rect -13354 -131795 -13310 -131751
rect -13254 -131795 -13210 -131751
rect -13154 -131795 -13110 -131751
rect -13054 -131795 -13010 -131751
rect -12954 -131795 -12910 -131751
rect -12854 -131795 -12810 -131751
rect -12754 -131795 -12710 -131751
rect -12654 -131795 -12610 -131751
rect -12554 -131795 -12510 -131751
rect -12454 -131795 -12410 -131751
rect -12354 -131795 -12310 -131751
rect -12254 -131795 -12210 -131751
rect -12154 -131795 -12110 -131751
rect -12054 -131795 -12010 -131751
rect -11954 -131795 -11910 -131751
rect -11854 -131795 -11810 -131751
rect -11354 -131795 -11310 -131751
rect -11254 -131795 -11210 -131751
rect -11154 -131795 -11110 -131751
rect -11054 -131795 -11010 -131751
rect -10954 -131795 -10910 -131751
rect -10854 -131795 -10810 -131751
rect -10754 -131795 -10710 -131751
rect -10654 -131795 -10610 -131751
rect -10554 -131795 -10510 -131751
rect -10454 -131795 -10410 -131751
rect -10354 -131795 -10310 -131751
rect -10254 -131795 -10210 -131751
rect -10154 -131795 -10110 -131751
rect -10054 -131795 -10010 -131751
rect -9954 -131795 -9910 -131751
rect -9854 -131795 -9810 -131751
rect -9354 -131795 -9310 -131751
rect -9254 -131795 -9210 -131751
rect -9154 -131795 -9110 -131751
rect -9054 -131795 -9010 -131751
rect -8954 -131795 -8910 -131751
rect -8854 -131795 -8810 -131751
rect -8754 -131795 -8710 -131751
rect -8654 -131795 -8610 -131751
rect -8554 -131795 -8510 -131751
rect -8454 -131795 -8410 -131751
rect -8354 -131795 -8310 -131751
rect -8254 -131795 -8210 -131751
rect -8154 -131795 -8110 -131751
rect -8054 -131795 -8010 -131751
rect -7954 -131795 -7910 -131751
rect -7854 -131795 -7810 -131751
rect -7354 -131795 -7310 -131751
rect -7254 -131795 -7210 -131751
rect -7154 -131795 -7110 -131751
rect -7054 -131795 -7010 -131751
rect -6954 -131795 -6910 -131751
rect -6854 -131795 -6810 -131751
rect -6754 -131795 -6710 -131751
rect -6654 -131795 -6610 -131751
rect -6554 -131795 -6510 -131751
rect -6454 -131795 -6410 -131751
rect -6354 -131795 -6310 -131751
rect -6254 -131795 -6210 -131751
rect -6154 -131795 -6110 -131751
rect -6054 -131795 -6010 -131751
rect -5954 -131795 -5910 -131751
rect -5854 -131795 -5810 -131751
rect 37387 -131829 37431 -131785
rect 37487 -131829 37531 -131785
rect 37587 -131829 37631 -131785
rect 37687 -131829 37731 -131785
rect 37787 -131829 37831 -131785
rect 37887 -131829 37931 -131785
rect 37987 -131829 38031 -131785
rect 38087 -131829 38131 -131785
rect 38187 -131829 38231 -131785
rect 38287 -131829 38331 -131785
rect 38387 -131829 38431 -131785
rect 38487 -131829 38531 -131785
rect 38587 -131829 38631 -131785
rect 38687 -131829 38731 -131785
rect 38787 -131829 38831 -131785
rect 38887 -131829 38931 -131785
rect 39387 -131829 39431 -131785
rect 39487 -131829 39531 -131785
rect 39587 -131829 39631 -131785
rect 39687 -131829 39731 -131785
rect 39787 -131829 39831 -131785
rect 39887 -131829 39931 -131785
rect 39987 -131829 40031 -131785
rect 40087 -131829 40131 -131785
rect 40187 -131829 40231 -131785
rect 40287 -131829 40331 -131785
rect 40387 -131829 40431 -131785
rect 40487 -131829 40531 -131785
rect 40587 -131829 40631 -131785
rect 40687 -131829 40731 -131785
rect 40787 -131829 40831 -131785
rect 40887 -131829 40931 -131785
rect 41387 -131829 41431 -131785
rect 41487 -131829 41531 -131785
rect 41587 -131829 41631 -131785
rect 41687 -131829 41731 -131785
rect 41787 -131829 41831 -131785
rect 41887 -131829 41931 -131785
rect 41987 -131829 42031 -131785
rect 42087 -131829 42131 -131785
rect 42187 -131829 42231 -131785
rect 42287 -131829 42331 -131785
rect 42387 -131829 42431 -131785
rect 42487 -131829 42531 -131785
rect 42587 -131829 42631 -131785
rect 42687 -131829 42731 -131785
rect 42787 -131829 42831 -131785
rect 42887 -131829 42931 -131785
rect 43387 -131829 43431 -131785
rect 43487 -131829 43531 -131785
rect 43587 -131829 43631 -131785
rect 43687 -131829 43731 -131785
rect 43787 -131829 43831 -131785
rect 43887 -131829 43931 -131785
rect 43987 -131829 44031 -131785
rect 44087 -131829 44131 -131785
rect 44187 -131829 44231 -131785
rect 44287 -131829 44331 -131785
rect 44387 -131829 44431 -131785
rect 44487 -131829 44531 -131785
rect 44587 -131829 44631 -131785
rect 44687 -131829 44731 -131785
rect 44787 -131829 44831 -131785
rect 44887 -131829 44931 -131785
rect -13354 -131895 -13310 -131851
rect -13254 -131895 -13210 -131851
rect -13154 -131895 -13110 -131851
rect -13054 -131895 -13010 -131851
rect -12954 -131895 -12910 -131851
rect -12854 -131895 -12810 -131851
rect -12754 -131895 -12710 -131851
rect -12654 -131895 -12610 -131851
rect -12554 -131895 -12510 -131851
rect -12454 -131895 -12410 -131851
rect -12354 -131895 -12310 -131851
rect -12254 -131895 -12210 -131851
rect -12154 -131895 -12110 -131851
rect -12054 -131895 -12010 -131851
rect -11954 -131895 -11910 -131851
rect -11854 -131895 -11810 -131851
rect -11354 -131895 -11310 -131851
rect -11254 -131895 -11210 -131851
rect -11154 -131895 -11110 -131851
rect -11054 -131895 -11010 -131851
rect -10954 -131895 -10910 -131851
rect -10854 -131895 -10810 -131851
rect -10754 -131895 -10710 -131851
rect -10654 -131895 -10610 -131851
rect -10554 -131895 -10510 -131851
rect -10454 -131895 -10410 -131851
rect -10354 -131895 -10310 -131851
rect -10254 -131895 -10210 -131851
rect -10154 -131895 -10110 -131851
rect -10054 -131895 -10010 -131851
rect -9954 -131895 -9910 -131851
rect -9854 -131895 -9810 -131851
rect -9354 -131895 -9310 -131851
rect -9254 -131895 -9210 -131851
rect -9154 -131895 -9110 -131851
rect -9054 -131895 -9010 -131851
rect -8954 -131895 -8910 -131851
rect -8854 -131895 -8810 -131851
rect -8754 -131895 -8710 -131851
rect -8654 -131895 -8610 -131851
rect -8554 -131895 -8510 -131851
rect -8454 -131895 -8410 -131851
rect -8354 -131895 -8310 -131851
rect -8254 -131895 -8210 -131851
rect -8154 -131895 -8110 -131851
rect -8054 -131895 -8010 -131851
rect -7954 -131895 -7910 -131851
rect -7854 -131895 -7810 -131851
rect -7354 -131895 -7310 -131851
rect -7254 -131895 -7210 -131851
rect -7154 -131895 -7110 -131851
rect -7054 -131895 -7010 -131851
rect -6954 -131895 -6910 -131851
rect -6854 -131895 -6810 -131851
rect -6754 -131895 -6710 -131851
rect -6654 -131895 -6610 -131851
rect -6554 -131895 -6510 -131851
rect -6454 -131895 -6410 -131851
rect -6354 -131895 -6310 -131851
rect -6254 -131895 -6210 -131851
rect -6154 -131895 -6110 -131851
rect -6054 -131895 -6010 -131851
rect -5954 -131895 -5910 -131851
rect -5854 -131895 -5810 -131851
rect 37387 -131929 37431 -131885
rect 37487 -131929 37531 -131885
rect 37587 -131929 37631 -131885
rect 37687 -131929 37731 -131885
rect 37787 -131929 37831 -131885
rect 37887 -131929 37931 -131885
rect 37987 -131929 38031 -131885
rect 38087 -131929 38131 -131885
rect 38187 -131929 38231 -131885
rect 38287 -131929 38331 -131885
rect 38387 -131929 38431 -131885
rect 38487 -131929 38531 -131885
rect 38587 -131929 38631 -131885
rect 38687 -131929 38731 -131885
rect 38787 -131929 38831 -131885
rect 38887 -131929 38931 -131885
rect 39387 -131929 39431 -131885
rect 39487 -131929 39531 -131885
rect 39587 -131929 39631 -131885
rect 39687 -131929 39731 -131885
rect 39787 -131929 39831 -131885
rect 39887 -131929 39931 -131885
rect 39987 -131929 40031 -131885
rect 40087 -131929 40131 -131885
rect 40187 -131929 40231 -131885
rect 40287 -131929 40331 -131885
rect 40387 -131929 40431 -131885
rect 40487 -131929 40531 -131885
rect 40587 -131929 40631 -131885
rect 40687 -131929 40731 -131885
rect 40787 -131929 40831 -131885
rect 40887 -131929 40931 -131885
rect 41387 -131929 41431 -131885
rect 41487 -131929 41531 -131885
rect 41587 -131929 41631 -131885
rect 41687 -131929 41731 -131885
rect 41787 -131929 41831 -131885
rect 41887 -131929 41931 -131885
rect 41987 -131929 42031 -131885
rect 42087 -131929 42131 -131885
rect 42187 -131929 42231 -131885
rect 42287 -131929 42331 -131885
rect 42387 -131929 42431 -131885
rect 42487 -131929 42531 -131885
rect 42587 -131929 42631 -131885
rect 42687 -131929 42731 -131885
rect 42787 -131929 42831 -131885
rect 42887 -131929 42931 -131885
rect 43387 -131929 43431 -131885
rect 43487 -131929 43531 -131885
rect 43587 -131929 43631 -131885
rect 43687 -131929 43731 -131885
rect 43787 -131929 43831 -131885
rect 43887 -131929 43931 -131885
rect 43987 -131929 44031 -131885
rect 44087 -131929 44131 -131885
rect 44187 -131929 44231 -131885
rect 44287 -131929 44331 -131885
rect 44387 -131929 44431 -131885
rect 44487 -131929 44531 -131885
rect 44587 -131929 44631 -131885
rect 44687 -131929 44731 -131885
rect 44787 -131929 44831 -131885
rect 44887 -131929 44931 -131885
rect -13354 -131995 -13310 -131951
rect -13254 -131995 -13210 -131951
rect -13154 -131995 -13110 -131951
rect -13054 -131995 -13010 -131951
rect -12954 -131995 -12910 -131951
rect -12854 -131995 -12810 -131951
rect -12754 -131995 -12710 -131951
rect -12654 -131995 -12610 -131951
rect -12554 -131995 -12510 -131951
rect -12454 -131995 -12410 -131951
rect -12354 -131995 -12310 -131951
rect -12254 -131995 -12210 -131951
rect -12154 -131995 -12110 -131951
rect -12054 -131995 -12010 -131951
rect -11954 -131995 -11910 -131951
rect -11854 -131995 -11810 -131951
rect -11354 -131995 -11310 -131951
rect -11254 -131995 -11210 -131951
rect -11154 -131995 -11110 -131951
rect -11054 -131995 -11010 -131951
rect -10954 -131995 -10910 -131951
rect -10854 -131995 -10810 -131951
rect -10754 -131995 -10710 -131951
rect -10654 -131995 -10610 -131951
rect -10554 -131995 -10510 -131951
rect -10454 -131995 -10410 -131951
rect -10354 -131995 -10310 -131951
rect -10254 -131995 -10210 -131951
rect -10154 -131995 -10110 -131951
rect -10054 -131995 -10010 -131951
rect -9954 -131995 -9910 -131951
rect -9854 -131995 -9810 -131951
rect -9354 -131995 -9310 -131951
rect -9254 -131995 -9210 -131951
rect -9154 -131995 -9110 -131951
rect -9054 -131995 -9010 -131951
rect -8954 -131995 -8910 -131951
rect -8854 -131995 -8810 -131951
rect -8754 -131995 -8710 -131951
rect -8654 -131995 -8610 -131951
rect -8554 -131995 -8510 -131951
rect -8454 -131995 -8410 -131951
rect -8354 -131995 -8310 -131951
rect -8254 -131995 -8210 -131951
rect -8154 -131995 -8110 -131951
rect -8054 -131995 -8010 -131951
rect -7954 -131995 -7910 -131951
rect -7854 -131995 -7810 -131951
rect -7354 -131995 -7310 -131951
rect -7254 -131995 -7210 -131951
rect -7154 -131995 -7110 -131951
rect -7054 -131995 -7010 -131951
rect -6954 -131995 -6910 -131951
rect -6854 -131995 -6810 -131951
rect -6754 -131995 -6710 -131951
rect -6654 -131995 -6610 -131951
rect -6554 -131995 -6510 -131951
rect -6454 -131995 -6410 -131951
rect -6354 -131995 -6310 -131951
rect -6254 -131995 -6210 -131951
rect -6154 -131995 -6110 -131951
rect -6054 -131995 -6010 -131951
rect -5954 -131995 -5910 -131951
rect -5854 -131995 -5810 -131951
rect 37387 -132029 37431 -131985
rect 37487 -132029 37531 -131985
rect 37587 -132029 37631 -131985
rect 37687 -132029 37731 -131985
rect 37787 -132029 37831 -131985
rect 37887 -132029 37931 -131985
rect 37987 -132029 38031 -131985
rect 38087 -132029 38131 -131985
rect 38187 -132029 38231 -131985
rect 38287 -132029 38331 -131985
rect 38387 -132029 38431 -131985
rect 38487 -132029 38531 -131985
rect 38587 -132029 38631 -131985
rect 38687 -132029 38731 -131985
rect 38787 -132029 38831 -131985
rect 38887 -132029 38931 -131985
rect 39387 -132029 39431 -131985
rect 39487 -132029 39531 -131985
rect 39587 -132029 39631 -131985
rect 39687 -132029 39731 -131985
rect 39787 -132029 39831 -131985
rect 39887 -132029 39931 -131985
rect 39987 -132029 40031 -131985
rect 40087 -132029 40131 -131985
rect 40187 -132029 40231 -131985
rect 40287 -132029 40331 -131985
rect 40387 -132029 40431 -131985
rect 40487 -132029 40531 -131985
rect 40587 -132029 40631 -131985
rect 40687 -132029 40731 -131985
rect 40787 -132029 40831 -131985
rect 40887 -132029 40931 -131985
rect 41387 -132029 41431 -131985
rect 41487 -132029 41531 -131985
rect 41587 -132029 41631 -131985
rect 41687 -132029 41731 -131985
rect 41787 -132029 41831 -131985
rect 41887 -132029 41931 -131985
rect 41987 -132029 42031 -131985
rect 42087 -132029 42131 -131985
rect 42187 -132029 42231 -131985
rect 42287 -132029 42331 -131985
rect 42387 -132029 42431 -131985
rect 42487 -132029 42531 -131985
rect 42587 -132029 42631 -131985
rect 42687 -132029 42731 -131985
rect 42787 -132029 42831 -131985
rect 42887 -132029 42931 -131985
rect 43387 -132029 43431 -131985
rect 43487 -132029 43531 -131985
rect 43587 -132029 43631 -131985
rect 43687 -132029 43731 -131985
rect 43787 -132029 43831 -131985
rect 43887 -132029 43931 -131985
rect 43987 -132029 44031 -131985
rect 44087 -132029 44131 -131985
rect 44187 -132029 44231 -131985
rect 44287 -132029 44331 -131985
rect 44387 -132029 44431 -131985
rect 44487 -132029 44531 -131985
rect 44587 -132029 44631 -131985
rect 44687 -132029 44731 -131985
rect 44787 -132029 44831 -131985
rect 44887 -132029 44931 -131985
rect -13354 -132095 -13310 -132051
rect -13254 -132095 -13210 -132051
rect -13154 -132095 -13110 -132051
rect -13054 -132095 -13010 -132051
rect -12954 -132095 -12910 -132051
rect -12854 -132095 -12810 -132051
rect -12754 -132095 -12710 -132051
rect -12654 -132095 -12610 -132051
rect -12554 -132095 -12510 -132051
rect -12454 -132095 -12410 -132051
rect -12354 -132095 -12310 -132051
rect -12254 -132095 -12210 -132051
rect -12154 -132095 -12110 -132051
rect -12054 -132095 -12010 -132051
rect -11954 -132095 -11910 -132051
rect -11854 -132095 -11810 -132051
rect -11354 -132095 -11310 -132051
rect -11254 -132095 -11210 -132051
rect -11154 -132095 -11110 -132051
rect -11054 -132095 -11010 -132051
rect -10954 -132095 -10910 -132051
rect -10854 -132095 -10810 -132051
rect -10754 -132095 -10710 -132051
rect -10654 -132095 -10610 -132051
rect -10554 -132095 -10510 -132051
rect -10454 -132095 -10410 -132051
rect -10354 -132095 -10310 -132051
rect -10254 -132095 -10210 -132051
rect -10154 -132095 -10110 -132051
rect -10054 -132095 -10010 -132051
rect -9954 -132095 -9910 -132051
rect -9854 -132095 -9810 -132051
rect -9354 -132095 -9310 -132051
rect -9254 -132095 -9210 -132051
rect -9154 -132095 -9110 -132051
rect -9054 -132095 -9010 -132051
rect -8954 -132095 -8910 -132051
rect -8854 -132095 -8810 -132051
rect -8754 -132095 -8710 -132051
rect -8654 -132095 -8610 -132051
rect -8554 -132095 -8510 -132051
rect -8454 -132095 -8410 -132051
rect -8354 -132095 -8310 -132051
rect -8254 -132095 -8210 -132051
rect -8154 -132095 -8110 -132051
rect -8054 -132095 -8010 -132051
rect -7954 -132095 -7910 -132051
rect -7854 -132095 -7810 -132051
rect -7354 -132095 -7310 -132051
rect -7254 -132095 -7210 -132051
rect -7154 -132095 -7110 -132051
rect -7054 -132095 -7010 -132051
rect -6954 -132095 -6910 -132051
rect -6854 -132095 -6810 -132051
rect -6754 -132095 -6710 -132051
rect -6654 -132095 -6610 -132051
rect -6554 -132095 -6510 -132051
rect -6454 -132095 -6410 -132051
rect -6354 -132095 -6310 -132051
rect -6254 -132095 -6210 -132051
rect -6154 -132095 -6110 -132051
rect -6054 -132095 -6010 -132051
rect -5954 -132095 -5910 -132051
rect -5854 -132095 -5810 -132051
rect 37387 -132129 37431 -132085
rect 37487 -132129 37531 -132085
rect 37587 -132129 37631 -132085
rect 37687 -132129 37731 -132085
rect 37787 -132129 37831 -132085
rect 37887 -132129 37931 -132085
rect 37987 -132129 38031 -132085
rect 38087 -132129 38131 -132085
rect 38187 -132129 38231 -132085
rect 38287 -132129 38331 -132085
rect 38387 -132129 38431 -132085
rect 38487 -132129 38531 -132085
rect 38587 -132129 38631 -132085
rect 38687 -132129 38731 -132085
rect 38787 -132129 38831 -132085
rect 38887 -132129 38931 -132085
rect 39387 -132129 39431 -132085
rect 39487 -132129 39531 -132085
rect 39587 -132129 39631 -132085
rect 39687 -132129 39731 -132085
rect 39787 -132129 39831 -132085
rect 39887 -132129 39931 -132085
rect 39987 -132129 40031 -132085
rect 40087 -132129 40131 -132085
rect 40187 -132129 40231 -132085
rect 40287 -132129 40331 -132085
rect 40387 -132129 40431 -132085
rect 40487 -132129 40531 -132085
rect 40587 -132129 40631 -132085
rect 40687 -132129 40731 -132085
rect 40787 -132129 40831 -132085
rect 40887 -132129 40931 -132085
rect 41387 -132129 41431 -132085
rect 41487 -132129 41531 -132085
rect 41587 -132129 41631 -132085
rect 41687 -132129 41731 -132085
rect 41787 -132129 41831 -132085
rect 41887 -132129 41931 -132085
rect 41987 -132129 42031 -132085
rect 42087 -132129 42131 -132085
rect 42187 -132129 42231 -132085
rect 42287 -132129 42331 -132085
rect 42387 -132129 42431 -132085
rect 42487 -132129 42531 -132085
rect 42587 -132129 42631 -132085
rect 42687 -132129 42731 -132085
rect 42787 -132129 42831 -132085
rect 42887 -132129 42931 -132085
rect 43387 -132129 43431 -132085
rect 43487 -132129 43531 -132085
rect 43587 -132129 43631 -132085
rect 43687 -132129 43731 -132085
rect 43787 -132129 43831 -132085
rect 43887 -132129 43931 -132085
rect 43987 -132129 44031 -132085
rect 44087 -132129 44131 -132085
rect 44187 -132129 44231 -132085
rect 44287 -132129 44331 -132085
rect 44387 -132129 44431 -132085
rect 44487 -132129 44531 -132085
rect 44587 -132129 44631 -132085
rect 44687 -132129 44731 -132085
rect 44787 -132129 44831 -132085
rect 44887 -132129 44931 -132085
rect -13354 -132195 -13310 -132151
rect -13254 -132195 -13210 -132151
rect -13154 -132195 -13110 -132151
rect -13054 -132195 -13010 -132151
rect -12954 -132195 -12910 -132151
rect -12854 -132195 -12810 -132151
rect -12754 -132195 -12710 -132151
rect -12654 -132195 -12610 -132151
rect -12554 -132195 -12510 -132151
rect -12454 -132195 -12410 -132151
rect -12354 -132195 -12310 -132151
rect -12254 -132195 -12210 -132151
rect -12154 -132195 -12110 -132151
rect -12054 -132195 -12010 -132151
rect -11954 -132195 -11910 -132151
rect -11854 -132195 -11810 -132151
rect -11354 -132195 -11310 -132151
rect -11254 -132195 -11210 -132151
rect -11154 -132195 -11110 -132151
rect -11054 -132195 -11010 -132151
rect -10954 -132195 -10910 -132151
rect -10854 -132195 -10810 -132151
rect -10754 -132195 -10710 -132151
rect -10654 -132195 -10610 -132151
rect -10554 -132195 -10510 -132151
rect -10454 -132195 -10410 -132151
rect -10354 -132195 -10310 -132151
rect -10254 -132195 -10210 -132151
rect -10154 -132195 -10110 -132151
rect -10054 -132195 -10010 -132151
rect -9954 -132195 -9910 -132151
rect -9854 -132195 -9810 -132151
rect -9354 -132195 -9310 -132151
rect -9254 -132195 -9210 -132151
rect -9154 -132195 -9110 -132151
rect -9054 -132195 -9010 -132151
rect -8954 -132195 -8910 -132151
rect -8854 -132195 -8810 -132151
rect -8754 -132195 -8710 -132151
rect -8654 -132195 -8610 -132151
rect -8554 -132195 -8510 -132151
rect -8454 -132195 -8410 -132151
rect -8354 -132195 -8310 -132151
rect -8254 -132195 -8210 -132151
rect -8154 -132195 -8110 -132151
rect -8054 -132195 -8010 -132151
rect -7954 -132195 -7910 -132151
rect -7854 -132195 -7810 -132151
rect -7354 -132195 -7310 -132151
rect -7254 -132195 -7210 -132151
rect -7154 -132195 -7110 -132151
rect -7054 -132195 -7010 -132151
rect -6954 -132195 -6910 -132151
rect -6854 -132195 -6810 -132151
rect -6754 -132195 -6710 -132151
rect -6654 -132195 -6610 -132151
rect -6554 -132195 -6510 -132151
rect -6454 -132195 -6410 -132151
rect -6354 -132195 -6310 -132151
rect -6254 -132195 -6210 -132151
rect -6154 -132195 -6110 -132151
rect -6054 -132195 -6010 -132151
rect -5954 -132195 -5910 -132151
rect -5854 -132195 -5810 -132151
rect 37387 -132229 37431 -132185
rect 37487 -132229 37531 -132185
rect 37587 -132229 37631 -132185
rect 37687 -132229 37731 -132185
rect 37787 -132229 37831 -132185
rect 37887 -132229 37931 -132185
rect 37987 -132229 38031 -132185
rect 38087 -132229 38131 -132185
rect 38187 -132229 38231 -132185
rect 38287 -132229 38331 -132185
rect 38387 -132229 38431 -132185
rect 38487 -132229 38531 -132185
rect 38587 -132229 38631 -132185
rect 38687 -132229 38731 -132185
rect 38787 -132229 38831 -132185
rect 38887 -132229 38931 -132185
rect 39387 -132229 39431 -132185
rect 39487 -132229 39531 -132185
rect 39587 -132229 39631 -132185
rect 39687 -132229 39731 -132185
rect 39787 -132229 39831 -132185
rect 39887 -132229 39931 -132185
rect 39987 -132229 40031 -132185
rect 40087 -132229 40131 -132185
rect 40187 -132229 40231 -132185
rect 40287 -132229 40331 -132185
rect 40387 -132229 40431 -132185
rect 40487 -132229 40531 -132185
rect 40587 -132229 40631 -132185
rect 40687 -132229 40731 -132185
rect 40787 -132229 40831 -132185
rect 40887 -132229 40931 -132185
rect 41387 -132229 41431 -132185
rect 41487 -132229 41531 -132185
rect 41587 -132229 41631 -132185
rect 41687 -132229 41731 -132185
rect 41787 -132229 41831 -132185
rect 41887 -132229 41931 -132185
rect 41987 -132229 42031 -132185
rect 42087 -132229 42131 -132185
rect 42187 -132229 42231 -132185
rect 42287 -132229 42331 -132185
rect 42387 -132229 42431 -132185
rect 42487 -132229 42531 -132185
rect 42587 -132229 42631 -132185
rect 42687 -132229 42731 -132185
rect 42787 -132229 42831 -132185
rect 42887 -132229 42931 -132185
rect 43387 -132229 43431 -132185
rect 43487 -132229 43531 -132185
rect 43587 -132229 43631 -132185
rect 43687 -132229 43731 -132185
rect 43787 -132229 43831 -132185
rect 43887 -132229 43931 -132185
rect 43987 -132229 44031 -132185
rect 44087 -132229 44131 -132185
rect 44187 -132229 44231 -132185
rect 44287 -132229 44331 -132185
rect 44387 -132229 44431 -132185
rect 44487 -132229 44531 -132185
rect 44587 -132229 44631 -132185
rect 44687 -132229 44731 -132185
rect 44787 -132229 44831 -132185
rect 44887 -132229 44931 -132185
rect -13354 -132295 -13310 -132251
rect -13254 -132295 -13210 -132251
rect -13154 -132295 -13110 -132251
rect -13054 -132295 -13010 -132251
rect -12954 -132295 -12910 -132251
rect -12854 -132295 -12810 -132251
rect -12754 -132295 -12710 -132251
rect -12654 -132295 -12610 -132251
rect -12554 -132295 -12510 -132251
rect -12454 -132295 -12410 -132251
rect -12354 -132295 -12310 -132251
rect -12254 -132295 -12210 -132251
rect -12154 -132295 -12110 -132251
rect -12054 -132295 -12010 -132251
rect -11954 -132295 -11910 -132251
rect -11854 -132295 -11810 -132251
rect -11354 -132295 -11310 -132251
rect -11254 -132295 -11210 -132251
rect -11154 -132295 -11110 -132251
rect -11054 -132295 -11010 -132251
rect -10954 -132295 -10910 -132251
rect -10854 -132295 -10810 -132251
rect -10754 -132295 -10710 -132251
rect -10654 -132295 -10610 -132251
rect -10554 -132295 -10510 -132251
rect -10454 -132295 -10410 -132251
rect -10354 -132295 -10310 -132251
rect -10254 -132295 -10210 -132251
rect -10154 -132295 -10110 -132251
rect -10054 -132295 -10010 -132251
rect -9954 -132295 -9910 -132251
rect -9854 -132295 -9810 -132251
rect -9354 -132295 -9310 -132251
rect -9254 -132295 -9210 -132251
rect -9154 -132295 -9110 -132251
rect -9054 -132295 -9010 -132251
rect -8954 -132295 -8910 -132251
rect -8854 -132295 -8810 -132251
rect -8754 -132295 -8710 -132251
rect -8654 -132295 -8610 -132251
rect -8554 -132295 -8510 -132251
rect -8454 -132295 -8410 -132251
rect -8354 -132295 -8310 -132251
rect -8254 -132295 -8210 -132251
rect -8154 -132295 -8110 -132251
rect -8054 -132295 -8010 -132251
rect -7954 -132295 -7910 -132251
rect -7854 -132295 -7810 -132251
rect -7354 -132295 -7310 -132251
rect -7254 -132295 -7210 -132251
rect -7154 -132295 -7110 -132251
rect -7054 -132295 -7010 -132251
rect -6954 -132295 -6910 -132251
rect -6854 -132295 -6810 -132251
rect -6754 -132295 -6710 -132251
rect -6654 -132295 -6610 -132251
rect -6554 -132295 -6510 -132251
rect -6454 -132295 -6410 -132251
rect -6354 -132295 -6310 -132251
rect -6254 -132295 -6210 -132251
rect -6154 -132295 -6110 -132251
rect -6054 -132295 -6010 -132251
rect -5954 -132295 -5910 -132251
rect -5854 -132295 -5810 -132251
rect 37387 -132329 37431 -132285
rect 37487 -132329 37531 -132285
rect 37587 -132329 37631 -132285
rect 37687 -132329 37731 -132285
rect 37787 -132329 37831 -132285
rect 37887 -132329 37931 -132285
rect 37987 -132329 38031 -132285
rect 38087 -132329 38131 -132285
rect 38187 -132329 38231 -132285
rect 38287 -132329 38331 -132285
rect 38387 -132329 38431 -132285
rect 38487 -132329 38531 -132285
rect 38587 -132329 38631 -132285
rect 38687 -132329 38731 -132285
rect 38787 -132329 38831 -132285
rect 38887 -132329 38931 -132285
rect 39387 -132329 39431 -132285
rect 39487 -132329 39531 -132285
rect 39587 -132329 39631 -132285
rect 39687 -132329 39731 -132285
rect 39787 -132329 39831 -132285
rect 39887 -132329 39931 -132285
rect 39987 -132329 40031 -132285
rect 40087 -132329 40131 -132285
rect 40187 -132329 40231 -132285
rect 40287 -132329 40331 -132285
rect 40387 -132329 40431 -132285
rect 40487 -132329 40531 -132285
rect 40587 -132329 40631 -132285
rect 40687 -132329 40731 -132285
rect 40787 -132329 40831 -132285
rect 40887 -132329 40931 -132285
rect 41387 -132329 41431 -132285
rect 41487 -132329 41531 -132285
rect 41587 -132329 41631 -132285
rect 41687 -132329 41731 -132285
rect 41787 -132329 41831 -132285
rect 41887 -132329 41931 -132285
rect 41987 -132329 42031 -132285
rect 42087 -132329 42131 -132285
rect 42187 -132329 42231 -132285
rect 42287 -132329 42331 -132285
rect 42387 -132329 42431 -132285
rect 42487 -132329 42531 -132285
rect 42587 -132329 42631 -132285
rect 42687 -132329 42731 -132285
rect 42787 -132329 42831 -132285
rect 42887 -132329 42931 -132285
rect 43387 -132329 43431 -132285
rect 43487 -132329 43531 -132285
rect 43587 -132329 43631 -132285
rect 43687 -132329 43731 -132285
rect 43787 -132329 43831 -132285
rect 43887 -132329 43931 -132285
rect 43987 -132329 44031 -132285
rect 44087 -132329 44131 -132285
rect 44187 -132329 44231 -132285
rect 44287 -132329 44331 -132285
rect 44387 -132329 44431 -132285
rect 44487 -132329 44531 -132285
rect 44587 -132329 44631 -132285
rect 44687 -132329 44731 -132285
rect 44787 -132329 44831 -132285
rect 44887 -132329 44931 -132285
rect -13354 -132395 -13310 -132351
rect -13254 -132395 -13210 -132351
rect -13154 -132395 -13110 -132351
rect -13054 -132395 -13010 -132351
rect -12954 -132395 -12910 -132351
rect -12854 -132395 -12810 -132351
rect -12754 -132395 -12710 -132351
rect -12654 -132395 -12610 -132351
rect -12554 -132395 -12510 -132351
rect -12454 -132395 -12410 -132351
rect -12354 -132395 -12310 -132351
rect -12254 -132395 -12210 -132351
rect -12154 -132395 -12110 -132351
rect -12054 -132395 -12010 -132351
rect -11954 -132395 -11910 -132351
rect -11854 -132395 -11810 -132351
rect -11354 -132395 -11310 -132351
rect -11254 -132395 -11210 -132351
rect -11154 -132395 -11110 -132351
rect -11054 -132395 -11010 -132351
rect -10954 -132395 -10910 -132351
rect -10854 -132395 -10810 -132351
rect -10754 -132395 -10710 -132351
rect -10654 -132395 -10610 -132351
rect -10554 -132395 -10510 -132351
rect -10454 -132395 -10410 -132351
rect -10354 -132395 -10310 -132351
rect -10254 -132395 -10210 -132351
rect -10154 -132395 -10110 -132351
rect -10054 -132395 -10010 -132351
rect -9954 -132395 -9910 -132351
rect -9854 -132395 -9810 -132351
rect -9354 -132395 -9310 -132351
rect -9254 -132395 -9210 -132351
rect -9154 -132395 -9110 -132351
rect -9054 -132395 -9010 -132351
rect -8954 -132395 -8910 -132351
rect -8854 -132395 -8810 -132351
rect -8754 -132395 -8710 -132351
rect -8654 -132395 -8610 -132351
rect -8554 -132395 -8510 -132351
rect -8454 -132395 -8410 -132351
rect -8354 -132395 -8310 -132351
rect -8254 -132395 -8210 -132351
rect -8154 -132395 -8110 -132351
rect -8054 -132395 -8010 -132351
rect -7954 -132395 -7910 -132351
rect -7854 -132395 -7810 -132351
rect -7354 -132395 -7310 -132351
rect -7254 -132395 -7210 -132351
rect -7154 -132395 -7110 -132351
rect -7054 -132395 -7010 -132351
rect -6954 -132395 -6910 -132351
rect -6854 -132395 -6810 -132351
rect -6754 -132395 -6710 -132351
rect -6654 -132395 -6610 -132351
rect -6554 -132395 -6510 -132351
rect -6454 -132395 -6410 -132351
rect -6354 -132395 -6310 -132351
rect -6254 -132395 -6210 -132351
rect -6154 -132395 -6110 -132351
rect -6054 -132395 -6010 -132351
rect -5954 -132395 -5910 -132351
rect -5854 -132395 -5810 -132351
rect 37387 -132429 37431 -132385
rect 37487 -132429 37531 -132385
rect 37587 -132429 37631 -132385
rect 37687 -132429 37731 -132385
rect 37787 -132429 37831 -132385
rect 37887 -132429 37931 -132385
rect 37987 -132429 38031 -132385
rect 38087 -132429 38131 -132385
rect 38187 -132429 38231 -132385
rect 38287 -132429 38331 -132385
rect 38387 -132429 38431 -132385
rect 38487 -132429 38531 -132385
rect 38587 -132429 38631 -132385
rect 38687 -132429 38731 -132385
rect 38787 -132429 38831 -132385
rect 38887 -132429 38931 -132385
rect 39387 -132429 39431 -132385
rect 39487 -132429 39531 -132385
rect 39587 -132429 39631 -132385
rect 39687 -132429 39731 -132385
rect 39787 -132429 39831 -132385
rect 39887 -132429 39931 -132385
rect 39987 -132429 40031 -132385
rect 40087 -132429 40131 -132385
rect 40187 -132429 40231 -132385
rect 40287 -132429 40331 -132385
rect 40387 -132429 40431 -132385
rect 40487 -132429 40531 -132385
rect 40587 -132429 40631 -132385
rect 40687 -132429 40731 -132385
rect 40787 -132429 40831 -132385
rect 40887 -132429 40931 -132385
rect 41387 -132429 41431 -132385
rect 41487 -132429 41531 -132385
rect 41587 -132429 41631 -132385
rect 41687 -132429 41731 -132385
rect 41787 -132429 41831 -132385
rect 41887 -132429 41931 -132385
rect 41987 -132429 42031 -132385
rect 42087 -132429 42131 -132385
rect 42187 -132429 42231 -132385
rect 42287 -132429 42331 -132385
rect 42387 -132429 42431 -132385
rect 42487 -132429 42531 -132385
rect 42587 -132429 42631 -132385
rect 42687 -132429 42731 -132385
rect 42787 -132429 42831 -132385
rect 42887 -132429 42931 -132385
rect 43387 -132429 43431 -132385
rect 43487 -132429 43531 -132385
rect 43587 -132429 43631 -132385
rect 43687 -132429 43731 -132385
rect 43787 -132429 43831 -132385
rect 43887 -132429 43931 -132385
rect 43987 -132429 44031 -132385
rect 44087 -132429 44131 -132385
rect 44187 -132429 44231 -132385
rect 44287 -132429 44331 -132385
rect 44387 -132429 44431 -132385
rect 44487 -132429 44531 -132385
rect 44587 -132429 44631 -132385
rect 44687 -132429 44731 -132385
rect 44787 -132429 44831 -132385
rect 44887 -132429 44931 -132385
rect -13354 -132495 -13310 -132451
rect -13254 -132495 -13210 -132451
rect -13154 -132495 -13110 -132451
rect -13054 -132495 -13010 -132451
rect -12954 -132495 -12910 -132451
rect -12854 -132495 -12810 -132451
rect -12754 -132495 -12710 -132451
rect -12654 -132495 -12610 -132451
rect -12554 -132495 -12510 -132451
rect -12454 -132495 -12410 -132451
rect -12354 -132495 -12310 -132451
rect -12254 -132495 -12210 -132451
rect -12154 -132495 -12110 -132451
rect -12054 -132495 -12010 -132451
rect -11954 -132495 -11910 -132451
rect -11854 -132495 -11810 -132451
rect -11354 -132495 -11310 -132451
rect -11254 -132495 -11210 -132451
rect -11154 -132495 -11110 -132451
rect -11054 -132495 -11010 -132451
rect -10954 -132495 -10910 -132451
rect -10854 -132495 -10810 -132451
rect -10754 -132495 -10710 -132451
rect -10654 -132495 -10610 -132451
rect -10554 -132495 -10510 -132451
rect -10454 -132495 -10410 -132451
rect -10354 -132495 -10310 -132451
rect -10254 -132495 -10210 -132451
rect -10154 -132495 -10110 -132451
rect -10054 -132495 -10010 -132451
rect -9954 -132495 -9910 -132451
rect -9854 -132495 -9810 -132451
rect -9354 -132495 -9310 -132451
rect -9254 -132495 -9210 -132451
rect -9154 -132495 -9110 -132451
rect -9054 -132495 -9010 -132451
rect -8954 -132495 -8910 -132451
rect -8854 -132495 -8810 -132451
rect -8754 -132495 -8710 -132451
rect -8654 -132495 -8610 -132451
rect -8554 -132495 -8510 -132451
rect -8454 -132495 -8410 -132451
rect -8354 -132495 -8310 -132451
rect -8254 -132495 -8210 -132451
rect -8154 -132495 -8110 -132451
rect -8054 -132495 -8010 -132451
rect -7954 -132495 -7910 -132451
rect -7854 -132495 -7810 -132451
rect -7354 -132495 -7310 -132451
rect -7254 -132495 -7210 -132451
rect -7154 -132495 -7110 -132451
rect -7054 -132495 -7010 -132451
rect -6954 -132495 -6910 -132451
rect -6854 -132495 -6810 -132451
rect -6754 -132495 -6710 -132451
rect -6654 -132495 -6610 -132451
rect -6554 -132495 -6510 -132451
rect -6454 -132495 -6410 -132451
rect -6354 -132495 -6310 -132451
rect -6254 -132495 -6210 -132451
rect -6154 -132495 -6110 -132451
rect -6054 -132495 -6010 -132451
rect -5954 -132495 -5910 -132451
rect -5854 -132495 -5810 -132451
rect 37387 -132529 37431 -132485
rect 37487 -132529 37531 -132485
rect 37587 -132529 37631 -132485
rect 37687 -132529 37731 -132485
rect 37787 -132529 37831 -132485
rect 37887 -132529 37931 -132485
rect 37987 -132529 38031 -132485
rect 38087 -132529 38131 -132485
rect 38187 -132529 38231 -132485
rect 38287 -132529 38331 -132485
rect 38387 -132529 38431 -132485
rect 38487 -132529 38531 -132485
rect 38587 -132529 38631 -132485
rect 38687 -132529 38731 -132485
rect 38787 -132529 38831 -132485
rect 38887 -132529 38931 -132485
rect 39387 -132529 39431 -132485
rect 39487 -132529 39531 -132485
rect 39587 -132529 39631 -132485
rect 39687 -132529 39731 -132485
rect 39787 -132529 39831 -132485
rect 39887 -132529 39931 -132485
rect 39987 -132529 40031 -132485
rect 40087 -132529 40131 -132485
rect 40187 -132529 40231 -132485
rect 40287 -132529 40331 -132485
rect 40387 -132529 40431 -132485
rect 40487 -132529 40531 -132485
rect 40587 -132529 40631 -132485
rect 40687 -132529 40731 -132485
rect 40787 -132529 40831 -132485
rect 40887 -132529 40931 -132485
rect 41387 -132529 41431 -132485
rect 41487 -132529 41531 -132485
rect 41587 -132529 41631 -132485
rect 41687 -132529 41731 -132485
rect 41787 -132529 41831 -132485
rect 41887 -132529 41931 -132485
rect 41987 -132529 42031 -132485
rect 42087 -132529 42131 -132485
rect 42187 -132529 42231 -132485
rect 42287 -132529 42331 -132485
rect 42387 -132529 42431 -132485
rect 42487 -132529 42531 -132485
rect 42587 -132529 42631 -132485
rect 42687 -132529 42731 -132485
rect 42787 -132529 42831 -132485
rect 42887 -132529 42931 -132485
rect 43387 -132529 43431 -132485
rect 43487 -132529 43531 -132485
rect 43587 -132529 43631 -132485
rect 43687 -132529 43731 -132485
rect 43787 -132529 43831 -132485
rect 43887 -132529 43931 -132485
rect 43987 -132529 44031 -132485
rect 44087 -132529 44131 -132485
rect 44187 -132529 44231 -132485
rect 44287 -132529 44331 -132485
rect 44387 -132529 44431 -132485
rect 44487 -132529 44531 -132485
rect 44587 -132529 44631 -132485
rect 44687 -132529 44731 -132485
rect 44787 -132529 44831 -132485
rect 44887 -132529 44931 -132485
rect -13354 -132595 -13310 -132551
rect -13254 -132595 -13210 -132551
rect -13154 -132595 -13110 -132551
rect -13054 -132595 -13010 -132551
rect -12954 -132595 -12910 -132551
rect -12854 -132595 -12810 -132551
rect -12754 -132595 -12710 -132551
rect -12654 -132595 -12610 -132551
rect -12554 -132595 -12510 -132551
rect -12454 -132595 -12410 -132551
rect -12354 -132595 -12310 -132551
rect -12254 -132595 -12210 -132551
rect -12154 -132595 -12110 -132551
rect -12054 -132595 -12010 -132551
rect -11954 -132595 -11910 -132551
rect -11854 -132595 -11810 -132551
rect -11354 -132595 -11310 -132551
rect -11254 -132595 -11210 -132551
rect -11154 -132595 -11110 -132551
rect -11054 -132595 -11010 -132551
rect -10954 -132595 -10910 -132551
rect -10854 -132595 -10810 -132551
rect -10754 -132595 -10710 -132551
rect -10654 -132595 -10610 -132551
rect -10554 -132595 -10510 -132551
rect -10454 -132595 -10410 -132551
rect -10354 -132595 -10310 -132551
rect -10254 -132595 -10210 -132551
rect -10154 -132595 -10110 -132551
rect -10054 -132595 -10010 -132551
rect -9954 -132595 -9910 -132551
rect -9854 -132595 -9810 -132551
rect -9354 -132595 -9310 -132551
rect -9254 -132595 -9210 -132551
rect -9154 -132595 -9110 -132551
rect -9054 -132595 -9010 -132551
rect -8954 -132595 -8910 -132551
rect -8854 -132595 -8810 -132551
rect -8754 -132595 -8710 -132551
rect -8654 -132595 -8610 -132551
rect -8554 -132595 -8510 -132551
rect -8454 -132595 -8410 -132551
rect -8354 -132595 -8310 -132551
rect -8254 -132595 -8210 -132551
rect -8154 -132595 -8110 -132551
rect -8054 -132595 -8010 -132551
rect -7954 -132595 -7910 -132551
rect -7854 -132595 -7810 -132551
rect -7354 -132595 -7310 -132551
rect -7254 -132595 -7210 -132551
rect -7154 -132595 -7110 -132551
rect -7054 -132595 -7010 -132551
rect -6954 -132595 -6910 -132551
rect -6854 -132595 -6810 -132551
rect -6754 -132595 -6710 -132551
rect -6654 -132595 -6610 -132551
rect -6554 -132595 -6510 -132551
rect -6454 -132595 -6410 -132551
rect -6354 -132595 -6310 -132551
rect -6254 -132595 -6210 -132551
rect -6154 -132595 -6110 -132551
rect -6054 -132595 -6010 -132551
rect -5954 -132595 -5910 -132551
rect -5854 -132595 -5810 -132551
rect 37387 -132629 37431 -132585
rect 37487 -132629 37531 -132585
rect 37587 -132629 37631 -132585
rect 37687 -132629 37731 -132585
rect 37787 -132629 37831 -132585
rect 37887 -132629 37931 -132585
rect 37987 -132629 38031 -132585
rect 38087 -132629 38131 -132585
rect 38187 -132629 38231 -132585
rect 38287 -132629 38331 -132585
rect 38387 -132629 38431 -132585
rect 38487 -132629 38531 -132585
rect 38587 -132629 38631 -132585
rect 38687 -132629 38731 -132585
rect 38787 -132629 38831 -132585
rect 38887 -132629 38931 -132585
rect 39387 -132629 39431 -132585
rect 39487 -132629 39531 -132585
rect 39587 -132629 39631 -132585
rect 39687 -132629 39731 -132585
rect 39787 -132629 39831 -132585
rect 39887 -132629 39931 -132585
rect 39987 -132629 40031 -132585
rect 40087 -132629 40131 -132585
rect 40187 -132629 40231 -132585
rect 40287 -132629 40331 -132585
rect 40387 -132629 40431 -132585
rect 40487 -132629 40531 -132585
rect 40587 -132629 40631 -132585
rect 40687 -132629 40731 -132585
rect 40787 -132629 40831 -132585
rect 40887 -132629 40931 -132585
rect 41387 -132629 41431 -132585
rect 41487 -132629 41531 -132585
rect 41587 -132629 41631 -132585
rect 41687 -132629 41731 -132585
rect 41787 -132629 41831 -132585
rect 41887 -132629 41931 -132585
rect 41987 -132629 42031 -132585
rect 42087 -132629 42131 -132585
rect 42187 -132629 42231 -132585
rect 42287 -132629 42331 -132585
rect 42387 -132629 42431 -132585
rect 42487 -132629 42531 -132585
rect 42587 -132629 42631 -132585
rect 42687 -132629 42731 -132585
rect 42787 -132629 42831 -132585
rect 42887 -132629 42931 -132585
rect 43387 -132629 43431 -132585
rect 43487 -132629 43531 -132585
rect 43587 -132629 43631 -132585
rect 43687 -132629 43731 -132585
rect 43787 -132629 43831 -132585
rect 43887 -132629 43931 -132585
rect 43987 -132629 44031 -132585
rect 44087 -132629 44131 -132585
rect 44187 -132629 44231 -132585
rect 44287 -132629 44331 -132585
rect 44387 -132629 44431 -132585
rect 44487 -132629 44531 -132585
rect 44587 -132629 44631 -132585
rect 44687 -132629 44731 -132585
rect 44787 -132629 44831 -132585
rect 44887 -132629 44931 -132585
rect -13354 -132695 -13310 -132651
rect -13254 -132695 -13210 -132651
rect -13154 -132695 -13110 -132651
rect -13054 -132695 -13010 -132651
rect -12954 -132695 -12910 -132651
rect -12854 -132695 -12810 -132651
rect -12754 -132695 -12710 -132651
rect -12654 -132695 -12610 -132651
rect -12554 -132695 -12510 -132651
rect -12454 -132695 -12410 -132651
rect -12354 -132695 -12310 -132651
rect -12254 -132695 -12210 -132651
rect -12154 -132695 -12110 -132651
rect -12054 -132695 -12010 -132651
rect -11954 -132695 -11910 -132651
rect -11854 -132695 -11810 -132651
rect -11354 -132695 -11310 -132651
rect -11254 -132695 -11210 -132651
rect -11154 -132695 -11110 -132651
rect -11054 -132695 -11010 -132651
rect -10954 -132695 -10910 -132651
rect -10854 -132695 -10810 -132651
rect -10754 -132695 -10710 -132651
rect -10654 -132695 -10610 -132651
rect -10554 -132695 -10510 -132651
rect -10454 -132695 -10410 -132651
rect -10354 -132695 -10310 -132651
rect -10254 -132695 -10210 -132651
rect -10154 -132695 -10110 -132651
rect -10054 -132695 -10010 -132651
rect -9954 -132695 -9910 -132651
rect -9854 -132695 -9810 -132651
rect -9354 -132695 -9310 -132651
rect -9254 -132695 -9210 -132651
rect -9154 -132695 -9110 -132651
rect -9054 -132695 -9010 -132651
rect -8954 -132695 -8910 -132651
rect -8854 -132695 -8810 -132651
rect -8754 -132695 -8710 -132651
rect -8654 -132695 -8610 -132651
rect -8554 -132695 -8510 -132651
rect -8454 -132695 -8410 -132651
rect -8354 -132695 -8310 -132651
rect -8254 -132695 -8210 -132651
rect -8154 -132695 -8110 -132651
rect -8054 -132695 -8010 -132651
rect -7954 -132695 -7910 -132651
rect -7854 -132695 -7810 -132651
rect -7354 -132695 -7310 -132651
rect -7254 -132695 -7210 -132651
rect -7154 -132695 -7110 -132651
rect -7054 -132695 -7010 -132651
rect -6954 -132695 -6910 -132651
rect -6854 -132695 -6810 -132651
rect -6754 -132695 -6710 -132651
rect -6654 -132695 -6610 -132651
rect -6554 -132695 -6510 -132651
rect -6454 -132695 -6410 -132651
rect -6354 -132695 -6310 -132651
rect -6254 -132695 -6210 -132651
rect -6154 -132695 -6110 -132651
rect -6054 -132695 -6010 -132651
rect -5954 -132695 -5910 -132651
rect -5854 -132695 -5810 -132651
rect 37387 -132729 37431 -132685
rect 37487 -132729 37531 -132685
rect 37587 -132729 37631 -132685
rect 37687 -132729 37731 -132685
rect 37787 -132729 37831 -132685
rect 37887 -132729 37931 -132685
rect 37987 -132729 38031 -132685
rect 38087 -132729 38131 -132685
rect 38187 -132729 38231 -132685
rect 38287 -132729 38331 -132685
rect 38387 -132729 38431 -132685
rect 38487 -132729 38531 -132685
rect 38587 -132729 38631 -132685
rect 38687 -132729 38731 -132685
rect 38787 -132729 38831 -132685
rect 38887 -132729 38931 -132685
rect 39387 -132729 39431 -132685
rect 39487 -132729 39531 -132685
rect 39587 -132729 39631 -132685
rect 39687 -132729 39731 -132685
rect 39787 -132729 39831 -132685
rect 39887 -132729 39931 -132685
rect 39987 -132729 40031 -132685
rect 40087 -132729 40131 -132685
rect 40187 -132729 40231 -132685
rect 40287 -132729 40331 -132685
rect 40387 -132729 40431 -132685
rect 40487 -132729 40531 -132685
rect 40587 -132729 40631 -132685
rect 40687 -132729 40731 -132685
rect 40787 -132729 40831 -132685
rect 40887 -132729 40931 -132685
rect 41387 -132729 41431 -132685
rect 41487 -132729 41531 -132685
rect 41587 -132729 41631 -132685
rect 41687 -132729 41731 -132685
rect 41787 -132729 41831 -132685
rect 41887 -132729 41931 -132685
rect 41987 -132729 42031 -132685
rect 42087 -132729 42131 -132685
rect 42187 -132729 42231 -132685
rect 42287 -132729 42331 -132685
rect 42387 -132729 42431 -132685
rect 42487 -132729 42531 -132685
rect 42587 -132729 42631 -132685
rect 42687 -132729 42731 -132685
rect 42787 -132729 42831 -132685
rect 42887 -132729 42931 -132685
rect 43387 -132729 43431 -132685
rect 43487 -132729 43531 -132685
rect 43587 -132729 43631 -132685
rect 43687 -132729 43731 -132685
rect 43787 -132729 43831 -132685
rect 43887 -132729 43931 -132685
rect 43987 -132729 44031 -132685
rect 44087 -132729 44131 -132685
rect 44187 -132729 44231 -132685
rect 44287 -132729 44331 -132685
rect 44387 -132729 44431 -132685
rect 44487 -132729 44531 -132685
rect 44587 -132729 44631 -132685
rect 44687 -132729 44731 -132685
rect 44787 -132729 44831 -132685
rect 44887 -132729 44931 -132685
rect -13354 -132795 -13310 -132751
rect -13254 -132795 -13210 -132751
rect -13154 -132795 -13110 -132751
rect -13054 -132795 -13010 -132751
rect -12954 -132795 -12910 -132751
rect -12854 -132795 -12810 -132751
rect -12754 -132795 -12710 -132751
rect -12654 -132795 -12610 -132751
rect -12554 -132795 -12510 -132751
rect -12454 -132795 -12410 -132751
rect -12354 -132795 -12310 -132751
rect -12254 -132795 -12210 -132751
rect -12154 -132795 -12110 -132751
rect -12054 -132795 -12010 -132751
rect -11954 -132795 -11910 -132751
rect -11854 -132795 -11810 -132751
rect -11354 -132795 -11310 -132751
rect -11254 -132795 -11210 -132751
rect -11154 -132795 -11110 -132751
rect -11054 -132795 -11010 -132751
rect -10954 -132795 -10910 -132751
rect -10854 -132795 -10810 -132751
rect -10754 -132795 -10710 -132751
rect -10654 -132795 -10610 -132751
rect -10554 -132795 -10510 -132751
rect -10454 -132795 -10410 -132751
rect -10354 -132795 -10310 -132751
rect -10254 -132795 -10210 -132751
rect -10154 -132795 -10110 -132751
rect -10054 -132795 -10010 -132751
rect -9954 -132795 -9910 -132751
rect -9854 -132795 -9810 -132751
rect -9354 -132795 -9310 -132751
rect -9254 -132795 -9210 -132751
rect -9154 -132795 -9110 -132751
rect -9054 -132795 -9010 -132751
rect -8954 -132795 -8910 -132751
rect -8854 -132795 -8810 -132751
rect -8754 -132795 -8710 -132751
rect -8654 -132795 -8610 -132751
rect -8554 -132795 -8510 -132751
rect -8454 -132795 -8410 -132751
rect -8354 -132795 -8310 -132751
rect -8254 -132795 -8210 -132751
rect -8154 -132795 -8110 -132751
rect -8054 -132795 -8010 -132751
rect -7954 -132795 -7910 -132751
rect -7854 -132795 -7810 -132751
rect -7354 -132795 -7310 -132751
rect -7254 -132795 -7210 -132751
rect -7154 -132795 -7110 -132751
rect -7054 -132795 -7010 -132751
rect -6954 -132795 -6910 -132751
rect -6854 -132795 -6810 -132751
rect -6754 -132795 -6710 -132751
rect -6654 -132795 -6610 -132751
rect -6554 -132795 -6510 -132751
rect -6454 -132795 -6410 -132751
rect -6354 -132795 -6310 -132751
rect -6254 -132795 -6210 -132751
rect -6154 -132795 -6110 -132751
rect -6054 -132795 -6010 -132751
rect -5954 -132795 -5910 -132751
rect -5854 -132795 -5810 -132751
rect 37387 -132829 37431 -132785
rect 37487 -132829 37531 -132785
rect 37587 -132829 37631 -132785
rect 37687 -132829 37731 -132785
rect 37787 -132829 37831 -132785
rect 37887 -132829 37931 -132785
rect 37987 -132829 38031 -132785
rect 38087 -132829 38131 -132785
rect 38187 -132829 38231 -132785
rect 38287 -132829 38331 -132785
rect 38387 -132829 38431 -132785
rect 38487 -132829 38531 -132785
rect 38587 -132829 38631 -132785
rect 38687 -132829 38731 -132785
rect 38787 -132829 38831 -132785
rect 38887 -132829 38931 -132785
rect 39387 -132829 39431 -132785
rect 39487 -132829 39531 -132785
rect 39587 -132829 39631 -132785
rect 39687 -132829 39731 -132785
rect 39787 -132829 39831 -132785
rect 39887 -132829 39931 -132785
rect 39987 -132829 40031 -132785
rect 40087 -132829 40131 -132785
rect 40187 -132829 40231 -132785
rect 40287 -132829 40331 -132785
rect 40387 -132829 40431 -132785
rect 40487 -132829 40531 -132785
rect 40587 -132829 40631 -132785
rect 40687 -132829 40731 -132785
rect 40787 -132829 40831 -132785
rect 40887 -132829 40931 -132785
rect 41387 -132829 41431 -132785
rect 41487 -132829 41531 -132785
rect 41587 -132829 41631 -132785
rect 41687 -132829 41731 -132785
rect 41787 -132829 41831 -132785
rect 41887 -132829 41931 -132785
rect 41987 -132829 42031 -132785
rect 42087 -132829 42131 -132785
rect 42187 -132829 42231 -132785
rect 42287 -132829 42331 -132785
rect 42387 -132829 42431 -132785
rect 42487 -132829 42531 -132785
rect 42587 -132829 42631 -132785
rect 42687 -132829 42731 -132785
rect 42787 -132829 42831 -132785
rect 42887 -132829 42931 -132785
rect 43387 -132829 43431 -132785
rect 43487 -132829 43531 -132785
rect 43587 -132829 43631 -132785
rect 43687 -132829 43731 -132785
rect 43787 -132829 43831 -132785
rect 43887 -132829 43931 -132785
rect 43987 -132829 44031 -132785
rect 44087 -132829 44131 -132785
rect 44187 -132829 44231 -132785
rect 44287 -132829 44331 -132785
rect 44387 -132829 44431 -132785
rect 44487 -132829 44531 -132785
rect 44587 -132829 44631 -132785
rect 44687 -132829 44731 -132785
rect 44787 -132829 44831 -132785
rect 44887 -132829 44931 -132785
rect 37387 -132929 37431 -132885
rect 37487 -132929 37531 -132885
rect 37587 -132929 37631 -132885
rect 37687 -132929 37731 -132885
rect 37787 -132929 37831 -132885
rect 37887 -132929 37931 -132885
rect 37987 -132929 38031 -132885
rect 38087 -132929 38131 -132885
rect 38187 -132929 38231 -132885
rect 38287 -132929 38331 -132885
rect 38387 -132929 38431 -132885
rect 38487 -132929 38531 -132885
rect 38587 -132929 38631 -132885
rect 38687 -132929 38731 -132885
rect 38787 -132929 38831 -132885
rect 38887 -132929 38931 -132885
rect 39387 -132929 39431 -132885
rect 39487 -132929 39531 -132885
rect 39587 -132929 39631 -132885
rect 39687 -132929 39731 -132885
rect 39787 -132929 39831 -132885
rect 39887 -132929 39931 -132885
rect 39987 -132929 40031 -132885
rect 40087 -132929 40131 -132885
rect 40187 -132929 40231 -132885
rect 40287 -132929 40331 -132885
rect 40387 -132929 40431 -132885
rect 40487 -132929 40531 -132885
rect 40587 -132929 40631 -132885
rect 40687 -132929 40731 -132885
rect 40787 -132929 40831 -132885
rect 40887 -132929 40931 -132885
rect 41387 -132929 41431 -132885
rect 41487 -132929 41531 -132885
rect 41587 -132929 41631 -132885
rect 41687 -132929 41731 -132885
rect 41787 -132929 41831 -132885
rect 41887 -132929 41931 -132885
rect 41987 -132929 42031 -132885
rect 42087 -132929 42131 -132885
rect 42187 -132929 42231 -132885
rect 42287 -132929 42331 -132885
rect 42387 -132929 42431 -132885
rect 42487 -132929 42531 -132885
rect 42587 -132929 42631 -132885
rect 42687 -132929 42731 -132885
rect 42787 -132929 42831 -132885
rect 42887 -132929 42931 -132885
rect 43387 -132929 43431 -132885
rect 43487 -132929 43531 -132885
rect 43587 -132929 43631 -132885
rect 43687 -132929 43731 -132885
rect 43787 -132929 43831 -132885
rect 43887 -132929 43931 -132885
rect 43987 -132929 44031 -132885
rect 44087 -132929 44131 -132885
rect 44187 -132929 44231 -132885
rect 44287 -132929 44331 -132885
rect 44387 -132929 44431 -132885
rect 44487 -132929 44531 -132885
rect 44587 -132929 44631 -132885
rect 44687 -132929 44731 -132885
rect 44787 -132929 44831 -132885
rect 44887 -132929 44931 -132885
rect -104783 -135358 -104739 -135314
rect -104683 -135358 -104639 -135314
rect -104583 -135358 -104539 -135314
rect -104483 -135358 -104439 -135314
rect -104383 -135358 -104339 -135314
rect -104283 -135358 -104239 -135314
rect -104183 -135358 -104139 -135314
rect -104083 -135358 -104039 -135314
rect -103983 -135358 -103939 -135314
rect -103883 -135358 -103839 -135314
rect -103783 -135358 -103739 -135314
rect -103683 -135358 -103639 -135314
rect -103583 -135358 -103539 -135314
rect -103483 -135358 -103439 -135314
rect -103383 -135358 -103339 -135314
rect -103283 -135358 -103239 -135314
rect -102783 -135358 -102739 -135314
rect -102683 -135358 -102639 -135314
rect -102583 -135358 -102539 -135314
rect -102483 -135358 -102439 -135314
rect -102383 -135358 -102339 -135314
rect -102283 -135358 -102239 -135314
rect -102183 -135358 -102139 -135314
rect -102083 -135358 -102039 -135314
rect -101983 -135358 -101939 -135314
rect -101883 -135358 -101839 -135314
rect -101783 -135358 -101739 -135314
rect -101683 -135358 -101639 -135314
rect -101583 -135358 -101539 -135314
rect -101483 -135358 -101439 -135314
rect -101383 -135358 -101339 -135314
rect -101283 -135358 -101239 -135314
rect -100783 -135358 -100739 -135314
rect -100683 -135358 -100639 -135314
rect -100583 -135358 -100539 -135314
rect -100483 -135358 -100439 -135314
rect -100383 -135358 -100339 -135314
rect -100283 -135358 -100239 -135314
rect -100183 -135358 -100139 -135314
rect -100083 -135358 -100039 -135314
rect -99983 -135358 -99939 -135314
rect -99883 -135358 -99839 -135314
rect -99783 -135358 -99739 -135314
rect -99683 -135358 -99639 -135314
rect -99583 -135358 -99539 -135314
rect -99483 -135358 -99439 -135314
rect -99383 -135358 -99339 -135314
rect -99283 -135358 -99239 -135314
rect -98783 -135358 -98739 -135314
rect -98683 -135358 -98639 -135314
rect -98583 -135358 -98539 -135314
rect -98483 -135358 -98439 -135314
rect -98383 -135358 -98339 -135314
rect -98283 -135358 -98239 -135314
rect -98183 -135358 -98139 -135314
rect -98083 -135358 -98039 -135314
rect -97983 -135358 -97939 -135314
rect -97883 -135358 -97839 -135314
rect -97783 -135358 -97739 -135314
rect -97683 -135358 -97639 -135314
rect -97583 -135358 -97539 -135314
rect -97483 -135358 -97439 -135314
rect -97383 -135358 -97339 -135314
rect -97283 -135358 -97239 -135314
rect -104783 -135458 -104739 -135414
rect -104683 -135458 -104639 -135414
rect -104583 -135458 -104539 -135414
rect -104483 -135458 -104439 -135414
rect -104383 -135458 -104339 -135414
rect -104283 -135458 -104239 -135414
rect -104183 -135458 -104139 -135414
rect -104083 -135458 -104039 -135414
rect -103983 -135458 -103939 -135414
rect -103883 -135458 -103839 -135414
rect -103783 -135458 -103739 -135414
rect -103683 -135458 -103639 -135414
rect -103583 -135458 -103539 -135414
rect -103483 -135458 -103439 -135414
rect -103383 -135458 -103339 -135414
rect -103283 -135458 -103239 -135414
rect -102783 -135458 -102739 -135414
rect -102683 -135458 -102639 -135414
rect -102583 -135458 -102539 -135414
rect -102483 -135458 -102439 -135414
rect -102383 -135458 -102339 -135414
rect -102283 -135458 -102239 -135414
rect -102183 -135458 -102139 -135414
rect -102083 -135458 -102039 -135414
rect -101983 -135458 -101939 -135414
rect -101883 -135458 -101839 -135414
rect -101783 -135458 -101739 -135414
rect -101683 -135458 -101639 -135414
rect -101583 -135458 -101539 -135414
rect -101483 -135458 -101439 -135414
rect -101383 -135458 -101339 -135414
rect -101283 -135458 -101239 -135414
rect -100783 -135458 -100739 -135414
rect -100683 -135458 -100639 -135414
rect -100583 -135458 -100539 -135414
rect -100483 -135458 -100439 -135414
rect -100383 -135458 -100339 -135414
rect -100283 -135458 -100239 -135414
rect -100183 -135458 -100139 -135414
rect -100083 -135458 -100039 -135414
rect -99983 -135458 -99939 -135414
rect -99883 -135458 -99839 -135414
rect -99783 -135458 -99739 -135414
rect -99683 -135458 -99639 -135414
rect -99583 -135458 -99539 -135414
rect -99483 -135458 -99439 -135414
rect -99383 -135458 -99339 -135414
rect -99283 -135458 -99239 -135414
rect -98783 -135458 -98739 -135414
rect -98683 -135458 -98639 -135414
rect -98583 -135458 -98539 -135414
rect -98483 -135458 -98439 -135414
rect -98383 -135458 -98339 -135414
rect -98283 -135458 -98239 -135414
rect -98183 -135458 -98139 -135414
rect -98083 -135458 -98039 -135414
rect -97983 -135458 -97939 -135414
rect -97883 -135458 -97839 -135414
rect -97783 -135458 -97739 -135414
rect -97683 -135458 -97639 -135414
rect -97583 -135458 -97539 -135414
rect -97483 -135458 -97439 -135414
rect -97383 -135458 -97339 -135414
rect -97283 -135458 -97239 -135414
rect -104783 -135558 -104739 -135514
rect -104683 -135558 -104639 -135514
rect -104583 -135558 -104539 -135514
rect -104483 -135558 -104439 -135514
rect -104383 -135558 -104339 -135514
rect -104283 -135558 -104239 -135514
rect -104183 -135558 -104139 -135514
rect -104083 -135558 -104039 -135514
rect -103983 -135558 -103939 -135514
rect -103883 -135558 -103839 -135514
rect -103783 -135558 -103739 -135514
rect -103683 -135558 -103639 -135514
rect -103583 -135558 -103539 -135514
rect -103483 -135558 -103439 -135514
rect -103383 -135558 -103339 -135514
rect -103283 -135558 -103239 -135514
rect -102783 -135558 -102739 -135514
rect -102683 -135558 -102639 -135514
rect -102583 -135558 -102539 -135514
rect -102483 -135558 -102439 -135514
rect -102383 -135558 -102339 -135514
rect -102283 -135558 -102239 -135514
rect -102183 -135558 -102139 -135514
rect -102083 -135558 -102039 -135514
rect -101983 -135558 -101939 -135514
rect -101883 -135558 -101839 -135514
rect -101783 -135558 -101739 -135514
rect -101683 -135558 -101639 -135514
rect -101583 -135558 -101539 -135514
rect -101483 -135558 -101439 -135514
rect -101383 -135558 -101339 -135514
rect -101283 -135558 -101239 -135514
rect -100783 -135558 -100739 -135514
rect -100683 -135558 -100639 -135514
rect -100583 -135558 -100539 -135514
rect -100483 -135558 -100439 -135514
rect -100383 -135558 -100339 -135514
rect -100283 -135558 -100239 -135514
rect -100183 -135558 -100139 -135514
rect -100083 -135558 -100039 -135514
rect -99983 -135558 -99939 -135514
rect -99883 -135558 -99839 -135514
rect -99783 -135558 -99739 -135514
rect -99683 -135558 -99639 -135514
rect -99583 -135558 -99539 -135514
rect -99483 -135558 -99439 -135514
rect -99383 -135558 -99339 -135514
rect -99283 -135558 -99239 -135514
rect -98783 -135558 -98739 -135514
rect -98683 -135558 -98639 -135514
rect -98583 -135558 -98539 -135514
rect -98483 -135558 -98439 -135514
rect -98383 -135558 -98339 -135514
rect -98283 -135558 -98239 -135514
rect -98183 -135558 -98139 -135514
rect -98083 -135558 -98039 -135514
rect -97983 -135558 -97939 -135514
rect -97883 -135558 -97839 -135514
rect -97783 -135558 -97739 -135514
rect -97683 -135558 -97639 -135514
rect -97583 -135558 -97539 -135514
rect -97483 -135558 -97439 -135514
rect -97383 -135558 -97339 -135514
rect -97283 -135558 -97239 -135514
rect -104783 -135658 -104739 -135614
rect -104683 -135658 -104639 -135614
rect -104583 -135658 -104539 -135614
rect -104483 -135658 -104439 -135614
rect -104383 -135658 -104339 -135614
rect -104283 -135658 -104239 -135614
rect -104183 -135658 -104139 -135614
rect -104083 -135658 -104039 -135614
rect -103983 -135658 -103939 -135614
rect -103883 -135658 -103839 -135614
rect -103783 -135658 -103739 -135614
rect -103683 -135658 -103639 -135614
rect -103583 -135658 -103539 -135614
rect -103483 -135658 -103439 -135614
rect -103383 -135658 -103339 -135614
rect -103283 -135658 -103239 -135614
rect -102783 -135658 -102739 -135614
rect -102683 -135658 -102639 -135614
rect -102583 -135658 -102539 -135614
rect -102483 -135658 -102439 -135614
rect -102383 -135658 -102339 -135614
rect -102283 -135658 -102239 -135614
rect -102183 -135658 -102139 -135614
rect -102083 -135658 -102039 -135614
rect -101983 -135658 -101939 -135614
rect -101883 -135658 -101839 -135614
rect -101783 -135658 -101739 -135614
rect -101683 -135658 -101639 -135614
rect -101583 -135658 -101539 -135614
rect -101483 -135658 -101439 -135614
rect -101383 -135658 -101339 -135614
rect -101283 -135658 -101239 -135614
rect -100783 -135658 -100739 -135614
rect -100683 -135658 -100639 -135614
rect -100583 -135658 -100539 -135614
rect -100483 -135658 -100439 -135614
rect -100383 -135658 -100339 -135614
rect -100283 -135658 -100239 -135614
rect -100183 -135658 -100139 -135614
rect -100083 -135658 -100039 -135614
rect -99983 -135658 -99939 -135614
rect -99883 -135658 -99839 -135614
rect -99783 -135658 -99739 -135614
rect -99683 -135658 -99639 -135614
rect -99583 -135658 -99539 -135614
rect -99483 -135658 -99439 -135614
rect -99383 -135658 -99339 -135614
rect -99283 -135658 -99239 -135614
rect -98783 -135658 -98739 -135614
rect -98683 -135658 -98639 -135614
rect -98583 -135658 -98539 -135614
rect -98483 -135658 -98439 -135614
rect -98383 -135658 -98339 -135614
rect -98283 -135658 -98239 -135614
rect -98183 -135658 -98139 -135614
rect -98083 -135658 -98039 -135614
rect -97983 -135658 -97939 -135614
rect -97883 -135658 -97839 -135614
rect -97783 -135658 -97739 -135614
rect -97683 -135658 -97639 -135614
rect -97583 -135658 -97539 -135614
rect -97483 -135658 -97439 -135614
rect -97383 -135658 -97339 -135614
rect -97283 -135658 -97239 -135614
rect -104783 -135758 -104739 -135714
rect -104683 -135758 -104639 -135714
rect -104583 -135758 -104539 -135714
rect -104483 -135758 -104439 -135714
rect -104383 -135758 -104339 -135714
rect -104283 -135758 -104239 -135714
rect -104183 -135758 -104139 -135714
rect -104083 -135758 -104039 -135714
rect -103983 -135758 -103939 -135714
rect -103883 -135758 -103839 -135714
rect -103783 -135758 -103739 -135714
rect -103683 -135758 -103639 -135714
rect -103583 -135758 -103539 -135714
rect -103483 -135758 -103439 -135714
rect -103383 -135758 -103339 -135714
rect -103283 -135758 -103239 -135714
rect -102783 -135758 -102739 -135714
rect -102683 -135758 -102639 -135714
rect -102583 -135758 -102539 -135714
rect -102483 -135758 -102439 -135714
rect -102383 -135758 -102339 -135714
rect -102283 -135758 -102239 -135714
rect -102183 -135758 -102139 -135714
rect -102083 -135758 -102039 -135714
rect -101983 -135758 -101939 -135714
rect -101883 -135758 -101839 -135714
rect -101783 -135758 -101739 -135714
rect -101683 -135758 -101639 -135714
rect -101583 -135758 -101539 -135714
rect -101483 -135758 -101439 -135714
rect -101383 -135758 -101339 -135714
rect -101283 -135758 -101239 -135714
rect -100783 -135758 -100739 -135714
rect -100683 -135758 -100639 -135714
rect -100583 -135758 -100539 -135714
rect -100483 -135758 -100439 -135714
rect -100383 -135758 -100339 -135714
rect -100283 -135758 -100239 -135714
rect -100183 -135758 -100139 -135714
rect -100083 -135758 -100039 -135714
rect -99983 -135758 -99939 -135714
rect -99883 -135758 -99839 -135714
rect -99783 -135758 -99739 -135714
rect -99683 -135758 -99639 -135714
rect -99583 -135758 -99539 -135714
rect -99483 -135758 -99439 -135714
rect -99383 -135758 -99339 -135714
rect -99283 -135758 -99239 -135714
rect -98783 -135758 -98739 -135714
rect -98683 -135758 -98639 -135714
rect -98583 -135758 -98539 -135714
rect -98483 -135758 -98439 -135714
rect -98383 -135758 -98339 -135714
rect -98283 -135758 -98239 -135714
rect -98183 -135758 -98139 -135714
rect -98083 -135758 -98039 -135714
rect -97983 -135758 -97939 -135714
rect -97883 -135758 -97839 -135714
rect -97783 -135758 -97739 -135714
rect -97683 -135758 -97639 -135714
rect -97583 -135758 -97539 -135714
rect -97483 -135758 -97439 -135714
rect -97383 -135758 -97339 -135714
rect -97283 -135758 -97239 -135714
rect -104783 -135858 -104739 -135814
rect -104683 -135858 -104639 -135814
rect -104583 -135858 -104539 -135814
rect -104483 -135858 -104439 -135814
rect -104383 -135858 -104339 -135814
rect -104283 -135858 -104239 -135814
rect -104183 -135858 -104139 -135814
rect -104083 -135858 -104039 -135814
rect -103983 -135858 -103939 -135814
rect -103883 -135858 -103839 -135814
rect -103783 -135858 -103739 -135814
rect -103683 -135858 -103639 -135814
rect -103583 -135858 -103539 -135814
rect -103483 -135858 -103439 -135814
rect -103383 -135858 -103339 -135814
rect -103283 -135858 -103239 -135814
rect -102783 -135858 -102739 -135814
rect -102683 -135858 -102639 -135814
rect -102583 -135858 -102539 -135814
rect -102483 -135858 -102439 -135814
rect -102383 -135858 -102339 -135814
rect -102283 -135858 -102239 -135814
rect -102183 -135858 -102139 -135814
rect -102083 -135858 -102039 -135814
rect -101983 -135858 -101939 -135814
rect -101883 -135858 -101839 -135814
rect -101783 -135858 -101739 -135814
rect -101683 -135858 -101639 -135814
rect -101583 -135858 -101539 -135814
rect -101483 -135858 -101439 -135814
rect -101383 -135858 -101339 -135814
rect -101283 -135858 -101239 -135814
rect -100783 -135858 -100739 -135814
rect -100683 -135858 -100639 -135814
rect -100583 -135858 -100539 -135814
rect -100483 -135858 -100439 -135814
rect -100383 -135858 -100339 -135814
rect -100283 -135858 -100239 -135814
rect -100183 -135858 -100139 -135814
rect -100083 -135858 -100039 -135814
rect -99983 -135858 -99939 -135814
rect -99883 -135858 -99839 -135814
rect -99783 -135858 -99739 -135814
rect -99683 -135858 -99639 -135814
rect -99583 -135858 -99539 -135814
rect -99483 -135858 -99439 -135814
rect -99383 -135858 -99339 -135814
rect -99283 -135858 -99239 -135814
rect -98783 -135858 -98739 -135814
rect -98683 -135858 -98639 -135814
rect -98583 -135858 -98539 -135814
rect -98483 -135858 -98439 -135814
rect -98383 -135858 -98339 -135814
rect -98283 -135858 -98239 -135814
rect -98183 -135858 -98139 -135814
rect -98083 -135858 -98039 -135814
rect -97983 -135858 -97939 -135814
rect -97883 -135858 -97839 -135814
rect -97783 -135858 -97739 -135814
rect -97683 -135858 -97639 -135814
rect -97583 -135858 -97539 -135814
rect -97483 -135858 -97439 -135814
rect -97383 -135858 -97339 -135814
rect -97283 -135858 -97239 -135814
rect -104783 -135958 -104739 -135914
rect -104683 -135958 -104639 -135914
rect -104583 -135958 -104539 -135914
rect -104483 -135958 -104439 -135914
rect -104383 -135958 -104339 -135914
rect -104283 -135958 -104239 -135914
rect -104183 -135958 -104139 -135914
rect -104083 -135958 -104039 -135914
rect -103983 -135958 -103939 -135914
rect -103883 -135958 -103839 -135914
rect -103783 -135958 -103739 -135914
rect -103683 -135958 -103639 -135914
rect -103583 -135958 -103539 -135914
rect -103483 -135958 -103439 -135914
rect -103383 -135958 -103339 -135914
rect -103283 -135958 -103239 -135914
rect -102783 -135958 -102739 -135914
rect -102683 -135958 -102639 -135914
rect -102583 -135958 -102539 -135914
rect -102483 -135958 -102439 -135914
rect -102383 -135958 -102339 -135914
rect -102283 -135958 -102239 -135914
rect -102183 -135958 -102139 -135914
rect -102083 -135958 -102039 -135914
rect -101983 -135958 -101939 -135914
rect -101883 -135958 -101839 -135914
rect -101783 -135958 -101739 -135914
rect -101683 -135958 -101639 -135914
rect -101583 -135958 -101539 -135914
rect -101483 -135958 -101439 -135914
rect -101383 -135958 -101339 -135914
rect -101283 -135958 -101239 -135914
rect -100783 -135958 -100739 -135914
rect -100683 -135958 -100639 -135914
rect -100583 -135958 -100539 -135914
rect -100483 -135958 -100439 -135914
rect -100383 -135958 -100339 -135914
rect -100283 -135958 -100239 -135914
rect -100183 -135958 -100139 -135914
rect -100083 -135958 -100039 -135914
rect -99983 -135958 -99939 -135914
rect -99883 -135958 -99839 -135914
rect -99783 -135958 -99739 -135914
rect -99683 -135958 -99639 -135914
rect -99583 -135958 -99539 -135914
rect -99483 -135958 -99439 -135914
rect -99383 -135958 -99339 -135914
rect -99283 -135958 -99239 -135914
rect -98783 -135958 -98739 -135914
rect -98683 -135958 -98639 -135914
rect -98583 -135958 -98539 -135914
rect -98483 -135958 -98439 -135914
rect -98383 -135958 -98339 -135914
rect -98283 -135958 -98239 -135914
rect -98183 -135958 -98139 -135914
rect -98083 -135958 -98039 -135914
rect -97983 -135958 -97939 -135914
rect -97883 -135958 -97839 -135914
rect -97783 -135958 -97739 -135914
rect -97683 -135958 -97639 -135914
rect -97583 -135958 -97539 -135914
rect -97483 -135958 -97439 -135914
rect -97383 -135958 -97339 -135914
rect -97283 -135958 -97239 -135914
rect -104783 -136058 -104739 -136014
rect -104683 -136058 -104639 -136014
rect -104583 -136058 -104539 -136014
rect -104483 -136058 -104439 -136014
rect -104383 -136058 -104339 -136014
rect -104283 -136058 -104239 -136014
rect -104183 -136058 -104139 -136014
rect -104083 -136058 -104039 -136014
rect -103983 -136058 -103939 -136014
rect -103883 -136058 -103839 -136014
rect -103783 -136058 -103739 -136014
rect -103683 -136058 -103639 -136014
rect -103583 -136058 -103539 -136014
rect -103483 -136058 -103439 -136014
rect -103383 -136058 -103339 -136014
rect -103283 -136058 -103239 -136014
rect -102783 -136058 -102739 -136014
rect -102683 -136058 -102639 -136014
rect -102583 -136058 -102539 -136014
rect -102483 -136058 -102439 -136014
rect -102383 -136058 -102339 -136014
rect -102283 -136058 -102239 -136014
rect -102183 -136058 -102139 -136014
rect -102083 -136058 -102039 -136014
rect -101983 -136058 -101939 -136014
rect -101883 -136058 -101839 -136014
rect -101783 -136058 -101739 -136014
rect -101683 -136058 -101639 -136014
rect -101583 -136058 -101539 -136014
rect -101483 -136058 -101439 -136014
rect -101383 -136058 -101339 -136014
rect -101283 -136058 -101239 -136014
rect -100783 -136058 -100739 -136014
rect -100683 -136058 -100639 -136014
rect -100583 -136058 -100539 -136014
rect -100483 -136058 -100439 -136014
rect -100383 -136058 -100339 -136014
rect -100283 -136058 -100239 -136014
rect -100183 -136058 -100139 -136014
rect -100083 -136058 -100039 -136014
rect -99983 -136058 -99939 -136014
rect -99883 -136058 -99839 -136014
rect -99783 -136058 -99739 -136014
rect -99683 -136058 -99639 -136014
rect -99583 -136058 -99539 -136014
rect -99483 -136058 -99439 -136014
rect -99383 -136058 -99339 -136014
rect -99283 -136058 -99239 -136014
rect -98783 -136058 -98739 -136014
rect -98683 -136058 -98639 -136014
rect -98583 -136058 -98539 -136014
rect -98483 -136058 -98439 -136014
rect -98383 -136058 -98339 -136014
rect -98283 -136058 -98239 -136014
rect -98183 -136058 -98139 -136014
rect -98083 -136058 -98039 -136014
rect -97983 -136058 -97939 -136014
rect -97883 -136058 -97839 -136014
rect -97783 -136058 -97739 -136014
rect -97683 -136058 -97639 -136014
rect -97583 -136058 -97539 -136014
rect -97483 -136058 -97439 -136014
rect -97383 -136058 -97339 -136014
rect -97283 -136058 -97239 -136014
rect -104783 -136158 -104739 -136114
rect -104683 -136158 -104639 -136114
rect -104583 -136158 -104539 -136114
rect -104483 -136158 -104439 -136114
rect -104383 -136158 -104339 -136114
rect -104283 -136158 -104239 -136114
rect -104183 -136158 -104139 -136114
rect -104083 -136158 -104039 -136114
rect -103983 -136158 -103939 -136114
rect -103883 -136158 -103839 -136114
rect -103783 -136158 -103739 -136114
rect -103683 -136158 -103639 -136114
rect -103583 -136158 -103539 -136114
rect -103483 -136158 -103439 -136114
rect -103383 -136158 -103339 -136114
rect -103283 -136158 -103239 -136114
rect -102783 -136158 -102739 -136114
rect -102683 -136158 -102639 -136114
rect -102583 -136158 -102539 -136114
rect -102483 -136158 -102439 -136114
rect -102383 -136158 -102339 -136114
rect -102283 -136158 -102239 -136114
rect -102183 -136158 -102139 -136114
rect -102083 -136158 -102039 -136114
rect -101983 -136158 -101939 -136114
rect -101883 -136158 -101839 -136114
rect -101783 -136158 -101739 -136114
rect -101683 -136158 -101639 -136114
rect -101583 -136158 -101539 -136114
rect -101483 -136158 -101439 -136114
rect -101383 -136158 -101339 -136114
rect -101283 -136158 -101239 -136114
rect -100783 -136158 -100739 -136114
rect -100683 -136158 -100639 -136114
rect -100583 -136158 -100539 -136114
rect -100483 -136158 -100439 -136114
rect -100383 -136158 -100339 -136114
rect -100283 -136158 -100239 -136114
rect -100183 -136158 -100139 -136114
rect -100083 -136158 -100039 -136114
rect -99983 -136158 -99939 -136114
rect -99883 -136158 -99839 -136114
rect -99783 -136158 -99739 -136114
rect -99683 -136158 -99639 -136114
rect -99583 -136158 -99539 -136114
rect -99483 -136158 -99439 -136114
rect -99383 -136158 -99339 -136114
rect -99283 -136158 -99239 -136114
rect -98783 -136158 -98739 -136114
rect -98683 -136158 -98639 -136114
rect -98583 -136158 -98539 -136114
rect -98483 -136158 -98439 -136114
rect -98383 -136158 -98339 -136114
rect -98283 -136158 -98239 -136114
rect -98183 -136158 -98139 -136114
rect -98083 -136158 -98039 -136114
rect -97983 -136158 -97939 -136114
rect -97883 -136158 -97839 -136114
rect -97783 -136158 -97739 -136114
rect -97683 -136158 -97639 -136114
rect -97583 -136158 -97539 -136114
rect -97483 -136158 -97439 -136114
rect -97383 -136158 -97339 -136114
rect -97283 -136158 -97239 -136114
rect -104783 -136258 -104739 -136214
rect -104683 -136258 -104639 -136214
rect -104583 -136258 -104539 -136214
rect -104483 -136258 -104439 -136214
rect -104383 -136258 -104339 -136214
rect -104283 -136258 -104239 -136214
rect -104183 -136258 -104139 -136214
rect -104083 -136258 -104039 -136214
rect -103983 -136258 -103939 -136214
rect -103883 -136258 -103839 -136214
rect -103783 -136258 -103739 -136214
rect -103683 -136258 -103639 -136214
rect -103583 -136258 -103539 -136214
rect -103483 -136258 -103439 -136214
rect -103383 -136258 -103339 -136214
rect -103283 -136258 -103239 -136214
rect -102783 -136258 -102739 -136214
rect -102683 -136258 -102639 -136214
rect -102583 -136258 -102539 -136214
rect -102483 -136258 -102439 -136214
rect -102383 -136258 -102339 -136214
rect -102283 -136258 -102239 -136214
rect -102183 -136258 -102139 -136214
rect -102083 -136258 -102039 -136214
rect -101983 -136258 -101939 -136214
rect -101883 -136258 -101839 -136214
rect -101783 -136258 -101739 -136214
rect -101683 -136258 -101639 -136214
rect -101583 -136258 -101539 -136214
rect -101483 -136258 -101439 -136214
rect -101383 -136258 -101339 -136214
rect -101283 -136258 -101239 -136214
rect -100783 -136258 -100739 -136214
rect -100683 -136258 -100639 -136214
rect -100583 -136258 -100539 -136214
rect -100483 -136258 -100439 -136214
rect -100383 -136258 -100339 -136214
rect -100283 -136258 -100239 -136214
rect -100183 -136258 -100139 -136214
rect -100083 -136258 -100039 -136214
rect -99983 -136258 -99939 -136214
rect -99883 -136258 -99839 -136214
rect -99783 -136258 -99739 -136214
rect -99683 -136258 -99639 -136214
rect -99583 -136258 -99539 -136214
rect -99483 -136258 -99439 -136214
rect -99383 -136258 -99339 -136214
rect -99283 -136258 -99239 -136214
rect -98783 -136258 -98739 -136214
rect -98683 -136258 -98639 -136214
rect -98583 -136258 -98539 -136214
rect -98483 -136258 -98439 -136214
rect -98383 -136258 -98339 -136214
rect -98283 -136258 -98239 -136214
rect -98183 -136258 -98139 -136214
rect -98083 -136258 -98039 -136214
rect -97983 -136258 -97939 -136214
rect -97883 -136258 -97839 -136214
rect -97783 -136258 -97739 -136214
rect -97683 -136258 -97639 -136214
rect -97583 -136258 -97539 -136214
rect -97483 -136258 -97439 -136214
rect -97383 -136258 -97339 -136214
rect -97283 -136258 -97239 -136214
rect -104783 -136358 -104739 -136314
rect -104683 -136358 -104639 -136314
rect -104583 -136358 -104539 -136314
rect -104483 -136358 -104439 -136314
rect -104383 -136358 -104339 -136314
rect -104283 -136358 -104239 -136314
rect -104183 -136358 -104139 -136314
rect -104083 -136358 -104039 -136314
rect -103983 -136358 -103939 -136314
rect -103883 -136358 -103839 -136314
rect -103783 -136358 -103739 -136314
rect -103683 -136358 -103639 -136314
rect -103583 -136358 -103539 -136314
rect -103483 -136358 -103439 -136314
rect -103383 -136358 -103339 -136314
rect -103283 -136358 -103239 -136314
rect -102783 -136358 -102739 -136314
rect -102683 -136358 -102639 -136314
rect -102583 -136358 -102539 -136314
rect -102483 -136358 -102439 -136314
rect -102383 -136358 -102339 -136314
rect -102283 -136358 -102239 -136314
rect -102183 -136358 -102139 -136314
rect -102083 -136358 -102039 -136314
rect -101983 -136358 -101939 -136314
rect -101883 -136358 -101839 -136314
rect -101783 -136358 -101739 -136314
rect -101683 -136358 -101639 -136314
rect -101583 -136358 -101539 -136314
rect -101483 -136358 -101439 -136314
rect -101383 -136358 -101339 -136314
rect -101283 -136358 -101239 -136314
rect -100783 -136358 -100739 -136314
rect -100683 -136358 -100639 -136314
rect -100583 -136358 -100539 -136314
rect -100483 -136358 -100439 -136314
rect -100383 -136358 -100339 -136314
rect -100283 -136358 -100239 -136314
rect -100183 -136358 -100139 -136314
rect -100083 -136358 -100039 -136314
rect -99983 -136358 -99939 -136314
rect -99883 -136358 -99839 -136314
rect -99783 -136358 -99739 -136314
rect -99683 -136358 -99639 -136314
rect -99583 -136358 -99539 -136314
rect -99483 -136358 -99439 -136314
rect -99383 -136358 -99339 -136314
rect -99283 -136358 -99239 -136314
rect -98783 -136358 -98739 -136314
rect -98683 -136358 -98639 -136314
rect -98583 -136358 -98539 -136314
rect -98483 -136358 -98439 -136314
rect -98383 -136358 -98339 -136314
rect -98283 -136358 -98239 -136314
rect -98183 -136358 -98139 -136314
rect -98083 -136358 -98039 -136314
rect -97983 -136358 -97939 -136314
rect -97883 -136358 -97839 -136314
rect -97783 -136358 -97739 -136314
rect -97683 -136358 -97639 -136314
rect -97583 -136358 -97539 -136314
rect -97483 -136358 -97439 -136314
rect -97383 -136358 -97339 -136314
rect -97283 -136358 -97239 -136314
rect -104783 -136458 -104739 -136414
rect -104683 -136458 -104639 -136414
rect -104583 -136458 -104539 -136414
rect -104483 -136458 -104439 -136414
rect -104383 -136458 -104339 -136414
rect -104283 -136458 -104239 -136414
rect -104183 -136458 -104139 -136414
rect -104083 -136458 -104039 -136414
rect -103983 -136458 -103939 -136414
rect -103883 -136458 -103839 -136414
rect -103783 -136458 -103739 -136414
rect -103683 -136458 -103639 -136414
rect -103583 -136458 -103539 -136414
rect -103483 -136458 -103439 -136414
rect -103383 -136458 -103339 -136414
rect -103283 -136458 -103239 -136414
rect -102783 -136458 -102739 -136414
rect -102683 -136458 -102639 -136414
rect -102583 -136458 -102539 -136414
rect -102483 -136458 -102439 -136414
rect -102383 -136458 -102339 -136414
rect -102283 -136458 -102239 -136414
rect -102183 -136458 -102139 -136414
rect -102083 -136458 -102039 -136414
rect -101983 -136458 -101939 -136414
rect -101883 -136458 -101839 -136414
rect -101783 -136458 -101739 -136414
rect -101683 -136458 -101639 -136414
rect -101583 -136458 -101539 -136414
rect -101483 -136458 -101439 -136414
rect -101383 -136458 -101339 -136414
rect -101283 -136458 -101239 -136414
rect -100783 -136458 -100739 -136414
rect -100683 -136458 -100639 -136414
rect -100583 -136458 -100539 -136414
rect -100483 -136458 -100439 -136414
rect -100383 -136458 -100339 -136414
rect -100283 -136458 -100239 -136414
rect -100183 -136458 -100139 -136414
rect -100083 -136458 -100039 -136414
rect -99983 -136458 -99939 -136414
rect -99883 -136458 -99839 -136414
rect -99783 -136458 -99739 -136414
rect -99683 -136458 -99639 -136414
rect -99583 -136458 -99539 -136414
rect -99483 -136458 -99439 -136414
rect -99383 -136458 -99339 -136414
rect -99283 -136458 -99239 -136414
rect -98783 -136458 -98739 -136414
rect -98683 -136458 -98639 -136414
rect -98583 -136458 -98539 -136414
rect -98483 -136458 -98439 -136414
rect -98383 -136458 -98339 -136414
rect -98283 -136458 -98239 -136414
rect -98183 -136458 -98139 -136414
rect -98083 -136458 -98039 -136414
rect -97983 -136458 -97939 -136414
rect -97883 -136458 -97839 -136414
rect -97783 -136458 -97739 -136414
rect -97683 -136458 -97639 -136414
rect -97583 -136458 -97539 -136414
rect -97483 -136458 -97439 -136414
rect -97383 -136458 -97339 -136414
rect -97283 -136458 -97239 -136414
rect -104783 -136558 -104739 -136514
rect -104683 -136558 -104639 -136514
rect -104583 -136558 -104539 -136514
rect -104483 -136558 -104439 -136514
rect -104383 -136558 -104339 -136514
rect -104283 -136558 -104239 -136514
rect -104183 -136558 -104139 -136514
rect -104083 -136558 -104039 -136514
rect -103983 -136558 -103939 -136514
rect -103883 -136558 -103839 -136514
rect -103783 -136558 -103739 -136514
rect -103683 -136558 -103639 -136514
rect -103583 -136558 -103539 -136514
rect -103483 -136558 -103439 -136514
rect -103383 -136558 -103339 -136514
rect -103283 -136558 -103239 -136514
rect -102783 -136558 -102739 -136514
rect -102683 -136558 -102639 -136514
rect -102583 -136558 -102539 -136514
rect -102483 -136558 -102439 -136514
rect -102383 -136558 -102339 -136514
rect -102283 -136558 -102239 -136514
rect -102183 -136558 -102139 -136514
rect -102083 -136558 -102039 -136514
rect -101983 -136558 -101939 -136514
rect -101883 -136558 -101839 -136514
rect -101783 -136558 -101739 -136514
rect -101683 -136558 -101639 -136514
rect -101583 -136558 -101539 -136514
rect -101483 -136558 -101439 -136514
rect -101383 -136558 -101339 -136514
rect -101283 -136558 -101239 -136514
rect -100783 -136558 -100739 -136514
rect -100683 -136558 -100639 -136514
rect -100583 -136558 -100539 -136514
rect -100483 -136558 -100439 -136514
rect -100383 -136558 -100339 -136514
rect -100283 -136558 -100239 -136514
rect -100183 -136558 -100139 -136514
rect -100083 -136558 -100039 -136514
rect -99983 -136558 -99939 -136514
rect -99883 -136558 -99839 -136514
rect -99783 -136558 -99739 -136514
rect -99683 -136558 -99639 -136514
rect -99583 -136558 -99539 -136514
rect -99483 -136558 -99439 -136514
rect -99383 -136558 -99339 -136514
rect -99283 -136558 -99239 -136514
rect -98783 -136558 -98739 -136514
rect -98683 -136558 -98639 -136514
rect -98583 -136558 -98539 -136514
rect -98483 -136558 -98439 -136514
rect -98383 -136558 -98339 -136514
rect -98283 -136558 -98239 -136514
rect -98183 -136558 -98139 -136514
rect -98083 -136558 -98039 -136514
rect -97983 -136558 -97939 -136514
rect -97883 -136558 -97839 -136514
rect -97783 -136558 -97739 -136514
rect -97683 -136558 -97639 -136514
rect -97583 -136558 -97539 -136514
rect -97483 -136558 -97439 -136514
rect -97383 -136558 -97339 -136514
rect -97283 -136558 -97239 -136514
rect -104783 -136658 -104739 -136614
rect -104683 -136658 -104639 -136614
rect -104583 -136658 -104539 -136614
rect -104483 -136658 -104439 -136614
rect -104383 -136658 -104339 -136614
rect -104283 -136658 -104239 -136614
rect -104183 -136658 -104139 -136614
rect -104083 -136658 -104039 -136614
rect -103983 -136658 -103939 -136614
rect -103883 -136658 -103839 -136614
rect -103783 -136658 -103739 -136614
rect -103683 -136658 -103639 -136614
rect -103583 -136658 -103539 -136614
rect -103483 -136658 -103439 -136614
rect -103383 -136658 -103339 -136614
rect -103283 -136658 -103239 -136614
rect -102783 -136658 -102739 -136614
rect -102683 -136658 -102639 -136614
rect -102583 -136658 -102539 -136614
rect -102483 -136658 -102439 -136614
rect -102383 -136658 -102339 -136614
rect -102283 -136658 -102239 -136614
rect -102183 -136658 -102139 -136614
rect -102083 -136658 -102039 -136614
rect -101983 -136658 -101939 -136614
rect -101883 -136658 -101839 -136614
rect -101783 -136658 -101739 -136614
rect -101683 -136658 -101639 -136614
rect -101583 -136658 -101539 -136614
rect -101483 -136658 -101439 -136614
rect -101383 -136658 -101339 -136614
rect -101283 -136658 -101239 -136614
rect -100783 -136658 -100739 -136614
rect -100683 -136658 -100639 -136614
rect -100583 -136658 -100539 -136614
rect -100483 -136658 -100439 -136614
rect -100383 -136658 -100339 -136614
rect -100283 -136658 -100239 -136614
rect -100183 -136658 -100139 -136614
rect -100083 -136658 -100039 -136614
rect -99983 -136658 -99939 -136614
rect -99883 -136658 -99839 -136614
rect -99783 -136658 -99739 -136614
rect -99683 -136658 -99639 -136614
rect -99583 -136658 -99539 -136614
rect -99483 -136658 -99439 -136614
rect -99383 -136658 -99339 -136614
rect -99283 -136658 -99239 -136614
rect -98783 -136658 -98739 -136614
rect -98683 -136658 -98639 -136614
rect -98583 -136658 -98539 -136614
rect -98483 -136658 -98439 -136614
rect -98383 -136658 -98339 -136614
rect -98283 -136658 -98239 -136614
rect -98183 -136658 -98139 -136614
rect -98083 -136658 -98039 -136614
rect -97983 -136658 -97939 -136614
rect -97883 -136658 -97839 -136614
rect -97783 -136658 -97739 -136614
rect -97683 -136658 -97639 -136614
rect -97583 -136658 -97539 -136614
rect -97483 -136658 -97439 -136614
rect -97383 -136658 -97339 -136614
rect -97283 -136658 -97239 -136614
rect -104783 -136758 -104739 -136714
rect -104683 -136758 -104639 -136714
rect -104583 -136758 -104539 -136714
rect -104483 -136758 -104439 -136714
rect -104383 -136758 -104339 -136714
rect -104283 -136758 -104239 -136714
rect -104183 -136758 -104139 -136714
rect -104083 -136758 -104039 -136714
rect -103983 -136758 -103939 -136714
rect -103883 -136758 -103839 -136714
rect -103783 -136758 -103739 -136714
rect -103683 -136758 -103639 -136714
rect -103583 -136758 -103539 -136714
rect -103483 -136758 -103439 -136714
rect -103383 -136758 -103339 -136714
rect -103283 -136758 -103239 -136714
rect -102783 -136758 -102739 -136714
rect -102683 -136758 -102639 -136714
rect -102583 -136758 -102539 -136714
rect -102483 -136758 -102439 -136714
rect -102383 -136758 -102339 -136714
rect -102283 -136758 -102239 -136714
rect -102183 -136758 -102139 -136714
rect -102083 -136758 -102039 -136714
rect -101983 -136758 -101939 -136714
rect -101883 -136758 -101839 -136714
rect -101783 -136758 -101739 -136714
rect -101683 -136758 -101639 -136714
rect -101583 -136758 -101539 -136714
rect -101483 -136758 -101439 -136714
rect -101383 -136758 -101339 -136714
rect -101283 -136758 -101239 -136714
rect -100783 -136758 -100739 -136714
rect -100683 -136758 -100639 -136714
rect -100583 -136758 -100539 -136714
rect -100483 -136758 -100439 -136714
rect -100383 -136758 -100339 -136714
rect -100283 -136758 -100239 -136714
rect -100183 -136758 -100139 -136714
rect -100083 -136758 -100039 -136714
rect -99983 -136758 -99939 -136714
rect -99883 -136758 -99839 -136714
rect -99783 -136758 -99739 -136714
rect -99683 -136758 -99639 -136714
rect -99583 -136758 -99539 -136714
rect -99483 -136758 -99439 -136714
rect -99383 -136758 -99339 -136714
rect -99283 -136758 -99239 -136714
rect -98783 -136758 -98739 -136714
rect -98683 -136758 -98639 -136714
rect -98583 -136758 -98539 -136714
rect -98483 -136758 -98439 -136714
rect -98383 -136758 -98339 -136714
rect -98283 -136758 -98239 -136714
rect -98183 -136758 -98139 -136714
rect -98083 -136758 -98039 -136714
rect -97983 -136758 -97939 -136714
rect -97883 -136758 -97839 -136714
rect -97783 -136758 -97739 -136714
rect -97683 -136758 -97639 -136714
rect -97583 -136758 -97539 -136714
rect -97483 -136758 -97439 -136714
rect -97383 -136758 -97339 -136714
rect -97283 -136758 -97239 -136714
rect -104783 -136858 -104739 -136814
rect -104683 -136858 -104639 -136814
rect -104583 -136858 -104539 -136814
rect -104483 -136858 -104439 -136814
rect -104383 -136858 -104339 -136814
rect -104283 -136858 -104239 -136814
rect -104183 -136858 -104139 -136814
rect -104083 -136858 -104039 -136814
rect -103983 -136858 -103939 -136814
rect -103883 -136858 -103839 -136814
rect -103783 -136858 -103739 -136814
rect -103683 -136858 -103639 -136814
rect -103583 -136858 -103539 -136814
rect -103483 -136858 -103439 -136814
rect -103383 -136858 -103339 -136814
rect -103283 -136858 -103239 -136814
rect -102783 -136858 -102739 -136814
rect -102683 -136858 -102639 -136814
rect -102583 -136858 -102539 -136814
rect -102483 -136858 -102439 -136814
rect -102383 -136858 -102339 -136814
rect -102283 -136858 -102239 -136814
rect -102183 -136858 -102139 -136814
rect -102083 -136858 -102039 -136814
rect -101983 -136858 -101939 -136814
rect -101883 -136858 -101839 -136814
rect -101783 -136858 -101739 -136814
rect -101683 -136858 -101639 -136814
rect -101583 -136858 -101539 -136814
rect -101483 -136858 -101439 -136814
rect -101383 -136858 -101339 -136814
rect -101283 -136858 -101239 -136814
rect -100783 -136858 -100739 -136814
rect -100683 -136858 -100639 -136814
rect -100583 -136858 -100539 -136814
rect -100483 -136858 -100439 -136814
rect -100383 -136858 -100339 -136814
rect -100283 -136858 -100239 -136814
rect -100183 -136858 -100139 -136814
rect -100083 -136858 -100039 -136814
rect -99983 -136858 -99939 -136814
rect -99883 -136858 -99839 -136814
rect -99783 -136858 -99739 -136814
rect -99683 -136858 -99639 -136814
rect -99583 -136858 -99539 -136814
rect -99483 -136858 -99439 -136814
rect -99383 -136858 -99339 -136814
rect -99283 -136858 -99239 -136814
rect -98783 -136858 -98739 -136814
rect -98683 -136858 -98639 -136814
rect -98583 -136858 -98539 -136814
rect -98483 -136858 -98439 -136814
rect -98383 -136858 -98339 -136814
rect -98283 -136858 -98239 -136814
rect -98183 -136858 -98139 -136814
rect -98083 -136858 -98039 -136814
rect -97983 -136858 -97939 -136814
rect -97883 -136858 -97839 -136814
rect -97783 -136858 -97739 -136814
rect -97683 -136858 -97639 -136814
rect -97583 -136858 -97539 -136814
rect -97483 -136858 -97439 -136814
rect -97383 -136858 -97339 -136814
rect -97283 -136858 -97239 -136814
rect 81632 -138010 81676 -137966
rect 81732 -138010 81776 -137966
rect 81832 -138010 81876 -137966
rect 81932 -138010 81976 -137966
rect 82032 -138010 82076 -137966
rect 82132 -138010 82176 -137966
rect 82232 -138010 82276 -137966
rect 82332 -138010 82376 -137966
rect 82432 -138010 82476 -137966
rect 82532 -138010 82576 -137966
rect 82632 -138010 82676 -137966
rect 82732 -138010 82776 -137966
rect 82832 -138010 82876 -137966
rect 82932 -138010 82976 -137966
rect 83032 -138010 83076 -137966
rect 83132 -138010 83176 -137966
rect 83632 -138010 83676 -137966
rect 83732 -138010 83776 -137966
rect 83832 -138010 83876 -137966
rect 83932 -138010 83976 -137966
rect 84032 -138010 84076 -137966
rect 84132 -138010 84176 -137966
rect 84232 -138010 84276 -137966
rect 84332 -138010 84376 -137966
rect 84432 -138010 84476 -137966
rect 84532 -138010 84576 -137966
rect 84632 -138010 84676 -137966
rect 84732 -138010 84776 -137966
rect 84832 -138010 84876 -137966
rect 84932 -138010 84976 -137966
rect 85032 -138010 85076 -137966
rect 85132 -138010 85176 -137966
rect 85632 -138010 85676 -137966
rect 85732 -138010 85776 -137966
rect 85832 -138010 85876 -137966
rect 85932 -138010 85976 -137966
rect 86032 -138010 86076 -137966
rect 86132 -138010 86176 -137966
rect 86232 -138010 86276 -137966
rect 86332 -138010 86376 -137966
rect 86432 -138010 86476 -137966
rect 86532 -138010 86576 -137966
rect 86632 -138010 86676 -137966
rect 86732 -138010 86776 -137966
rect 86832 -138010 86876 -137966
rect 86932 -138010 86976 -137966
rect 87032 -138010 87076 -137966
rect 87132 -138010 87176 -137966
rect 87632 -138010 87676 -137966
rect 87732 -138010 87776 -137966
rect 87832 -138010 87876 -137966
rect 87932 -138010 87976 -137966
rect 88032 -138010 88076 -137966
rect 88132 -138010 88176 -137966
rect 88232 -138010 88276 -137966
rect 88332 -138010 88376 -137966
rect 88432 -138010 88476 -137966
rect 88532 -138010 88576 -137966
rect 88632 -138010 88676 -137966
rect 88732 -138010 88776 -137966
rect 88832 -138010 88876 -137966
rect 88932 -138010 88976 -137966
rect 89032 -138010 89076 -137966
rect 89132 -138010 89176 -137966
rect 81632 -138110 81676 -138066
rect 81732 -138110 81776 -138066
rect 81832 -138110 81876 -138066
rect 81932 -138110 81976 -138066
rect 82032 -138110 82076 -138066
rect 82132 -138110 82176 -138066
rect 82232 -138110 82276 -138066
rect 82332 -138110 82376 -138066
rect 82432 -138110 82476 -138066
rect 82532 -138110 82576 -138066
rect 82632 -138110 82676 -138066
rect 82732 -138110 82776 -138066
rect 82832 -138110 82876 -138066
rect 82932 -138110 82976 -138066
rect 83032 -138110 83076 -138066
rect 83132 -138110 83176 -138066
rect 83632 -138110 83676 -138066
rect 83732 -138110 83776 -138066
rect 83832 -138110 83876 -138066
rect 83932 -138110 83976 -138066
rect 84032 -138110 84076 -138066
rect 84132 -138110 84176 -138066
rect 84232 -138110 84276 -138066
rect 84332 -138110 84376 -138066
rect 84432 -138110 84476 -138066
rect 84532 -138110 84576 -138066
rect 84632 -138110 84676 -138066
rect 84732 -138110 84776 -138066
rect 84832 -138110 84876 -138066
rect 84932 -138110 84976 -138066
rect 85032 -138110 85076 -138066
rect 85132 -138110 85176 -138066
rect 85632 -138110 85676 -138066
rect 85732 -138110 85776 -138066
rect 85832 -138110 85876 -138066
rect 85932 -138110 85976 -138066
rect 86032 -138110 86076 -138066
rect 86132 -138110 86176 -138066
rect 86232 -138110 86276 -138066
rect 86332 -138110 86376 -138066
rect 86432 -138110 86476 -138066
rect 86532 -138110 86576 -138066
rect 86632 -138110 86676 -138066
rect 86732 -138110 86776 -138066
rect 86832 -138110 86876 -138066
rect 86932 -138110 86976 -138066
rect 87032 -138110 87076 -138066
rect 87132 -138110 87176 -138066
rect 87632 -138110 87676 -138066
rect 87732 -138110 87776 -138066
rect 87832 -138110 87876 -138066
rect 87932 -138110 87976 -138066
rect 88032 -138110 88076 -138066
rect 88132 -138110 88176 -138066
rect 88232 -138110 88276 -138066
rect 88332 -138110 88376 -138066
rect 88432 -138110 88476 -138066
rect 88532 -138110 88576 -138066
rect 88632 -138110 88676 -138066
rect 88732 -138110 88776 -138066
rect 88832 -138110 88876 -138066
rect 88932 -138110 88976 -138066
rect 89032 -138110 89076 -138066
rect 89132 -138110 89176 -138066
rect 81632 -138210 81676 -138166
rect 81732 -138210 81776 -138166
rect 81832 -138210 81876 -138166
rect 81932 -138210 81976 -138166
rect 82032 -138210 82076 -138166
rect 82132 -138210 82176 -138166
rect 82232 -138210 82276 -138166
rect 82332 -138210 82376 -138166
rect 82432 -138210 82476 -138166
rect 82532 -138210 82576 -138166
rect 82632 -138210 82676 -138166
rect 82732 -138210 82776 -138166
rect 82832 -138210 82876 -138166
rect 82932 -138210 82976 -138166
rect 83032 -138210 83076 -138166
rect 83132 -138210 83176 -138166
rect 83632 -138210 83676 -138166
rect 83732 -138210 83776 -138166
rect 83832 -138210 83876 -138166
rect 83932 -138210 83976 -138166
rect 84032 -138210 84076 -138166
rect 84132 -138210 84176 -138166
rect 84232 -138210 84276 -138166
rect 84332 -138210 84376 -138166
rect 84432 -138210 84476 -138166
rect 84532 -138210 84576 -138166
rect 84632 -138210 84676 -138166
rect 84732 -138210 84776 -138166
rect 84832 -138210 84876 -138166
rect 84932 -138210 84976 -138166
rect 85032 -138210 85076 -138166
rect 85132 -138210 85176 -138166
rect 85632 -138210 85676 -138166
rect 85732 -138210 85776 -138166
rect 85832 -138210 85876 -138166
rect 85932 -138210 85976 -138166
rect 86032 -138210 86076 -138166
rect 86132 -138210 86176 -138166
rect 86232 -138210 86276 -138166
rect 86332 -138210 86376 -138166
rect 86432 -138210 86476 -138166
rect 86532 -138210 86576 -138166
rect 86632 -138210 86676 -138166
rect 86732 -138210 86776 -138166
rect 86832 -138210 86876 -138166
rect 86932 -138210 86976 -138166
rect 87032 -138210 87076 -138166
rect 87132 -138210 87176 -138166
rect 87632 -138210 87676 -138166
rect 87732 -138210 87776 -138166
rect 87832 -138210 87876 -138166
rect 87932 -138210 87976 -138166
rect 88032 -138210 88076 -138166
rect 88132 -138210 88176 -138166
rect 88232 -138210 88276 -138166
rect 88332 -138210 88376 -138166
rect 88432 -138210 88476 -138166
rect 88532 -138210 88576 -138166
rect 88632 -138210 88676 -138166
rect 88732 -138210 88776 -138166
rect 88832 -138210 88876 -138166
rect 88932 -138210 88976 -138166
rect 89032 -138210 89076 -138166
rect 89132 -138210 89176 -138166
rect -83265 -140275 -83221 -140231
rect -83165 -140275 -83121 -140231
rect -83065 -140275 -83021 -140231
rect -82965 -140275 -82921 -140231
rect -82865 -140275 -82821 -140231
rect -82765 -140275 -82721 -140231
rect -82665 -140275 -82621 -140231
rect -82565 -140275 -82521 -140231
rect -82465 -140275 -82421 -140231
rect -82365 -140275 -82321 -140231
rect -82265 -140275 -82221 -140231
rect -82165 -140275 -82121 -140231
rect -82065 -140275 -82021 -140231
rect -81965 -140275 -81921 -140231
rect -81865 -140275 -81821 -140231
rect -81765 -140275 -81721 -140231
rect -81265 -140275 -81221 -140231
rect -81165 -140275 -81121 -140231
rect -81065 -140275 -81021 -140231
rect -80965 -140275 -80921 -140231
rect -80865 -140275 -80821 -140231
rect -80765 -140275 -80721 -140231
rect -80665 -140275 -80621 -140231
rect -80565 -140275 -80521 -140231
rect -80465 -140275 -80421 -140231
rect -80365 -140275 -80321 -140231
rect -80265 -140275 -80221 -140231
rect -80165 -140275 -80121 -140231
rect -80065 -140275 -80021 -140231
rect -79965 -140275 -79921 -140231
rect -79865 -140275 -79821 -140231
rect -79765 -140275 -79721 -140231
rect -79265 -140275 -79221 -140231
rect -79165 -140275 -79121 -140231
rect -79065 -140275 -79021 -140231
rect -78965 -140275 -78921 -140231
rect -78865 -140275 -78821 -140231
rect -78765 -140275 -78721 -140231
rect -78665 -140275 -78621 -140231
rect -78565 -140275 -78521 -140231
rect -78465 -140275 -78421 -140231
rect -78365 -140275 -78321 -140231
rect -78265 -140275 -78221 -140231
rect -78165 -140275 -78121 -140231
rect -78065 -140275 -78021 -140231
rect -77965 -140275 -77921 -140231
rect -77865 -140275 -77821 -140231
rect -77765 -140275 -77721 -140231
rect -77265 -140275 -77221 -140231
rect -77165 -140275 -77121 -140231
rect -77065 -140275 -77021 -140231
rect -76965 -140275 -76921 -140231
rect -76865 -140275 -76821 -140231
rect -76765 -140275 -76721 -140231
rect -76665 -140275 -76621 -140231
rect -76565 -140275 -76521 -140231
rect -76465 -140275 -76421 -140231
rect -76365 -140275 -76321 -140231
rect -76265 -140275 -76221 -140231
rect -76165 -140275 -76121 -140231
rect -76065 -140275 -76021 -140231
rect -75965 -140275 -75921 -140231
rect -75865 -140275 -75821 -140231
rect -75765 -140275 -75721 -140231
rect -83265 -140375 -83221 -140331
rect -83165 -140375 -83121 -140331
rect -83065 -140375 -83021 -140331
rect -82965 -140375 -82921 -140331
rect -82865 -140375 -82821 -140331
rect -82765 -140375 -82721 -140331
rect -82665 -140375 -82621 -140331
rect -82565 -140375 -82521 -140331
rect -82465 -140375 -82421 -140331
rect -82365 -140375 -82321 -140331
rect -82265 -140375 -82221 -140331
rect -82165 -140375 -82121 -140331
rect -82065 -140375 -82021 -140331
rect -81965 -140375 -81921 -140331
rect -81865 -140375 -81821 -140331
rect -81765 -140375 -81721 -140331
rect -81265 -140375 -81221 -140331
rect -81165 -140375 -81121 -140331
rect -81065 -140375 -81021 -140331
rect -80965 -140375 -80921 -140331
rect -80865 -140375 -80821 -140331
rect -80765 -140375 -80721 -140331
rect -80665 -140375 -80621 -140331
rect -80565 -140375 -80521 -140331
rect -80465 -140375 -80421 -140331
rect -80365 -140375 -80321 -140331
rect -80265 -140375 -80221 -140331
rect -80165 -140375 -80121 -140331
rect -80065 -140375 -80021 -140331
rect -79965 -140375 -79921 -140331
rect -79865 -140375 -79821 -140331
rect -79765 -140375 -79721 -140331
rect -79265 -140375 -79221 -140331
rect -79165 -140375 -79121 -140331
rect -79065 -140375 -79021 -140331
rect -78965 -140375 -78921 -140331
rect -78865 -140375 -78821 -140331
rect -78765 -140375 -78721 -140331
rect -78665 -140375 -78621 -140331
rect -78565 -140375 -78521 -140331
rect -78465 -140375 -78421 -140331
rect -78365 -140375 -78321 -140331
rect -78265 -140375 -78221 -140331
rect -78165 -140375 -78121 -140331
rect -78065 -140375 -78021 -140331
rect -77965 -140375 -77921 -140331
rect -77865 -140375 -77821 -140331
rect -77765 -140375 -77721 -140331
rect -77265 -140375 -77221 -140331
rect -77165 -140375 -77121 -140331
rect -77065 -140375 -77021 -140331
rect -76965 -140375 -76921 -140331
rect -76865 -140375 -76821 -140331
rect -76765 -140375 -76721 -140331
rect -76665 -140375 -76621 -140331
rect -76565 -140375 -76521 -140331
rect -76465 -140375 -76421 -140331
rect -76365 -140375 -76321 -140331
rect -76265 -140375 -76221 -140331
rect -76165 -140375 -76121 -140331
rect -76065 -140375 -76021 -140331
rect -75965 -140375 -75921 -140331
rect -75865 -140375 -75821 -140331
rect -75765 -140375 -75721 -140331
rect -83265 -140475 -83221 -140431
rect -83165 -140475 -83121 -140431
rect -83065 -140475 -83021 -140431
rect -82965 -140475 -82921 -140431
rect -82865 -140475 -82821 -140431
rect -82765 -140475 -82721 -140431
rect -82665 -140475 -82621 -140431
rect -82565 -140475 -82521 -140431
rect -82465 -140475 -82421 -140431
rect -82365 -140475 -82321 -140431
rect -82265 -140475 -82221 -140431
rect -82165 -140475 -82121 -140431
rect -82065 -140475 -82021 -140431
rect -81965 -140475 -81921 -140431
rect -81865 -140475 -81821 -140431
rect -81765 -140475 -81721 -140431
rect -81265 -140475 -81221 -140431
rect -81165 -140475 -81121 -140431
rect -81065 -140475 -81021 -140431
rect -80965 -140475 -80921 -140431
rect -80865 -140475 -80821 -140431
rect -80765 -140475 -80721 -140431
rect -80665 -140475 -80621 -140431
rect -80565 -140475 -80521 -140431
rect -80465 -140475 -80421 -140431
rect -80365 -140475 -80321 -140431
rect -80265 -140475 -80221 -140431
rect -80165 -140475 -80121 -140431
rect -80065 -140475 -80021 -140431
rect -79965 -140475 -79921 -140431
rect -79865 -140475 -79821 -140431
rect -79765 -140475 -79721 -140431
rect -79265 -140475 -79221 -140431
rect -79165 -140475 -79121 -140431
rect -79065 -140475 -79021 -140431
rect -78965 -140475 -78921 -140431
rect -78865 -140475 -78821 -140431
rect -78765 -140475 -78721 -140431
rect -78665 -140475 -78621 -140431
rect -78565 -140475 -78521 -140431
rect -78465 -140475 -78421 -140431
rect -78365 -140475 -78321 -140431
rect -78265 -140475 -78221 -140431
rect -78165 -140475 -78121 -140431
rect -78065 -140475 -78021 -140431
rect -77965 -140475 -77921 -140431
rect -77865 -140475 -77821 -140431
rect -77765 -140475 -77721 -140431
rect -77265 -140475 -77221 -140431
rect -77165 -140475 -77121 -140431
rect -77065 -140475 -77021 -140431
rect -76965 -140475 -76921 -140431
rect -76865 -140475 -76821 -140431
rect -76765 -140475 -76721 -140431
rect -76665 -140475 -76621 -140431
rect -76565 -140475 -76521 -140431
rect -76465 -140475 -76421 -140431
rect -76365 -140475 -76321 -140431
rect -76265 -140475 -76221 -140431
rect -76165 -140475 -76121 -140431
rect -76065 -140475 -76021 -140431
rect -75965 -140475 -75921 -140431
rect -75865 -140475 -75821 -140431
rect -75765 -140475 -75721 -140431
rect -83265 -140575 -83221 -140531
rect -83165 -140575 -83121 -140531
rect -83065 -140575 -83021 -140531
rect -82965 -140575 -82921 -140531
rect -82865 -140575 -82821 -140531
rect -82765 -140575 -82721 -140531
rect -82665 -140575 -82621 -140531
rect -82565 -140575 -82521 -140531
rect -82465 -140575 -82421 -140531
rect -82365 -140575 -82321 -140531
rect -82265 -140575 -82221 -140531
rect -82165 -140575 -82121 -140531
rect -82065 -140575 -82021 -140531
rect -81965 -140575 -81921 -140531
rect -81865 -140575 -81821 -140531
rect -81765 -140575 -81721 -140531
rect -81265 -140575 -81221 -140531
rect -81165 -140575 -81121 -140531
rect -81065 -140575 -81021 -140531
rect -80965 -140575 -80921 -140531
rect -80865 -140575 -80821 -140531
rect -80765 -140575 -80721 -140531
rect -80665 -140575 -80621 -140531
rect -80565 -140575 -80521 -140531
rect -80465 -140575 -80421 -140531
rect -80365 -140575 -80321 -140531
rect -80265 -140575 -80221 -140531
rect -80165 -140575 -80121 -140531
rect -80065 -140575 -80021 -140531
rect -79965 -140575 -79921 -140531
rect -79865 -140575 -79821 -140531
rect -79765 -140575 -79721 -140531
rect -79265 -140575 -79221 -140531
rect -79165 -140575 -79121 -140531
rect -79065 -140575 -79021 -140531
rect -78965 -140575 -78921 -140531
rect -78865 -140575 -78821 -140531
rect -78765 -140575 -78721 -140531
rect -78665 -140575 -78621 -140531
rect -78565 -140575 -78521 -140531
rect -78465 -140575 -78421 -140531
rect -78365 -140575 -78321 -140531
rect -78265 -140575 -78221 -140531
rect -78165 -140575 -78121 -140531
rect -78065 -140575 -78021 -140531
rect -77965 -140575 -77921 -140531
rect -77865 -140575 -77821 -140531
rect -77765 -140575 -77721 -140531
rect -77265 -140575 -77221 -140531
rect -77165 -140575 -77121 -140531
rect -77065 -140575 -77021 -140531
rect -76965 -140575 -76921 -140531
rect -76865 -140575 -76821 -140531
rect -76765 -140575 -76721 -140531
rect -76665 -140575 -76621 -140531
rect -76565 -140575 -76521 -140531
rect -76465 -140575 -76421 -140531
rect -76365 -140575 -76321 -140531
rect -76265 -140575 -76221 -140531
rect -76165 -140575 -76121 -140531
rect -76065 -140575 -76021 -140531
rect -75965 -140575 -75921 -140531
rect -75865 -140575 -75821 -140531
rect -75765 -140575 -75721 -140531
rect -83265 -140675 -83221 -140631
rect -83165 -140675 -83121 -140631
rect -83065 -140675 -83021 -140631
rect -82965 -140675 -82921 -140631
rect -82865 -140675 -82821 -140631
rect -82765 -140675 -82721 -140631
rect -82665 -140675 -82621 -140631
rect -82565 -140675 -82521 -140631
rect -82465 -140675 -82421 -140631
rect -82365 -140675 -82321 -140631
rect -82265 -140675 -82221 -140631
rect -82165 -140675 -82121 -140631
rect -82065 -140675 -82021 -140631
rect -81965 -140675 -81921 -140631
rect -81865 -140675 -81821 -140631
rect -81765 -140675 -81721 -140631
rect -81265 -140675 -81221 -140631
rect -81165 -140675 -81121 -140631
rect -81065 -140675 -81021 -140631
rect -80965 -140675 -80921 -140631
rect -80865 -140675 -80821 -140631
rect -80765 -140675 -80721 -140631
rect -80665 -140675 -80621 -140631
rect -80565 -140675 -80521 -140631
rect -80465 -140675 -80421 -140631
rect -80365 -140675 -80321 -140631
rect -80265 -140675 -80221 -140631
rect -80165 -140675 -80121 -140631
rect -80065 -140675 -80021 -140631
rect -79965 -140675 -79921 -140631
rect -79865 -140675 -79821 -140631
rect -79765 -140675 -79721 -140631
rect -79265 -140675 -79221 -140631
rect -79165 -140675 -79121 -140631
rect -79065 -140675 -79021 -140631
rect -78965 -140675 -78921 -140631
rect -78865 -140675 -78821 -140631
rect -78765 -140675 -78721 -140631
rect -78665 -140675 -78621 -140631
rect -78565 -140675 -78521 -140631
rect -78465 -140675 -78421 -140631
rect -78365 -140675 -78321 -140631
rect -78265 -140675 -78221 -140631
rect -78165 -140675 -78121 -140631
rect -78065 -140675 -78021 -140631
rect -77965 -140675 -77921 -140631
rect -77865 -140675 -77821 -140631
rect -77765 -140675 -77721 -140631
rect -77265 -140675 -77221 -140631
rect -77165 -140675 -77121 -140631
rect -77065 -140675 -77021 -140631
rect -76965 -140675 -76921 -140631
rect -76865 -140675 -76821 -140631
rect -76765 -140675 -76721 -140631
rect -76665 -140675 -76621 -140631
rect -76565 -140675 -76521 -140631
rect -76465 -140675 -76421 -140631
rect -76365 -140675 -76321 -140631
rect -76265 -140675 -76221 -140631
rect -76165 -140675 -76121 -140631
rect -76065 -140675 -76021 -140631
rect -75965 -140675 -75921 -140631
rect -75865 -140675 -75821 -140631
rect -75765 -140675 -75721 -140631
rect -83265 -140775 -83221 -140731
rect -83165 -140775 -83121 -140731
rect -83065 -140775 -83021 -140731
rect -82965 -140775 -82921 -140731
rect -82865 -140775 -82821 -140731
rect -82765 -140775 -82721 -140731
rect -82665 -140775 -82621 -140731
rect -82565 -140775 -82521 -140731
rect -82465 -140775 -82421 -140731
rect -82365 -140775 -82321 -140731
rect -82265 -140775 -82221 -140731
rect -82165 -140775 -82121 -140731
rect -82065 -140775 -82021 -140731
rect -81965 -140775 -81921 -140731
rect -81865 -140775 -81821 -140731
rect -81765 -140775 -81721 -140731
rect -81265 -140775 -81221 -140731
rect -81165 -140775 -81121 -140731
rect -81065 -140775 -81021 -140731
rect -80965 -140775 -80921 -140731
rect -80865 -140775 -80821 -140731
rect -80765 -140775 -80721 -140731
rect -80665 -140775 -80621 -140731
rect -80565 -140775 -80521 -140731
rect -80465 -140775 -80421 -140731
rect -80365 -140775 -80321 -140731
rect -80265 -140775 -80221 -140731
rect -80165 -140775 -80121 -140731
rect -80065 -140775 -80021 -140731
rect -79965 -140775 -79921 -140731
rect -79865 -140775 -79821 -140731
rect -79765 -140775 -79721 -140731
rect -79265 -140775 -79221 -140731
rect -79165 -140775 -79121 -140731
rect -79065 -140775 -79021 -140731
rect -78965 -140775 -78921 -140731
rect -78865 -140775 -78821 -140731
rect -78765 -140775 -78721 -140731
rect -78665 -140775 -78621 -140731
rect -78565 -140775 -78521 -140731
rect -78465 -140775 -78421 -140731
rect -78365 -140775 -78321 -140731
rect -78265 -140775 -78221 -140731
rect -78165 -140775 -78121 -140731
rect -78065 -140775 -78021 -140731
rect -77965 -140775 -77921 -140731
rect -77865 -140775 -77821 -140731
rect -77765 -140775 -77721 -140731
rect -77265 -140775 -77221 -140731
rect -77165 -140775 -77121 -140731
rect -77065 -140775 -77021 -140731
rect -76965 -140775 -76921 -140731
rect -76865 -140775 -76821 -140731
rect -76765 -140775 -76721 -140731
rect -76665 -140775 -76621 -140731
rect -76565 -140775 -76521 -140731
rect -76465 -140775 -76421 -140731
rect -76365 -140775 -76321 -140731
rect -76265 -140775 -76221 -140731
rect -76165 -140775 -76121 -140731
rect -76065 -140775 -76021 -140731
rect -75965 -140775 -75921 -140731
rect -75865 -140775 -75821 -140731
rect -75765 -140775 -75721 -140731
rect -83265 -140875 -83221 -140831
rect -83165 -140875 -83121 -140831
rect -83065 -140875 -83021 -140831
rect -82965 -140875 -82921 -140831
rect -82865 -140875 -82821 -140831
rect -82765 -140875 -82721 -140831
rect -82665 -140875 -82621 -140831
rect -82565 -140875 -82521 -140831
rect -82465 -140875 -82421 -140831
rect -82365 -140875 -82321 -140831
rect -82265 -140875 -82221 -140831
rect -82165 -140875 -82121 -140831
rect -82065 -140875 -82021 -140831
rect -81965 -140875 -81921 -140831
rect -81865 -140875 -81821 -140831
rect -81765 -140875 -81721 -140831
rect -81265 -140875 -81221 -140831
rect -81165 -140875 -81121 -140831
rect -81065 -140875 -81021 -140831
rect -80965 -140875 -80921 -140831
rect -80865 -140875 -80821 -140831
rect -80765 -140875 -80721 -140831
rect -80665 -140875 -80621 -140831
rect -80565 -140875 -80521 -140831
rect -80465 -140875 -80421 -140831
rect -80365 -140875 -80321 -140831
rect -80265 -140875 -80221 -140831
rect -80165 -140875 -80121 -140831
rect -80065 -140875 -80021 -140831
rect -79965 -140875 -79921 -140831
rect -79865 -140875 -79821 -140831
rect -79765 -140875 -79721 -140831
rect -79265 -140875 -79221 -140831
rect -79165 -140875 -79121 -140831
rect -79065 -140875 -79021 -140831
rect -78965 -140875 -78921 -140831
rect -78865 -140875 -78821 -140831
rect -78765 -140875 -78721 -140831
rect -78665 -140875 -78621 -140831
rect -78565 -140875 -78521 -140831
rect -78465 -140875 -78421 -140831
rect -78365 -140875 -78321 -140831
rect -78265 -140875 -78221 -140831
rect -78165 -140875 -78121 -140831
rect -78065 -140875 -78021 -140831
rect -77965 -140875 -77921 -140831
rect -77865 -140875 -77821 -140831
rect -77765 -140875 -77721 -140831
rect -77265 -140875 -77221 -140831
rect -77165 -140875 -77121 -140831
rect -77065 -140875 -77021 -140831
rect -76965 -140875 -76921 -140831
rect -76865 -140875 -76821 -140831
rect -76765 -140875 -76721 -140831
rect -76665 -140875 -76621 -140831
rect -76565 -140875 -76521 -140831
rect -76465 -140875 -76421 -140831
rect -76365 -140875 -76321 -140831
rect -76265 -140875 -76221 -140831
rect -76165 -140875 -76121 -140831
rect -76065 -140875 -76021 -140831
rect -75965 -140875 -75921 -140831
rect -75865 -140875 -75821 -140831
rect -75765 -140875 -75721 -140831
rect -83265 -140975 -83221 -140931
rect -83165 -140975 -83121 -140931
rect -83065 -140975 -83021 -140931
rect -82965 -140975 -82921 -140931
rect -82865 -140975 -82821 -140931
rect -82765 -140975 -82721 -140931
rect -82665 -140975 -82621 -140931
rect -82565 -140975 -82521 -140931
rect -82465 -140975 -82421 -140931
rect -82365 -140975 -82321 -140931
rect -82265 -140975 -82221 -140931
rect -82165 -140975 -82121 -140931
rect -82065 -140975 -82021 -140931
rect -81965 -140975 -81921 -140931
rect -81865 -140975 -81821 -140931
rect -81765 -140975 -81721 -140931
rect -81265 -140975 -81221 -140931
rect -81165 -140975 -81121 -140931
rect -81065 -140975 -81021 -140931
rect -80965 -140975 -80921 -140931
rect -80865 -140975 -80821 -140931
rect -80765 -140975 -80721 -140931
rect -80665 -140975 -80621 -140931
rect -80565 -140975 -80521 -140931
rect -80465 -140975 -80421 -140931
rect -80365 -140975 -80321 -140931
rect -80265 -140975 -80221 -140931
rect -80165 -140975 -80121 -140931
rect -80065 -140975 -80021 -140931
rect -79965 -140975 -79921 -140931
rect -79865 -140975 -79821 -140931
rect -79765 -140975 -79721 -140931
rect -79265 -140975 -79221 -140931
rect -79165 -140975 -79121 -140931
rect -79065 -140975 -79021 -140931
rect -78965 -140975 -78921 -140931
rect -78865 -140975 -78821 -140931
rect -78765 -140975 -78721 -140931
rect -78665 -140975 -78621 -140931
rect -78565 -140975 -78521 -140931
rect -78465 -140975 -78421 -140931
rect -78365 -140975 -78321 -140931
rect -78265 -140975 -78221 -140931
rect -78165 -140975 -78121 -140931
rect -78065 -140975 -78021 -140931
rect -77965 -140975 -77921 -140931
rect -77865 -140975 -77821 -140931
rect -77765 -140975 -77721 -140931
rect -77265 -140975 -77221 -140931
rect -77165 -140975 -77121 -140931
rect -77065 -140975 -77021 -140931
rect -76965 -140975 -76921 -140931
rect -76865 -140975 -76821 -140931
rect -76765 -140975 -76721 -140931
rect -76665 -140975 -76621 -140931
rect -76565 -140975 -76521 -140931
rect -76465 -140975 -76421 -140931
rect -76365 -140975 -76321 -140931
rect -76265 -140975 -76221 -140931
rect -76165 -140975 -76121 -140931
rect -76065 -140975 -76021 -140931
rect -75965 -140975 -75921 -140931
rect -75865 -140975 -75821 -140931
rect -75765 -140975 -75721 -140931
rect -83265 -141075 -83221 -141031
rect -83165 -141075 -83121 -141031
rect -83065 -141075 -83021 -141031
rect -82965 -141075 -82921 -141031
rect -82865 -141075 -82821 -141031
rect -82765 -141075 -82721 -141031
rect -82665 -141075 -82621 -141031
rect -82565 -141075 -82521 -141031
rect -82465 -141075 -82421 -141031
rect -82365 -141075 -82321 -141031
rect -82265 -141075 -82221 -141031
rect -82165 -141075 -82121 -141031
rect -82065 -141075 -82021 -141031
rect -81965 -141075 -81921 -141031
rect -81865 -141075 -81821 -141031
rect -81765 -141075 -81721 -141031
rect -81265 -141075 -81221 -141031
rect -81165 -141075 -81121 -141031
rect -81065 -141075 -81021 -141031
rect -80965 -141075 -80921 -141031
rect -80865 -141075 -80821 -141031
rect -80765 -141075 -80721 -141031
rect -80665 -141075 -80621 -141031
rect -80565 -141075 -80521 -141031
rect -80465 -141075 -80421 -141031
rect -80365 -141075 -80321 -141031
rect -80265 -141075 -80221 -141031
rect -80165 -141075 -80121 -141031
rect -80065 -141075 -80021 -141031
rect -79965 -141075 -79921 -141031
rect -79865 -141075 -79821 -141031
rect -79765 -141075 -79721 -141031
rect -79265 -141075 -79221 -141031
rect -79165 -141075 -79121 -141031
rect -79065 -141075 -79021 -141031
rect -78965 -141075 -78921 -141031
rect -78865 -141075 -78821 -141031
rect -78765 -141075 -78721 -141031
rect -78665 -141075 -78621 -141031
rect -78565 -141075 -78521 -141031
rect -78465 -141075 -78421 -141031
rect -78365 -141075 -78321 -141031
rect -78265 -141075 -78221 -141031
rect -78165 -141075 -78121 -141031
rect -78065 -141075 -78021 -141031
rect -77965 -141075 -77921 -141031
rect -77865 -141075 -77821 -141031
rect -77765 -141075 -77721 -141031
rect -77265 -141075 -77221 -141031
rect -77165 -141075 -77121 -141031
rect -77065 -141075 -77021 -141031
rect -76965 -141075 -76921 -141031
rect -76865 -141075 -76821 -141031
rect -76765 -141075 -76721 -141031
rect -76665 -141075 -76621 -141031
rect -76565 -141075 -76521 -141031
rect -76465 -141075 -76421 -141031
rect -76365 -141075 -76321 -141031
rect -76265 -141075 -76221 -141031
rect -76165 -141075 -76121 -141031
rect -76065 -141075 -76021 -141031
rect -75965 -141075 -75921 -141031
rect -75865 -141075 -75821 -141031
rect -75765 -141075 -75721 -141031
rect -83265 -141175 -83221 -141131
rect -83165 -141175 -83121 -141131
rect -83065 -141175 -83021 -141131
rect -82965 -141175 -82921 -141131
rect -82865 -141175 -82821 -141131
rect -82765 -141175 -82721 -141131
rect -82665 -141175 -82621 -141131
rect -82565 -141175 -82521 -141131
rect -82465 -141175 -82421 -141131
rect -82365 -141175 -82321 -141131
rect -82265 -141175 -82221 -141131
rect -82165 -141175 -82121 -141131
rect -82065 -141175 -82021 -141131
rect -81965 -141175 -81921 -141131
rect -81865 -141175 -81821 -141131
rect -81765 -141175 -81721 -141131
rect -81265 -141175 -81221 -141131
rect -81165 -141175 -81121 -141131
rect -81065 -141175 -81021 -141131
rect -80965 -141175 -80921 -141131
rect -80865 -141175 -80821 -141131
rect -80765 -141175 -80721 -141131
rect -80665 -141175 -80621 -141131
rect -80565 -141175 -80521 -141131
rect -80465 -141175 -80421 -141131
rect -80365 -141175 -80321 -141131
rect -80265 -141175 -80221 -141131
rect -80165 -141175 -80121 -141131
rect -80065 -141175 -80021 -141131
rect -79965 -141175 -79921 -141131
rect -79865 -141175 -79821 -141131
rect -79765 -141175 -79721 -141131
rect -79265 -141175 -79221 -141131
rect -79165 -141175 -79121 -141131
rect -79065 -141175 -79021 -141131
rect -78965 -141175 -78921 -141131
rect -78865 -141175 -78821 -141131
rect -78765 -141175 -78721 -141131
rect -78665 -141175 -78621 -141131
rect -78565 -141175 -78521 -141131
rect -78465 -141175 -78421 -141131
rect -78365 -141175 -78321 -141131
rect -78265 -141175 -78221 -141131
rect -78165 -141175 -78121 -141131
rect -78065 -141175 -78021 -141131
rect -77965 -141175 -77921 -141131
rect -77865 -141175 -77821 -141131
rect -77765 -141175 -77721 -141131
rect -77265 -141175 -77221 -141131
rect -77165 -141175 -77121 -141131
rect -77065 -141175 -77021 -141131
rect -76965 -141175 -76921 -141131
rect -76865 -141175 -76821 -141131
rect -76765 -141175 -76721 -141131
rect -76665 -141175 -76621 -141131
rect -76565 -141175 -76521 -141131
rect -76465 -141175 -76421 -141131
rect -76365 -141175 -76321 -141131
rect -76265 -141175 -76221 -141131
rect -76165 -141175 -76121 -141131
rect -76065 -141175 -76021 -141131
rect -75965 -141175 -75921 -141131
rect -75865 -141175 -75821 -141131
rect -75765 -141175 -75721 -141131
rect -83265 -141275 -83221 -141231
rect -83165 -141275 -83121 -141231
rect -83065 -141275 -83021 -141231
rect -82965 -141275 -82921 -141231
rect -82865 -141275 -82821 -141231
rect -82765 -141275 -82721 -141231
rect -82665 -141275 -82621 -141231
rect -82565 -141275 -82521 -141231
rect -82465 -141275 -82421 -141231
rect -82365 -141275 -82321 -141231
rect -82265 -141275 -82221 -141231
rect -82165 -141275 -82121 -141231
rect -82065 -141275 -82021 -141231
rect -81965 -141275 -81921 -141231
rect -81865 -141275 -81821 -141231
rect -81765 -141275 -81721 -141231
rect -81265 -141275 -81221 -141231
rect -81165 -141275 -81121 -141231
rect -81065 -141275 -81021 -141231
rect -80965 -141275 -80921 -141231
rect -80865 -141275 -80821 -141231
rect -80765 -141275 -80721 -141231
rect -80665 -141275 -80621 -141231
rect -80565 -141275 -80521 -141231
rect -80465 -141275 -80421 -141231
rect -80365 -141275 -80321 -141231
rect -80265 -141275 -80221 -141231
rect -80165 -141275 -80121 -141231
rect -80065 -141275 -80021 -141231
rect -79965 -141275 -79921 -141231
rect -79865 -141275 -79821 -141231
rect -79765 -141275 -79721 -141231
rect -79265 -141275 -79221 -141231
rect -79165 -141275 -79121 -141231
rect -79065 -141275 -79021 -141231
rect -78965 -141275 -78921 -141231
rect -78865 -141275 -78821 -141231
rect -78765 -141275 -78721 -141231
rect -78665 -141275 -78621 -141231
rect -78565 -141275 -78521 -141231
rect -78465 -141275 -78421 -141231
rect -78365 -141275 -78321 -141231
rect -78265 -141275 -78221 -141231
rect -78165 -141275 -78121 -141231
rect -78065 -141275 -78021 -141231
rect -77965 -141275 -77921 -141231
rect -77865 -141275 -77821 -141231
rect -77765 -141275 -77721 -141231
rect -77265 -141275 -77221 -141231
rect -77165 -141275 -77121 -141231
rect -77065 -141275 -77021 -141231
rect -76965 -141275 -76921 -141231
rect -76865 -141275 -76821 -141231
rect -76765 -141275 -76721 -141231
rect -76665 -141275 -76621 -141231
rect -76565 -141275 -76521 -141231
rect -76465 -141275 -76421 -141231
rect -76365 -141275 -76321 -141231
rect -76265 -141275 -76221 -141231
rect -76165 -141275 -76121 -141231
rect -76065 -141275 -76021 -141231
rect -75965 -141275 -75921 -141231
rect -75865 -141275 -75821 -141231
rect -75765 -141275 -75721 -141231
rect -83265 -141375 -83221 -141331
rect -83165 -141375 -83121 -141331
rect -83065 -141375 -83021 -141331
rect -82965 -141375 -82921 -141331
rect -82865 -141375 -82821 -141331
rect -82765 -141375 -82721 -141331
rect -82665 -141375 -82621 -141331
rect -82565 -141375 -82521 -141331
rect -82465 -141375 -82421 -141331
rect -82365 -141375 -82321 -141331
rect -82265 -141375 -82221 -141331
rect -82165 -141375 -82121 -141331
rect -82065 -141375 -82021 -141331
rect -81965 -141375 -81921 -141331
rect -81865 -141375 -81821 -141331
rect -81765 -141375 -81721 -141331
rect -81265 -141375 -81221 -141331
rect -81165 -141375 -81121 -141331
rect -81065 -141375 -81021 -141331
rect -80965 -141375 -80921 -141331
rect -80865 -141375 -80821 -141331
rect -80765 -141375 -80721 -141331
rect -80665 -141375 -80621 -141331
rect -80565 -141375 -80521 -141331
rect -80465 -141375 -80421 -141331
rect -80365 -141375 -80321 -141331
rect -80265 -141375 -80221 -141331
rect -80165 -141375 -80121 -141331
rect -80065 -141375 -80021 -141331
rect -79965 -141375 -79921 -141331
rect -79865 -141375 -79821 -141331
rect -79765 -141375 -79721 -141331
rect -79265 -141375 -79221 -141331
rect -79165 -141375 -79121 -141331
rect -79065 -141375 -79021 -141331
rect -78965 -141375 -78921 -141331
rect -78865 -141375 -78821 -141331
rect -78765 -141375 -78721 -141331
rect -78665 -141375 -78621 -141331
rect -78565 -141375 -78521 -141331
rect -78465 -141375 -78421 -141331
rect -78365 -141375 -78321 -141331
rect -78265 -141375 -78221 -141331
rect -78165 -141375 -78121 -141331
rect -78065 -141375 -78021 -141331
rect -77965 -141375 -77921 -141331
rect -77865 -141375 -77821 -141331
rect -77765 -141375 -77721 -141331
rect -77265 -141375 -77221 -141331
rect -77165 -141375 -77121 -141331
rect -77065 -141375 -77021 -141331
rect -76965 -141375 -76921 -141331
rect -76865 -141375 -76821 -141331
rect -76765 -141375 -76721 -141331
rect -76665 -141375 -76621 -141331
rect -76565 -141375 -76521 -141331
rect -76465 -141375 -76421 -141331
rect -76365 -141375 -76321 -141331
rect -76265 -141375 -76221 -141331
rect -76165 -141375 -76121 -141331
rect -76065 -141375 -76021 -141331
rect -75965 -141375 -75921 -141331
rect -75865 -141375 -75821 -141331
rect -75765 -141375 -75721 -141331
rect -83265 -141475 -83221 -141431
rect -83165 -141475 -83121 -141431
rect -83065 -141475 -83021 -141431
rect -82965 -141475 -82921 -141431
rect -82865 -141475 -82821 -141431
rect -82765 -141475 -82721 -141431
rect -82665 -141475 -82621 -141431
rect -82565 -141475 -82521 -141431
rect -82465 -141475 -82421 -141431
rect -82365 -141475 -82321 -141431
rect -82265 -141475 -82221 -141431
rect -82165 -141475 -82121 -141431
rect -82065 -141475 -82021 -141431
rect -81965 -141475 -81921 -141431
rect -81865 -141475 -81821 -141431
rect -81765 -141475 -81721 -141431
rect -81265 -141475 -81221 -141431
rect -81165 -141475 -81121 -141431
rect -81065 -141475 -81021 -141431
rect -80965 -141475 -80921 -141431
rect -80865 -141475 -80821 -141431
rect -80765 -141475 -80721 -141431
rect -80665 -141475 -80621 -141431
rect -80565 -141475 -80521 -141431
rect -80465 -141475 -80421 -141431
rect -80365 -141475 -80321 -141431
rect -80265 -141475 -80221 -141431
rect -80165 -141475 -80121 -141431
rect -80065 -141475 -80021 -141431
rect -79965 -141475 -79921 -141431
rect -79865 -141475 -79821 -141431
rect -79765 -141475 -79721 -141431
rect -79265 -141475 -79221 -141431
rect -79165 -141475 -79121 -141431
rect -79065 -141475 -79021 -141431
rect -78965 -141475 -78921 -141431
rect -78865 -141475 -78821 -141431
rect -78765 -141475 -78721 -141431
rect -78665 -141475 -78621 -141431
rect -78565 -141475 -78521 -141431
rect -78465 -141475 -78421 -141431
rect -78365 -141475 -78321 -141431
rect -78265 -141475 -78221 -141431
rect -78165 -141475 -78121 -141431
rect -78065 -141475 -78021 -141431
rect -77965 -141475 -77921 -141431
rect -77865 -141475 -77821 -141431
rect -77765 -141475 -77721 -141431
rect -77265 -141475 -77221 -141431
rect -77165 -141475 -77121 -141431
rect -77065 -141475 -77021 -141431
rect -76965 -141475 -76921 -141431
rect -76865 -141475 -76821 -141431
rect -76765 -141475 -76721 -141431
rect -76665 -141475 -76621 -141431
rect -76565 -141475 -76521 -141431
rect -76465 -141475 -76421 -141431
rect -76365 -141475 -76321 -141431
rect -76265 -141475 -76221 -141431
rect -76165 -141475 -76121 -141431
rect -76065 -141475 -76021 -141431
rect -75965 -141475 -75921 -141431
rect -75865 -141475 -75821 -141431
rect -75765 -141475 -75721 -141431
rect -83265 -141575 -83221 -141531
rect -83165 -141575 -83121 -141531
rect -83065 -141575 -83021 -141531
rect -82965 -141575 -82921 -141531
rect -82865 -141575 -82821 -141531
rect -82765 -141575 -82721 -141531
rect -82665 -141575 -82621 -141531
rect -82565 -141575 -82521 -141531
rect -82465 -141575 -82421 -141531
rect -82365 -141575 -82321 -141531
rect -82265 -141575 -82221 -141531
rect -82165 -141575 -82121 -141531
rect -82065 -141575 -82021 -141531
rect -81965 -141575 -81921 -141531
rect -81865 -141575 -81821 -141531
rect -81765 -141575 -81721 -141531
rect -81265 -141575 -81221 -141531
rect -81165 -141575 -81121 -141531
rect -81065 -141575 -81021 -141531
rect -80965 -141575 -80921 -141531
rect -80865 -141575 -80821 -141531
rect -80765 -141575 -80721 -141531
rect -80665 -141575 -80621 -141531
rect -80565 -141575 -80521 -141531
rect -80465 -141575 -80421 -141531
rect -80365 -141575 -80321 -141531
rect -80265 -141575 -80221 -141531
rect -80165 -141575 -80121 -141531
rect -80065 -141575 -80021 -141531
rect -79965 -141575 -79921 -141531
rect -79865 -141575 -79821 -141531
rect -79765 -141575 -79721 -141531
rect -79265 -141575 -79221 -141531
rect -79165 -141575 -79121 -141531
rect -79065 -141575 -79021 -141531
rect -78965 -141575 -78921 -141531
rect -78865 -141575 -78821 -141531
rect -78765 -141575 -78721 -141531
rect -78665 -141575 -78621 -141531
rect -78565 -141575 -78521 -141531
rect -78465 -141575 -78421 -141531
rect -78365 -141575 -78321 -141531
rect -78265 -141575 -78221 -141531
rect -78165 -141575 -78121 -141531
rect -78065 -141575 -78021 -141531
rect -77965 -141575 -77921 -141531
rect -77865 -141575 -77821 -141531
rect -77765 -141575 -77721 -141531
rect -77265 -141575 -77221 -141531
rect -77165 -141575 -77121 -141531
rect -77065 -141575 -77021 -141531
rect -76965 -141575 -76921 -141531
rect -76865 -141575 -76821 -141531
rect -76765 -141575 -76721 -141531
rect -76665 -141575 -76621 -141531
rect -76565 -141575 -76521 -141531
rect -76465 -141575 -76421 -141531
rect -76365 -141575 -76321 -141531
rect -76265 -141575 -76221 -141531
rect -76165 -141575 -76121 -141531
rect -76065 -141575 -76021 -141531
rect -75965 -141575 -75921 -141531
rect -75865 -141575 -75821 -141531
rect -75765 -141575 -75721 -141531
rect -83265 -141675 -83221 -141631
rect -83165 -141675 -83121 -141631
rect -83065 -141675 -83021 -141631
rect -82965 -141675 -82921 -141631
rect -82865 -141675 -82821 -141631
rect -82765 -141675 -82721 -141631
rect -82665 -141675 -82621 -141631
rect -82565 -141675 -82521 -141631
rect -82465 -141675 -82421 -141631
rect -82365 -141675 -82321 -141631
rect -82265 -141675 -82221 -141631
rect -82165 -141675 -82121 -141631
rect -82065 -141675 -82021 -141631
rect -81965 -141675 -81921 -141631
rect -81865 -141675 -81821 -141631
rect -81765 -141675 -81721 -141631
rect -81265 -141675 -81221 -141631
rect -81165 -141675 -81121 -141631
rect -81065 -141675 -81021 -141631
rect -80965 -141675 -80921 -141631
rect -80865 -141675 -80821 -141631
rect -80765 -141675 -80721 -141631
rect -80665 -141675 -80621 -141631
rect -80565 -141675 -80521 -141631
rect -80465 -141675 -80421 -141631
rect -80365 -141675 -80321 -141631
rect -80265 -141675 -80221 -141631
rect -80165 -141675 -80121 -141631
rect -80065 -141675 -80021 -141631
rect -79965 -141675 -79921 -141631
rect -79865 -141675 -79821 -141631
rect -79765 -141675 -79721 -141631
rect -79265 -141675 -79221 -141631
rect -79165 -141675 -79121 -141631
rect -79065 -141675 -79021 -141631
rect -78965 -141675 -78921 -141631
rect -78865 -141675 -78821 -141631
rect -78765 -141675 -78721 -141631
rect -78665 -141675 -78621 -141631
rect -78565 -141675 -78521 -141631
rect -78465 -141675 -78421 -141631
rect -78365 -141675 -78321 -141631
rect -78265 -141675 -78221 -141631
rect -78165 -141675 -78121 -141631
rect -78065 -141675 -78021 -141631
rect -77965 -141675 -77921 -141631
rect -77865 -141675 -77821 -141631
rect -77765 -141675 -77721 -141631
rect -77265 -141675 -77221 -141631
rect -77165 -141675 -77121 -141631
rect -77065 -141675 -77021 -141631
rect -76965 -141675 -76921 -141631
rect -76865 -141675 -76821 -141631
rect -76765 -141675 -76721 -141631
rect -76665 -141675 -76621 -141631
rect -76565 -141675 -76521 -141631
rect -76465 -141675 -76421 -141631
rect -76365 -141675 -76321 -141631
rect -76265 -141675 -76221 -141631
rect -76165 -141675 -76121 -141631
rect -76065 -141675 -76021 -141631
rect -75965 -141675 -75921 -141631
rect -75865 -141675 -75821 -141631
rect -75765 -141675 -75721 -141631
rect -83265 -141775 -83221 -141731
rect -83165 -141775 -83121 -141731
rect -83065 -141775 -83021 -141731
rect -82965 -141775 -82921 -141731
rect -82865 -141775 -82821 -141731
rect -82765 -141775 -82721 -141731
rect -82665 -141775 -82621 -141731
rect -82565 -141775 -82521 -141731
rect -82465 -141775 -82421 -141731
rect -82365 -141775 -82321 -141731
rect -82265 -141775 -82221 -141731
rect -82165 -141775 -82121 -141731
rect -82065 -141775 -82021 -141731
rect -81965 -141775 -81921 -141731
rect -81865 -141775 -81821 -141731
rect -81765 -141775 -81721 -141731
rect -81265 -141775 -81221 -141731
rect -81165 -141775 -81121 -141731
rect -81065 -141775 -81021 -141731
rect -80965 -141775 -80921 -141731
rect -80865 -141775 -80821 -141731
rect -80765 -141775 -80721 -141731
rect -80665 -141775 -80621 -141731
rect -80565 -141775 -80521 -141731
rect -80465 -141775 -80421 -141731
rect -80365 -141775 -80321 -141731
rect -80265 -141775 -80221 -141731
rect -80165 -141775 -80121 -141731
rect -80065 -141775 -80021 -141731
rect -79965 -141775 -79921 -141731
rect -79865 -141775 -79821 -141731
rect -79765 -141775 -79721 -141731
rect -79265 -141775 -79221 -141731
rect -79165 -141775 -79121 -141731
rect -79065 -141775 -79021 -141731
rect -78965 -141775 -78921 -141731
rect -78865 -141775 -78821 -141731
rect -78765 -141775 -78721 -141731
rect -78665 -141775 -78621 -141731
rect -78565 -141775 -78521 -141731
rect -78465 -141775 -78421 -141731
rect -78365 -141775 -78321 -141731
rect -78265 -141775 -78221 -141731
rect -78165 -141775 -78121 -141731
rect -78065 -141775 -78021 -141731
rect -77965 -141775 -77921 -141731
rect -77865 -141775 -77821 -141731
rect -77765 -141775 -77721 -141731
rect -77265 -141775 -77221 -141731
rect -77165 -141775 -77121 -141731
rect -77065 -141775 -77021 -141731
rect -76965 -141775 -76921 -141731
rect -76865 -141775 -76821 -141731
rect -76765 -141775 -76721 -141731
rect -76665 -141775 -76621 -141731
rect -76565 -141775 -76521 -141731
rect -76465 -141775 -76421 -141731
rect -76365 -141775 -76321 -141731
rect -76265 -141775 -76221 -141731
rect -76165 -141775 -76121 -141731
rect -76065 -141775 -76021 -141731
rect -75965 -141775 -75921 -141731
rect -75865 -141775 -75821 -141731
rect -75765 -141775 -75721 -141731
rect 81632 -138310 81676 -138266
rect 81732 -138310 81776 -138266
rect 81832 -138310 81876 -138266
rect 81932 -138310 81976 -138266
rect 82032 -138310 82076 -138266
rect 82132 -138310 82176 -138266
rect 82232 -138310 82276 -138266
rect 82332 -138310 82376 -138266
rect 82432 -138310 82476 -138266
rect 82532 -138310 82576 -138266
rect 82632 -138310 82676 -138266
rect 82732 -138310 82776 -138266
rect 82832 -138310 82876 -138266
rect 82932 -138310 82976 -138266
rect 83032 -138310 83076 -138266
rect 83132 -138310 83176 -138266
rect 83632 -138310 83676 -138266
rect 83732 -138310 83776 -138266
rect 83832 -138310 83876 -138266
rect 83932 -138310 83976 -138266
rect 84032 -138310 84076 -138266
rect 84132 -138310 84176 -138266
rect 84232 -138310 84276 -138266
rect 84332 -138310 84376 -138266
rect 84432 -138310 84476 -138266
rect 84532 -138310 84576 -138266
rect 84632 -138310 84676 -138266
rect 84732 -138310 84776 -138266
rect 84832 -138310 84876 -138266
rect 84932 -138310 84976 -138266
rect 85032 -138310 85076 -138266
rect 85132 -138310 85176 -138266
rect 85632 -138310 85676 -138266
rect 85732 -138310 85776 -138266
rect 85832 -138310 85876 -138266
rect 85932 -138310 85976 -138266
rect 86032 -138310 86076 -138266
rect 86132 -138310 86176 -138266
rect 86232 -138310 86276 -138266
rect 86332 -138310 86376 -138266
rect 86432 -138310 86476 -138266
rect 86532 -138310 86576 -138266
rect 86632 -138310 86676 -138266
rect 86732 -138310 86776 -138266
rect 86832 -138310 86876 -138266
rect 86932 -138310 86976 -138266
rect 87032 -138310 87076 -138266
rect 87132 -138310 87176 -138266
rect 87632 -138310 87676 -138266
rect 87732 -138310 87776 -138266
rect 87832 -138310 87876 -138266
rect 87932 -138310 87976 -138266
rect 88032 -138310 88076 -138266
rect 88132 -138310 88176 -138266
rect 88232 -138310 88276 -138266
rect 88332 -138310 88376 -138266
rect 88432 -138310 88476 -138266
rect 88532 -138310 88576 -138266
rect 88632 -138310 88676 -138266
rect 88732 -138310 88776 -138266
rect 88832 -138310 88876 -138266
rect 88932 -138310 88976 -138266
rect 89032 -138310 89076 -138266
rect 89132 -138310 89176 -138266
rect 81632 -138410 81676 -138366
rect 81732 -138410 81776 -138366
rect 81832 -138410 81876 -138366
rect 81932 -138410 81976 -138366
rect 82032 -138410 82076 -138366
rect 82132 -138410 82176 -138366
rect 82232 -138410 82276 -138366
rect 82332 -138410 82376 -138366
rect 82432 -138410 82476 -138366
rect 82532 -138410 82576 -138366
rect 82632 -138410 82676 -138366
rect 82732 -138410 82776 -138366
rect 82832 -138410 82876 -138366
rect 82932 -138410 82976 -138366
rect 83032 -138410 83076 -138366
rect 83132 -138410 83176 -138366
rect 83632 -138410 83676 -138366
rect 83732 -138410 83776 -138366
rect 83832 -138410 83876 -138366
rect 83932 -138410 83976 -138366
rect 84032 -138410 84076 -138366
rect 84132 -138410 84176 -138366
rect 84232 -138410 84276 -138366
rect 84332 -138410 84376 -138366
rect 84432 -138410 84476 -138366
rect 84532 -138410 84576 -138366
rect 84632 -138410 84676 -138366
rect 84732 -138410 84776 -138366
rect 84832 -138410 84876 -138366
rect 84932 -138410 84976 -138366
rect 85032 -138410 85076 -138366
rect 85132 -138410 85176 -138366
rect 85632 -138410 85676 -138366
rect 85732 -138410 85776 -138366
rect 85832 -138410 85876 -138366
rect 85932 -138410 85976 -138366
rect 86032 -138410 86076 -138366
rect 86132 -138410 86176 -138366
rect 86232 -138410 86276 -138366
rect 86332 -138410 86376 -138366
rect 86432 -138410 86476 -138366
rect 86532 -138410 86576 -138366
rect 86632 -138410 86676 -138366
rect 86732 -138410 86776 -138366
rect 86832 -138410 86876 -138366
rect 86932 -138410 86976 -138366
rect 87032 -138410 87076 -138366
rect 87132 -138410 87176 -138366
rect 87632 -138410 87676 -138366
rect 87732 -138410 87776 -138366
rect 87832 -138410 87876 -138366
rect 87932 -138410 87976 -138366
rect 88032 -138410 88076 -138366
rect 88132 -138410 88176 -138366
rect 88232 -138410 88276 -138366
rect 88332 -138410 88376 -138366
rect 88432 -138410 88476 -138366
rect 88532 -138410 88576 -138366
rect 88632 -138410 88676 -138366
rect 88732 -138410 88776 -138366
rect 88832 -138410 88876 -138366
rect 88932 -138410 88976 -138366
rect 89032 -138410 89076 -138366
rect 89132 -138410 89176 -138366
rect 81632 -138510 81676 -138466
rect 81732 -138510 81776 -138466
rect 81832 -138510 81876 -138466
rect 81932 -138510 81976 -138466
rect 82032 -138510 82076 -138466
rect 82132 -138510 82176 -138466
rect 82232 -138510 82276 -138466
rect 82332 -138510 82376 -138466
rect 82432 -138510 82476 -138466
rect 82532 -138510 82576 -138466
rect 82632 -138510 82676 -138466
rect 82732 -138510 82776 -138466
rect 82832 -138510 82876 -138466
rect 82932 -138510 82976 -138466
rect 83032 -138510 83076 -138466
rect 83132 -138510 83176 -138466
rect 83632 -138510 83676 -138466
rect 83732 -138510 83776 -138466
rect 83832 -138510 83876 -138466
rect 83932 -138510 83976 -138466
rect 84032 -138510 84076 -138466
rect 84132 -138510 84176 -138466
rect 84232 -138510 84276 -138466
rect 84332 -138510 84376 -138466
rect 84432 -138510 84476 -138466
rect 84532 -138510 84576 -138466
rect 84632 -138510 84676 -138466
rect 84732 -138510 84776 -138466
rect 84832 -138510 84876 -138466
rect 84932 -138510 84976 -138466
rect 85032 -138510 85076 -138466
rect 85132 -138510 85176 -138466
rect 85632 -138510 85676 -138466
rect 85732 -138510 85776 -138466
rect 85832 -138510 85876 -138466
rect 85932 -138510 85976 -138466
rect 86032 -138510 86076 -138466
rect 86132 -138510 86176 -138466
rect 86232 -138510 86276 -138466
rect 86332 -138510 86376 -138466
rect 86432 -138510 86476 -138466
rect 86532 -138510 86576 -138466
rect 86632 -138510 86676 -138466
rect 86732 -138510 86776 -138466
rect 86832 -138510 86876 -138466
rect 86932 -138510 86976 -138466
rect 87032 -138510 87076 -138466
rect 87132 -138510 87176 -138466
rect 87632 -138510 87676 -138466
rect 87732 -138510 87776 -138466
rect 87832 -138510 87876 -138466
rect 87932 -138510 87976 -138466
rect 88032 -138510 88076 -138466
rect 88132 -138510 88176 -138466
rect 88232 -138510 88276 -138466
rect 88332 -138510 88376 -138466
rect 88432 -138510 88476 -138466
rect 88532 -138510 88576 -138466
rect 88632 -138510 88676 -138466
rect 88732 -138510 88776 -138466
rect 88832 -138510 88876 -138466
rect 88932 -138510 88976 -138466
rect 89032 -138510 89076 -138466
rect 89132 -138510 89176 -138466
rect 81632 -138610 81676 -138566
rect 81732 -138610 81776 -138566
rect 81832 -138610 81876 -138566
rect 81932 -138610 81976 -138566
rect 82032 -138610 82076 -138566
rect 82132 -138610 82176 -138566
rect 82232 -138610 82276 -138566
rect 82332 -138610 82376 -138566
rect 82432 -138610 82476 -138566
rect 82532 -138610 82576 -138566
rect 82632 -138610 82676 -138566
rect 82732 -138610 82776 -138566
rect 82832 -138610 82876 -138566
rect 82932 -138610 82976 -138566
rect 83032 -138610 83076 -138566
rect 83132 -138610 83176 -138566
rect 83632 -138610 83676 -138566
rect 83732 -138610 83776 -138566
rect 83832 -138610 83876 -138566
rect 83932 -138610 83976 -138566
rect 84032 -138610 84076 -138566
rect 84132 -138610 84176 -138566
rect 84232 -138610 84276 -138566
rect 84332 -138610 84376 -138566
rect 84432 -138610 84476 -138566
rect 84532 -138610 84576 -138566
rect 84632 -138610 84676 -138566
rect 84732 -138610 84776 -138566
rect 84832 -138610 84876 -138566
rect 84932 -138610 84976 -138566
rect 85032 -138610 85076 -138566
rect 85132 -138610 85176 -138566
rect 85632 -138610 85676 -138566
rect 85732 -138610 85776 -138566
rect 85832 -138610 85876 -138566
rect 85932 -138610 85976 -138566
rect 86032 -138610 86076 -138566
rect 86132 -138610 86176 -138566
rect 86232 -138610 86276 -138566
rect 86332 -138610 86376 -138566
rect 86432 -138610 86476 -138566
rect 86532 -138610 86576 -138566
rect 86632 -138610 86676 -138566
rect 86732 -138610 86776 -138566
rect 86832 -138610 86876 -138566
rect 86932 -138610 86976 -138566
rect 87032 -138610 87076 -138566
rect 87132 -138610 87176 -138566
rect 87632 -138610 87676 -138566
rect 87732 -138610 87776 -138566
rect 87832 -138610 87876 -138566
rect 87932 -138610 87976 -138566
rect 88032 -138610 88076 -138566
rect 88132 -138610 88176 -138566
rect 88232 -138610 88276 -138566
rect 88332 -138610 88376 -138566
rect 88432 -138610 88476 -138566
rect 88532 -138610 88576 -138566
rect 88632 -138610 88676 -138566
rect 88732 -138610 88776 -138566
rect 88832 -138610 88876 -138566
rect 88932 -138610 88976 -138566
rect 89032 -138610 89076 -138566
rect 89132 -138610 89176 -138566
rect 81632 -138710 81676 -138666
rect 81732 -138710 81776 -138666
rect 81832 -138710 81876 -138666
rect 81932 -138710 81976 -138666
rect 82032 -138710 82076 -138666
rect 82132 -138710 82176 -138666
rect 82232 -138710 82276 -138666
rect 82332 -138710 82376 -138666
rect 82432 -138710 82476 -138666
rect 82532 -138710 82576 -138666
rect 82632 -138710 82676 -138666
rect 82732 -138710 82776 -138666
rect 82832 -138710 82876 -138666
rect 82932 -138710 82976 -138666
rect 83032 -138710 83076 -138666
rect 83132 -138710 83176 -138666
rect 83632 -138710 83676 -138666
rect 83732 -138710 83776 -138666
rect 83832 -138710 83876 -138666
rect 83932 -138710 83976 -138666
rect 84032 -138710 84076 -138666
rect 84132 -138710 84176 -138666
rect 84232 -138710 84276 -138666
rect 84332 -138710 84376 -138666
rect 84432 -138710 84476 -138666
rect 84532 -138710 84576 -138666
rect 84632 -138710 84676 -138666
rect 84732 -138710 84776 -138666
rect 84832 -138710 84876 -138666
rect 84932 -138710 84976 -138666
rect 85032 -138710 85076 -138666
rect 85132 -138710 85176 -138666
rect 85632 -138710 85676 -138666
rect 85732 -138710 85776 -138666
rect 85832 -138710 85876 -138666
rect 85932 -138710 85976 -138666
rect 86032 -138710 86076 -138666
rect 86132 -138710 86176 -138666
rect 86232 -138710 86276 -138666
rect 86332 -138710 86376 -138666
rect 86432 -138710 86476 -138666
rect 86532 -138710 86576 -138666
rect 86632 -138710 86676 -138666
rect 86732 -138710 86776 -138666
rect 86832 -138710 86876 -138666
rect 86932 -138710 86976 -138666
rect 87032 -138710 87076 -138666
rect 87132 -138710 87176 -138666
rect 87632 -138710 87676 -138666
rect 87732 -138710 87776 -138666
rect 87832 -138710 87876 -138666
rect 87932 -138710 87976 -138666
rect 88032 -138710 88076 -138666
rect 88132 -138710 88176 -138666
rect 88232 -138710 88276 -138666
rect 88332 -138710 88376 -138666
rect 88432 -138710 88476 -138666
rect 88532 -138710 88576 -138666
rect 88632 -138710 88676 -138666
rect 88732 -138710 88776 -138666
rect 88832 -138710 88876 -138666
rect 88932 -138710 88976 -138666
rect 89032 -138710 89076 -138666
rect 89132 -138710 89176 -138666
rect 81632 -138810 81676 -138766
rect 81732 -138810 81776 -138766
rect 81832 -138810 81876 -138766
rect 81932 -138810 81976 -138766
rect 82032 -138810 82076 -138766
rect 82132 -138810 82176 -138766
rect 82232 -138810 82276 -138766
rect 82332 -138810 82376 -138766
rect 82432 -138810 82476 -138766
rect 82532 -138810 82576 -138766
rect 82632 -138810 82676 -138766
rect 82732 -138810 82776 -138766
rect 82832 -138810 82876 -138766
rect 82932 -138810 82976 -138766
rect 83032 -138810 83076 -138766
rect 83132 -138810 83176 -138766
rect 83632 -138810 83676 -138766
rect 83732 -138810 83776 -138766
rect 83832 -138810 83876 -138766
rect 83932 -138810 83976 -138766
rect 84032 -138810 84076 -138766
rect 84132 -138810 84176 -138766
rect 84232 -138810 84276 -138766
rect 84332 -138810 84376 -138766
rect 84432 -138810 84476 -138766
rect 84532 -138810 84576 -138766
rect 84632 -138810 84676 -138766
rect 84732 -138810 84776 -138766
rect 84832 -138810 84876 -138766
rect 84932 -138810 84976 -138766
rect 85032 -138810 85076 -138766
rect 85132 -138810 85176 -138766
rect 85632 -138810 85676 -138766
rect 85732 -138810 85776 -138766
rect 85832 -138810 85876 -138766
rect 85932 -138810 85976 -138766
rect 86032 -138810 86076 -138766
rect 86132 -138810 86176 -138766
rect 86232 -138810 86276 -138766
rect 86332 -138810 86376 -138766
rect 86432 -138810 86476 -138766
rect 86532 -138810 86576 -138766
rect 86632 -138810 86676 -138766
rect 86732 -138810 86776 -138766
rect 86832 -138810 86876 -138766
rect 86932 -138810 86976 -138766
rect 87032 -138810 87076 -138766
rect 87132 -138810 87176 -138766
rect 87632 -138810 87676 -138766
rect 87732 -138810 87776 -138766
rect 87832 -138810 87876 -138766
rect 87932 -138810 87976 -138766
rect 88032 -138810 88076 -138766
rect 88132 -138810 88176 -138766
rect 88232 -138810 88276 -138766
rect 88332 -138810 88376 -138766
rect 88432 -138810 88476 -138766
rect 88532 -138810 88576 -138766
rect 88632 -138810 88676 -138766
rect 88732 -138810 88776 -138766
rect 88832 -138810 88876 -138766
rect 88932 -138810 88976 -138766
rect 89032 -138810 89076 -138766
rect 89132 -138810 89176 -138766
rect 81632 -138910 81676 -138866
rect 81732 -138910 81776 -138866
rect 81832 -138910 81876 -138866
rect 81932 -138910 81976 -138866
rect 82032 -138910 82076 -138866
rect 82132 -138910 82176 -138866
rect 82232 -138910 82276 -138866
rect 82332 -138910 82376 -138866
rect 82432 -138910 82476 -138866
rect 82532 -138910 82576 -138866
rect 82632 -138910 82676 -138866
rect 82732 -138910 82776 -138866
rect 82832 -138910 82876 -138866
rect 82932 -138910 82976 -138866
rect 83032 -138910 83076 -138866
rect 83132 -138910 83176 -138866
rect 83632 -138910 83676 -138866
rect 83732 -138910 83776 -138866
rect 83832 -138910 83876 -138866
rect 83932 -138910 83976 -138866
rect 84032 -138910 84076 -138866
rect 84132 -138910 84176 -138866
rect 84232 -138910 84276 -138866
rect 84332 -138910 84376 -138866
rect 84432 -138910 84476 -138866
rect 84532 -138910 84576 -138866
rect 84632 -138910 84676 -138866
rect 84732 -138910 84776 -138866
rect 84832 -138910 84876 -138866
rect 84932 -138910 84976 -138866
rect 85032 -138910 85076 -138866
rect 85132 -138910 85176 -138866
rect 85632 -138910 85676 -138866
rect 85732 -138910 85776 -138866
rect 85832 -138910 85876 -138866
rect 85932 -138910 85976 -138866
rect 86032 -138910 86076 -138866
rect 86132 -138910 86176 -138866
rect 86232 -138910 86276 -138866
rect 86332 -138910 86376 -138866
rect 86432 -138910 86476 -138866
rect 86532 -138910 86576 -138866
rect 86632 -138910 86676 -138866
rect 86732 -138910 86776 -138866
rect 86832 -138910 86876 -138866
rect 86932 -138910 86976 -138866
rect 87032 -138910 87076 -138866
rect 87132 -138910 87176 -138866
rect 87632 -138910 87676 -138866
rect 87732 -138910 87776 -138866
rect 87832 -138910 87876 -138866
rect 87932 -138910 87976 -138866
rect 88032 -138910 88076 -138866
rect 88132 -138910 88176 -138866
rect 88232 -138910 88276 -138866
rect 88332 -138910 88376 -138866
rect 88432 -138910 88476 -138866
rect 88532 -138910 88576 -138866
rect 88632 -138910 88676 -138866
rect 88732 -138910 88776 -138866
rect 88832 -138910 88876 -138866
rect 88932 -138910 88976 -138866
rect 89032 -138910 89076 -138866
rect 89132 -138910 89176 -138866
rect 81632 -139010 81676 -138966
rect 81732 -139010 81776 -138966
rect 81832 -139010 81876 -138966
rect 81932 -139010 81976 -138966
rect 82032 -139010 82076 -138966
rect 82132 -139010 82176 -138966
rect 82232 -139010 82276 -138966
rect 82332 -139010 82376 -138966
rect 82432 -139010 82476 -138966
rect 82532 -139010 82576 -138966
rect 82632 -139010 82676 -138966
rect 82732 -139010 82776 -138966
rect 82832 -139010 82876 -138966
rect 82932 -139010 82976 -138966
rect 83032 -139010 83076 -138966
rect 83132 -139010 83176 -138966
rect 83632 -139010 83676 -138966
rect 83732 -139010 83776 -138966
rect 83832 -139010 83876 -138966
rect 83932 -139010 83976 -138966
rect 84032 -139010 84076 -138966
rect 84132 -139010 84176 -138966
rect 84232 -139010 84276 -138966
rect 84332 -139010 84376 -138966
rect 84432 -139010 84476 -138966
rect 84532 -139010 84576 -138966
rect 84632 -139010 84676 -138966
rect 84732 -139010 84776 -138966
rect 84832 -139010 84876 -138966
rect 84932 -139010 84976 -138966
rect 85032 -139010 85076 -138966
rect 85132 -139010 85176 -138966
rect 85632 -139010 85676 -138966
rect 85732 -139010 85776 -138966
rect 85832 -139010 85876 -138966
rect 85932 -139010 85976 -138966
rect 86032 -139010 86076 -138966
rect 86132 -139010 86176 -138966
rect 86232 -139010 86276 -138966
rect 86332 -139010 86376 -138966
rect 86432 -139010 86476 -138966
rect 86532 -139010 86576 -138966
rect 86632 -139010 86676 -138966
rect 86732 -139010 86776 -138966
rect 86832 -139010 86876 -138966
rect 86932 -139010 86976 -138966
rect 87032 -139010 87076 -138966
rect 87132 -139010 87176 -138966
rect 87632 -139010 87676 -138966
rect 87732 -139010 87776 -138966
rect 87832 -139010 87876 -138966
rect 87932 -139010 87976 -138966
rect 88032 -139010 88076 -138966
rect 88132 -139010 88176 -138966
rect 88232 -139010 88276 -138966
rect 88332 -139010 88376 -138966
rect 88432 -139010 88476 -138966
rect 88532 -139010 88576 -138966
rect 88632 -139010 88676 -138966
rect 88732 -139010 88776 -138966
rect 88832 -139010 88876 -138966
rect 88932 -139010 88976 -138966
rect 89032 -139010 89076 -138966
rect 89132 -139010 89176 -138966
rect 81632 -139110 81676 -139066
rect 81732 -139110 81776 -139066
rect 81832 -139110 81876 -139066
rect 81932 -139110 81976 -139066
rect 82032 -139110 82076 -139066
rect 82132 -139110 82176 -139066
rect 82232 -139110 82276 -139066
rect 82332 -139110 82376 -139066
rect 82432 -139110 82476 -139066
rect 82532 -139110 82576 -139066
rect 82632 -139110 82676 -139066
rect 82732 -139110 82776 -139066
rect 82832 -139110 82876 -139066
rect 82932 -139110 82976 -139066
rect 83032 -139110 83076 -139066
rect 83132 -139110 83176 -139066
rect 83632 -139110 83676 -139066
rect 83732 -139110 83776 -139066
rect 83832 -139110 83876 -139066
rect 83932 -139110 83976 -139066
rect 84032 -139110 84076 -139066
rect 84132 -139110 84176 -139066
rect 84232 -139110 84276 -139066
rect 84332 -139110 84376 -139066
rect 84432 -139110 84476 -139066
rect 84532 -139110 84576 -139066
rect 84632 -139110 84676 -139066
rect 84732 -139110 84776 -139066
rect 84832 -139110 84876 -139066
rect 84932 -139110 84976 -139066
rect 85032 -139110 85076 -139066
rect 85132 -139110 85176 -139066
rect 85632 -139110 85676 -139066
rect 85732 -139110 85776 -139066
rect 85832 -139110 85876 -139066
rect 85932 -139110 85976 -139066
rect 86032 -139110 86076 -139066
rect 86132 -139110 86176 -139066
rect 86232 -139110 86276 -139066
rect 86332 -139110 86376 -139066
rect 86432 -139110 86476 -139066
rect 86532 -139110 86576 -139066
rect 86632 -139110 86676 -139066
rect 86732 -139110 86776 -139066
rect 86832 -139110 86876 -139066
rect 86932 -139110 86976 -139066
rect 87032 -139110 87076 -139066
rect 87132 -139110 87176 -139066
rect 87632 -139110 87676 -139066
rect 87732 -139110 87776 -139066
rect 87832 -139110 87876 -139066
rect 87932 -139110 87976 -139066
rect 88032 -139110 88076 -139066
rect 88132 -139110 88176 -139066
rect 88232 -139110 88276 -139066
rect 88332 -139110 88376 -139066
rect 88432 -139110 88476 -139066
rect 88532 -139110 88576 -139066
rect 88632 -139110 88676 -139066
rect 88732 -139110 88776 -139066
rect 88832 -139110 88876 -139066
rect 88932 -139110 88976 -139066
rect 89032 -139110 89076 -139066
rect 89132 -139110 89176 -139066
rect 81632 -139210 81676 -139166
rect 81732 -139210 81776 -139166
rect 81832 -139210 81876 -139166
rect 81932 -139210 81976 -139166
rect 82032 -139210 82076 -139166
rect 82132 -139210 82176 -139166
rect 82232 -139210 82276 -139166
rect 82332 -139210 82376 -139166
rect 82432 -139210 82476 -139166
rect 82532 -139210 82576 -139166
rect 82632 -139210 82676 -139166
rect 82732 -139210 82776 -139166
rect 82832 -139210 82876 -139166
rect 82932 -139210 82976 -139166
rect 83032 -139210 83076 -139166
rect 83132 -139210 83176 -139166
rect 83632 -139210 83676 -139166
rect 83732 -139210 83776 -139166
rect 83832 -139210 83876 -139166
rect 83932 -139210 83976 -139166
rect 84032 -139210 84076 -139166
rect 84132 -139210 84176 -139166
rect 84232 -139210 84276 -139166
rect 84332 -139210 84376 -139166
rect 84432 -139210 84476 -139166
rect 84532 -139210 84576 -139166
rect 84632 -139210 84676 -139166
rect 84732 -139210 84776 -139166
rect 84832 -139210 84876 -139166
rect 84932 -139210 84976 -139166
rect 85032 -139210 85076 -139166
rect 85132 -139210 85176 -139166
rect 85632 -139210 85676 -139166
rect 85732 -139210 85776 -139166
rect 85832 -139210 85876 -139166
rect 85932 -139210 85976 -139166
rect 86032 -139210 86076 -139166
rect 86132 -139210 86176 -139166
rect 86232 -139210 86276 -139166
rect 86332 -139210 86376 -139166
rect 86432 -139210 86476 -139166
rect 86532 -139210 86576 -139166
rect 86632 -139210 86676 -139166
rect 86732 -139210 86776 -139166
rect 86832 -139210 86876 -139166
rect 86932 -139210 86976 -139166
rect 87032 -139210 87076 -139166
rect 87132 -139210 87176 -139166
rect 87632 -139210 87676 -139166
rect 87732 -139210 87776 -139166
rect 87832 -139210 87876 -139166
rect 87932 -139210 87976 -139166
rect 88032 -139210 88076 -139166
rect 88132 -139210 88176 -139166
rect 88232 -139210 88276 -139166
rect 88332 -139210 88376 -139166
rect 88432 -139210 88476 -139166
rect 88532 -139210 88576 -139166
rect 88632 -139210 88676 -139166
rect 88732 -139210 88776 -139166
rect 88832 -139210 88876 -139166
rect 88932 -139210 88976 -139166
rect 89032 -139210 89076 -139166
rect 89132 -139210 89176 -139166
rect 81632 -139310 81676 -139266
rect 81732 -139310 81776 -139266
rect 81832 -139310 81876 -139266
rect 81932 -139310 81976 -139266
rect 82032 -139310 82076 -139266
rect 82132 -139310 82176 -139266
rect 82232 -139310 82276 -139266
rect 82332 -139310 82376 -139266
rect 82432 -139310 82476 -139266
rect 82532 -139310 82576 -139266
rect 82632 -139310 82676 -139266
rect 82732 -139310 82776 -139266
rect 82832 -139310 82876 -139266
rect 82932 -139310 82976 -139266
rect 83032 -139310 83076 -139266
rect 83132 -139310 83176 -139266
rect 83632 -139310 83676 -139266
rect 83732 -139310 83776 -139266
rect 83832 -139310 83876 -139266
rect 83932 -139310 83976 -139266
rect 84032 -139310 84076 -139266
rect 84132 -139310 84176 -139266
rect 84232 -139310 84276 -139266
rect 84332 -139310 84376 -139266
rect 84432 -139310 84476 -139266
rect 84532 -139310 84576 -139266
rect 84632 -139310 84676 -139266
rect 84732 -139310 84776 -139266
rect 84832 -139310 84876 -139266
rect 84932 -139310 84976 -139266
rect 85032 -139310 85076 -139266
rect 85132 -139310 85176 -139266
rect 85632 -139310 85676 -139266
rect 85732 -139310 85776 -139266
rect 85832 -139310 85876 -139266
rect 85932 -139310 85976 -139266
rect 86032 -139310 86076 -139266
rect 86132 -139310 86176 -139266
rect 86232 -139310 86276 -139266
rect 86332 -139310 86376 -139266
rect 86432 -139310 86476 -139266
rect 86532 -139310 86576 -139266
rect 86632 -139310 86676 -139266
rect 86732 -139310 86776 -139266
rect 86832 -139310 86876 -139266
rect 86932 -139310 86976 -139266
rect 87032 -139310 87076 -139266
rect 87132 -139310 87176 -139266
rect 87632 -139310 87676 -139266
rect 87732 -139310 87776 -139266
rect 87832 -139310 87876 -139266
rect 87932 -139310 87976 -139266
rect 88032 -139310 88076 -139266
rect 88132 -139310 88176 -139266
rect 88232 -139310 88276 -139266
rect 88332 -139310 88376 -139266
rect 88432 -139310 88476 -139266
rect 88532 -139310 88576 -139266
rect 88632 -139310 88676 -139266
rect 88732 -139310 88776 -139266
rect 88832 -139310 88876 -139266
rect 88932 -139310 88976 -139266
rect 89032 -139310 89076 -139266
rect 89132 -139310 89176 -139266
rect 81632 -139410 81676 -139366
rect 81732 -139410 81776 -139366
rect 81832 -139410 81876 -139366
rect 81932 -139410 81976 -139366
rect 82032 -139410 82076 -139366
rect 82132 -139410 82176 -139366
rect 82232 -139410 82276 -139366
rect 82332 -139410 82376 -139366
rect 82432 -139410 82476 -139366
rect 82532 -139410 82576 -139366
rect 82632 -139410 82676 -139366
rect 82732 -139410 82776 -139366
rect 82832 -139410 82876 -139366
rect 82932 -139410 82976 -139366
rect 83032 -139410 83076 -139366
rect 83132 -139410 83176 -139366
rect 83632 -139410 83676 -139366
rect 83732 -139410 83776 -139366
rect 83832 -139410 83876 -139366
rect 83932 -139410 83976 -139366
rect 84032 -139410 84076 -139366
rect 84132 -139410 84176 -139366
rect 84232 -139410 84276 -139366
rect 84332 -139410 84376 -139366
rect 84432 -139410 84476 -139366
rect 84532 -139410 84576 -139366
rect 84632 -139410 84676 -139366
rect 84732 -139410 84776 -139366
rect 84832 -139410 84876 -139366
rect 84932 -139410 84976 -139366
rect 85032 -139410 85076 -139366
rect 85132 -139410 85176 -139366
rect 85632 -139410 85676 -139366
rect 85732 -139410 85776 -139366
rect 85832 -139410 85876 -139366
rect 85932 -139410 85976 -139366
rect 86032 -139410 86076 -139366
rect 86132 -139410 86176 -139366
rect 86232 -139410 86276 -139366
rect 86332 -139410 86376 -139366
rect 86432 -139410 86476 -139366
rect 86532 -139410 86576 -139366
rect 86632 -139410 86676 -139366
rect 86732 -139410 86776 -139366
rect 86832 -139410 86876 -139366
rect 86932 -139410 86976 -139366
rect 87032 -139410 87076 -139366
rect 87132 -139410 87176 -139366
rect 87632 -139410 87676 -139366
rect 87732 -139410 87776 -139366
rect 87832 -139410 87876 -139366
rect 87932 -139410 87976 -139366
rect 88032 -139410 88076 -139366
rect 88132 -139410 88176 -139366
rect 88232 -139410 88276 -139366
rect 88332 -139410 88376 -139366
rect 88432 -139410 88476 -139366
rect 88532 -139410 88576 -139366
rect 88632 -139410 88676 -139366
rect 88732 -139410 88776 -139366
rect 88832 -139410 88876 -139366
rect 88932 -139410 88976 -139366
rect 89032 -139410 89076 -139366
rect 89132 -139410 89176 -139366
rect 81632 -139510 81676 -139466
rect 81732 -139510 81776 -139466
rect 81832 -139510 81876 -139466
rect 81932 -139510 81976 -139466
rect 82032 -139510 82076 -139466
rect 82132 -139510 82176 -139466
rect 82232 -139510 82276 -139466
rect 82332 -139510 82376 -139466
rect 82432 -139510 82476 -139466
rect 82532 -139510 82576 -139466
rect 82632 -139510 82676 -139466
rect 82732 -139510 82776 -139466
rect 82832 -139510 82876 -139466
rect 82932 -139510 82976 -139466
rect 83032 -139510 83076 -139466
rect 83132 -139510 83176 -139466
rect 83632 -139510 83676 -139466
rect 83732 -139510 83776 -139466
rect 83832 -139510 83876 -139466
rect 83932 -139510 83976 -139466
rect 84032 -139510 84076 -139466
rect 84132 -139510 84176 -139466
rect 84232 -139510 84276 -139466
rect 84332 -139510 84376 -139466
rect 84432 -139510 84476 -139466
rect 84532 -139510 84576 -139466
rect 84632 -139510 84676 -139466
rect 84732 -139510 84776 -139466
rect 84832 -139510 84876 -139466
rect 84932 -139510 84976 -139466
rect 85032 -139510 85076 -139466
rect 85132 -139510 85176 -139466
rect 85632 -139510 85676 -139466
rect 85732 -139510 85776 -139466
rect 85832 -139510 85876 -139466
rect 85932 -139510 85976 -139466
rect 86032 -139510 86076 -139466
rect 86132 -139510 86176 -139466
rect 86232 -139510 86276 -139466
rect 86332 -139510 86376 -139466
rect 86432 -139510 86476 -139466
rect 86532 -139510 86576 -139466
rect 86632 -139510 86676 -139466
rect 86732 -139510 86776 -139466
rect 86832 -139510 86876 -139466
rect 86932 -139510 86976 -139466
rect 87032 -139510 87076 -139466
rect 87132 -139510 87176 -139466
rect 87632 -139510 87676 -139466
rect 87732 -139510 87776 -139466
rect 87832 -139510 87876 -139466
rect 87932 -139510 87976 -139466
rect 88032 -139510 88076 -139466
rect 88132 -139510 88176 -139466
rect 88232 -139510 88276 -139466
rect 88332 -139510 88376 -139466
rect 88432 -139510 88476 -139466
rect 88532 -139510 88576 -139466
rect 88632 -139510 88676 -139466
rect 88732 -139510 88776 -139466
rect 88832 -139510 88876 -139466
rect 88932 -139510 88976 -139466
rect 89032 -139510 89076 -139466
rect 89132 -139510 89176 -139466
rect 145268 -165659 145312 -165615
rect 145368 -165659 145412 -165615
rect 145468 -165659 145512 -165615
rect 145568 -165659 145612 -165615
rect 145668 -165659 145712 -165615
rect 145768 -165659 145812 -165615
rect 145868 -165659 145912 -165615
rect 145968 -165659 146012 -165615
rect 146068 -165659 146112 -165615
rect 146168 -165659 146212 -165615
rect 146268 -165659 146312 -165615
rect 146368 -165659 146412 -165615
rect 146468 -165659 146512 -165615
rect 146568 -165659 146612 -165615
rect 146668 -165659 146712 -165615
rect 146768 -165659 146812 -165615
rect 147268 -165659 147312 -165615
rect 147368 -165659 147412 -165615
rect 147468 -165659 147512 -165615
rect 147568 -165659 147612 -165615
rect 147668 -165659 147712 -165615
rect 147768 -165659 147812 -165615
rect 147868 -165659 147912 -165615
rect 147968 -165659 148012 -165615
rect 148068 -165659 148112 -165615
rect 148168 -165659 148212 -165615
rect 148268 -165659 148312 -165615
rect 148368 -165659 148412 -165615
rect 148468 -165659 148512 -165615
rect 148568 -165659 148612 -165615
rect 148668 -165659 148712 -165615
rect 148768 -165659 148812 -165615
rect 149268 -165659 149312 -165615
rect 149368 -165659 149412 -165615
rect 149468 -165659 149512 -165615
rect 149568 -165659 149612 -165615
rect 149668 -165659 149712 -165615
rect 149768 -165659 149812 -165615
rect 149868 -165659 149912 -165615
rect 149968 -165659 150012 -165615
rect 150068 -165659 150112 -165615
rect 150168 -165659 150212 -165615
rect 150268 -165659 150312 -165615
rect 150368 -165659 150412 -165615
rect 150468 -165659 150512 -165615
rect 150568 -165659 150612 -165615
rect 150668 -165659 150712 -165615
rect 150768 -165659 150812 -165615
rect 151268 -165659 151312 -165615
rect 151368 -165659 151412 -165615
rect 151468 -165659 151512 -165615
rect 151568 -165659 151612 -165615
rect 151668 -165659 151712 -165615
rect 151768 -165659 151812 -165615
rect 151868 -165659 151912 -165615
rect 151968 -165659 152012 -165615
rect 152068 -165659 152112 -165615
rect 152168 -165659 152212 -165615
rect 152268 -165659 152312 -165615
rect 152368 -165659 152412 -165615
rect 152468 -165659 152512 -165615
rect 152568 -165659 152612 -165615
rect 152668 -165659 152712 -165615
rect 152768 -165659 152812 -165615
rect 145268 -165759 145312 -165715
rect 145368 -165759 145412 -165715
rect 145468 -165759 145512 -165715
rect 145568 -165759 145612 -165715
rect 145668 -165759 145712 -165715
rect 145768 -165759 145812 -165715
rect 145868 -165759 145912 -165715
rect 145968 -165759 146012 -165715
rect 146068 -165759 146112 -165715
rect 146168 -165759 146212 -165715
rect 146268 -165759 146312 -165715
rect 146368 -165759 146412 -165715
rect 146468 -165759 146512 -165715
rect 146568 -165759 146612 -165715
rect 146668 -165759 146712 -165715
rect 146768 -165759 146812 -165715
rect 147268 -165759 147312 -165715
rect 147368 -165759 147412 -165715
rect 147468 -165759 147512 -165715
rect 147568 -165759 147612 -165715
rect 147668 -165759 147712 -165715
rect 147768 -165759 147812 -165715
rect 147868 -165759 147912 -165715
rect 147968 -165759 148012 -165715
rect 148068 -165759 148112 -165715
rect 148168 -165759 148212 -165715
rect 148268 -165759 148312 -165715
rect 148368 -165759 148412 -165715
rect 148468 -165759 148512 -165715
rect 148568 -165759 148612 -165715
rect 148668 -165759 148712 -165715
rect 148768 -165759 148812 -165715
rect 149268 -165759 149312 -165715
rect 149368 -165759 149412 -165715
rect 149468 -165759 149512 -165715
rect 149568 -165759 149612 -165715
rect 149668 -165759 149712 -165715
rect 149768 -165759 149812 -165715
rect 149868 -165759 149912 -165715
rect 149968 -165759 150012 -165715
rect 150068 -165759 150112 -165715
rect 150168 -165759 150212 -165715
rect 150268 -165759 150312 -165715
rect 150368 -165759 150412 -165715
rect 150468 -165759 150512 -165715
rect 150568 -165759 150612 -165715
rect 150668 -165759 150712 -165715
rect 150768 -165759 150812 -165715
rect 151268 -165759 151312 -165715
rect 151368 -165759 151412 -165715
rect 151468 -165759 151512 -165715
rect 151568 -165759 151612 -165715
rect 151668 -165759 151712 -165715
rect 151768 -165759 151812 -165715
rect 151868 -165759 151912 -165715
rect 151968 -165759 152012 -165715
rect 152068 -165759 152112 -165715
rect 152168 -165759 152212 -165715
rect 152268 -165759 152312 -165715
rect 152368 -165759 152412 -165715
rect 152468 -165759 152512 -165715
rect 152568 -165759 152612 -165715
rect 152668 -165759 152712 -165715
rect 152768 -165759 152812 -165715
rect 145268 -165859 145312 -165815
rect 145368 -165859 145412 -165815
rect 145468 -165859 145512 -165815
rect 145568 -165859 145612 -165815
rect 145668 -165859 145712 -165815
rect 145768 -165859 145812 -165815
rect 145868 -165859 145912 -165815
rect 145968 -165859 146012 -165815
rect 146068 -165859 146112 -165815
rect 146168 -165859 146212 -165815
rect 146268 -165859 146312 -165815
rect 146368 -165859 146412 -165815
rect 146468 -165859 146512 -165815
rect 146568 -165859 146612 -165815
rect 146668 -165859 146712 -165815
rect 146768 -165859 146812 -165815
rect 147268 -165859 147312 -165815
rect 147368 -165859 147412 -165815
rect 147468 -165859 147512 -165815
rect 147568 -165859 147612 -165815
rect 147668 -165859 147712 -165815
rect 147768 -165859 147812 -165815
rect 147868 -165859 147912 -165815
rect 147968 -165859 148012 -165815
rect 148068 -165859 148112 -165815
rect 148168 -165859 148212 -165815
rect 148268 -165859 148312 -165815
rect 148368 -165859 148412 -165815
rect 148468 -165859 148512 -165815
rect 148568 -165859 148612 -165815
rect 148668 -165859 148712 -165815
rect 148768 -165859 148812 -165815
rect 149268 -165859 149312 -165815
rect 149368 -165859 149412 -165815
rect 149468 -165859 149512 -165815
rect 149568 -165859 149612 -165815
rect 149668 -165859 149712 -165815
rect 149768 -165859 149812 -165815
rect 149868 -165859 149912 -165815
rect 149968 -165859 150012 -165815
rect 150068 -165859 150112 -165815
rect 150168 -165859 150212 -165815
rect 150268 -165859 150312 -165815
rect 150368 -165859 150412 -165815
rect 150468 -165859 150512 -165815
rect 150568 -165859 150612 -165815
rect 150668 -165859 150712 -165815
rect 150768 -165859 150812 -165815
rect 151268 -165859 151312 -165815
rect 151368 -165859 151412 -165815
rect 151468 -165859 151512 -165815
rect 151568 -165859 151612 -165815
rect 151668 -165859 151712 -165815
rect 151768 -165859 151812 -165815
rect 151868 -165859 151912 -165815
rect 151968 -165859 152012 -165815
rect 152068 -165859 152112 -165815
rect 152168 -165859 152212 -165815
rect 152268 -165859 152312 -165815
rect 152368 -165859 152412 -165815
rect 152468 -165859 152512 -165815
rect 152568 -165859 152612 -165815
rect 152668 -165859 152712 -165815
rect 152768 -165859 152812 -165815
rect 145268 -165959 145312 -165915
rect 145368 -165959 145412 -165915
rect 145468 -165959 145512 -165915
rect 145568 -165959 145612 -165915
rect 145668 -165959 145712 -165915
rect 145768 -165959 145812 -165915
rect 145868 -165959 145912 -165915
rect 145968 -165959 146012 -165915
rect 146068 -165959 146112 -165915
rect 146168 -165959 146212 -165915
rect 146268 -165959 146312 -165915
rect 146368 -165959 146412 -165915
rect 146468 -165959 146512 -165915
rect 146568 -165959 146612 -165915
rect 146668 -165959 146712 -165915
rect 146768 -165959 146812 -165915
rect 147268 -165959 147312 -165915
rect 147368 -165959 147412 -165915
rect 147468 -165959 147512 -165915
rect 147568 -165959 147612 -165915
rect 147668 -165959 147712 -165915
rect 147768 -165959 147812 -165915
rect 147868 -165959 147912 -165915
rect 147968 -165959 148012 -165915
rect 148068 -165959 148112 -165915
rect 148168 -165959 148212 -165915
rect 148268 -165959 148312 -165915
rect 148368 -165959 148412 -165915
rect 148468 -165959 148512 -165915
rect 148568 -165959 148612 -165915
rect 148668 -165959 148712 -165915
rect 148768 -165959 148812 -165915
rect 149268 -165959 149312 -165915
rect 149368 -165959 149412 -165915
rect 149468 -165959 149512 -165915
rect 149568 -165959 149612 -165915
rect 149668 -165959 149712 -165915
rect 149768 -165959 149812 -165915
rect 149868 -165959 149912 -165915
rect 149968 -165959 150012 -165915
rect 150068 -165959 150112 -165915
rect 150168 -165959 150212 -165915
rect 150268 -165959 150312 -165915
rect 150368 -165959 150412 -165915
rect 150468 -165959 150512 -165915
rect 150568 -165959 150612 -165915
rect 150668 -165959 150712 -165915
rect 150768 -165959 150812 -165915
rect 151268 -165959 151312 -165915
rect 151368 -165959 151412 -165915
rect 151468 -165959 151512 -165915
rect 151568 -165959 151612 -165915
rect 151668 -165959 151712 -165915
rect 151768 -165959 151812 -165915
rect 151868 -165959 151912 -165915
rect 151968 -165959 152012 -165915
rect 152068 -165959 152112 -165915
rect 152168 -165959 152212 -165915
rect 152268 -165959 152312 -165915
rect 152368 -165959 152412 -165915
rect 152468 -165959 152512 -165915
rect 152568 -165959 152612 -165915
rect 152668 -165959 152712 -165915
rect 152768 -165959 152812 -165915
rect 145268 -166059 145312 -166015
rect 145368 -166059 145412 -166015
rect 145468 -166059 145512 -166015
rect 145568 -166059 145612 -166015
rect 145668 -166059 145712 -166015
rect 145768 -166059 145812 -166015
rect 145868 -166059 145912 -166015
rect 145968 -166059 146012 -166015
rect 146068 -166059 146112 -166015
rect 146168 -166059 146212 -166015
rect 146268 -166059 146312 -166015
rect 146368 -166059 146412 -166015
rect 146468 -166059 146512 -166015
rect 146568 -166059 146612 -166015
rect 146668 -166059 146712 -166015
rect 146768 -166059 146812 -166015
rect 147268 -166059 147312 -166015
rect 147368 -166059 147412 -166015
rect 147468 -166059 147512 -166015
rect 147568 -166059 147612 -166015
rect 147668 -166059 147712 -166015
rect 147768 -166059 147812 -166015
rect 147868 -166059 147912 -166015
rect 147968 -166059 148012 -166015
rect 148068 -166059 148112 -166015
rect 148168 -166059 148212 -166015
rect 148268 -166059 148312 -166015
rect 148368 -166059 148412 -166015
rect 148468 -166059 148512 -166015
rect 148568 -166059 148612 -166015
rect 148668 -166059 148712 -166015
rect 148768 -166059 148812 -166015
rect 149268 -166059 149312 -166015
rect 149368 -166059 149412 -166015
rect 149468 -166059 149512 -166015
rect 149568 -166059 149612 -166015
rect 149668 -166059 149712 -166015
rect 149768 -166059 149812 -166015
rect 149868 -166059 149912 -166015
rect 149968 -166059 150012 -166015
rect 150068 -166059 150112 -166015
rect 150168 -166059 150212 -166015
rect 150268 -166059 150312 -166015
rect 150368 -166059 150412 -166015
rect 150468 -166059 150512 -166015
rect 150568 -166059 150612 -166015
rect 150668 -166059 150712 -166015
rect 150768 -166059 150812 -166015
rect 151268 -166059 151312 -166015
rect 151368 -166059 151412 -166015
rect 151468 -166059 151512 -166015
rect 151568 -166059 151612 -166015
rect 151668 -166059 151712 -166015
rect 151768 -166059 151812 -166015
rect 151868 -166059 151912 -166015
rect 151968 -166059 152012 -166015
rect 152068 -166059 152112 -166015
rect 152168 -166059 152212 -166015
rect 152268 -166059 152312 -166015
rect 152368 -166059 152412 -166015
rect 152468 -166059 152512 -166015
rect 152568 -166059 152612 -166015
rect 152668 -166059 152712 -166015
rect 152768 -166059 152812 -166015
rect 145268 -166159 145312 -166115
rect 145368 -166159 145412 -166115
rect 145468 -166159 145512 -166115
rect 145568 -166159 145612 -166115
rect 145668 -166159 145712 -166115
rect 145768 -166159 145812 -166115
rect 145868 -166159 145912 -166115
rect 145968 -166159 146012 -166115
rect 146068 -166159 146112 -166115
rect 146168 -166159 146212 -166115
rect 146268 -166159 146312 -166115
rect 146368 -166159 146412 -166115
rect 146468 -166159 146512 -166115
rect 146568 -166159 146612 -166115
rect 146668 -166159 146712 -166115
rect 146768 -166159 146812 -166115
rect 147268 -166159 147312 -166115
rect 147368 -166159 147412 -166115
rect 147468 -166159 147512 -166115
rect 147568 -166159 147612 -166115
rect 147668 -166159 147712 -166115
rect 147768 -166159 147812 -166115
rect 147868 -166159 147912 -166115
rect 147968 -166159 148012 -166115
rect 148068 -166159 148112 -166115
rect 148168 -166159 148212 -166115
rect 148268 -166159 148312 -166115
rect 148368 -166159 148412 -166115
rect 148468 -166159 148512 -166115
rect 148568 -166159 148612 -166115
rect 148668 -166159 148712 -166115
rect 148768 -166159 148812 -166115
rect 149268 -166159 149312 -166115
rect 149368 -166159 149412 -166115
rect 149468 -166159 149512 -166115
rect 149568 -166159 149612 -166115
rect 149668 -166159 149712 -166115
rect 149768 -166159 149812 -166115
rect 149868 -166159 149912 -166115
rect 149968 -166159 150012 -166115
rect 150068 -166159 150112 -166115
rect 150168 -166159 150212 -166115
rect 150268 -166159 150312 -166115
rect 150368 -166159 150412 -166115
rect 150468 -166159 150512 -166115
rect 150568 -166159 150612 -166115
rect 150668 -166159 150712 -166115
rect 150768 -166159 150812 -166115
rect 151268 -166159 151312 -166115
rect 151368 -166159 151412 -166115
rect 151468 -166159 151512 -166115
rect 151568 -166159 151612 -166115
rect 151668 -166159 151712 -166115
rect 151768 -166159 151812 -166115
rect 151868 -166159 151912 -166115
rect 151968 -166159 152012 -166115
rect 152068 -166159 152112 -166115
rect 152168 -166159 152212 -166115
rect 152268 -166159 152312 -166115
rect 152368 -166159 152412 -166115
rect 152468 -166159 152512 -166115
rect 152568 -166159 152612 -166115
rect 152668 -166159 152712 -166115
rect 152768 -166159 152812 -166115
rect 145268 -166259 145312 -166215
rect 145368 -166259 145412 -166215
rect 145468 -166259 145512 -166215
rect 145568 -166259 145612 -166215
rect 145668 -166259 145712 -166215
rect 145768 -166259 145812 -166215
rect 145868 -166259 145912 -166215
rect 145968 -166259 146012 -166215
rect 146068 -166259 146112 -166215
rect 146168 -166259 146212 -166215
rect 146268 -166259 146312 -166215
rect 146368 -166259 146412 -166215
rect 146468 -166259 146512 -166215
rect 146568 -166259 146612 -166215
rect 146668 -166259 146712 -166215
rect 146768 -166259 146812 -166215
rect 147268 -166259 147312 -166215
rect 147368 -166259 147412 -166215
rect 147468 -166259 147512 -166215
rect 147568 -166259 147612 -166215
rect 147668 -166259 147712 -166215
rect 147768 -166259 147812 -166215
rect 147868 -166259 147912 -166215
rect 147968 -166259 148012 -166215
rect 148068 -166259 148112 -166215
rect 148168 -166259 148212 -166215
rect 148268 -166259 148312 -166215
rect 148368 -166259 148412 -166215
rect 148468 -166259 148512 -166215
rect 148568 -166259 148612 -166215
rect 148668 -166259 148712 -166215
rect 148768 -166259 148812 -166215
rect 149268 -166259 149312 -166215
rect 149368 -166259 149412 -166215
rect 149468 -166259 149512 -166215
rect 149568 -166259 149612 -166215
rect 149668 -166259 149712 -166215
rect 149768 -166259 149812 -166215
rect 149868 -166259 149912 -166215
rect 149968 -166259 150012 -166215
rect 150068 -166259 150112 -166215
rect 150168 -166259 150212 -166215
rect 150268 -166259 150312 -166215
rect 150368 -166259 150412 -166215
rect 150468 -166259 150512 -166215
rect 150568 -166259 150612 -166215
rect 150668 -166259 150712 -166215
rect 150768 -166259 150812 -166215
rect 151268 -166259 151312 -166215
rect 151368 -166259 151412 -166215
rect 151468 -166259 151512 -166215
rect 151568 -166259 151612 -166215
rect 151668 -166259 151712 -166215
rect 151768 -166259 151812 -166215
rect 151868 -166259 151912 -166215
rect 151968 -166259 152012 -166215
rect 152068 -166259 152112 -166215
rect 152168 -166259 152212 -166215
rect 152268 -166259 152312 -166215
rect 152368 -166259 152412 -166215
rect 152468 -166259 152512 -166215
rect 152568 -166259 152612 -166215
rect 152668 -166259 152712 -166215
rect 152768 -166259 152812 -166215
rect 145268 -166359 145312 -166315
rect 145368 -166359 145412 -166315
rect 145468 -166359 145512 -166315
rect 145568 -166359 145612 -166315
rect 145668 -166359 145712 -166315
rect 145768 -166359 145812 -166315
rect 145868 -166359 145912 -166315
rect 145968 -166359 146012 -166315
rect 146068 -166359 146112 -166315
rect 146168 -166359 146212 -166315
rect 146268 -166359 146312 -166315
rect 146368 -166359 146412 -166315
rect 146468 -166359 146512 -166315
rect 146568 -166359 146612 -166315
rect 146668 -166359 146712 -166315
rect 146768 -166359 146812 -166315
rect 147268 -166359 147312 -166315
rect 147368 -166359 147412 -166315
rect 147468 -166359 147512 -166315
rect 147568 -166359 147612 -166315
rect 147668 -166359 147712 -166315
rect 147768 -166359 147812 -166315
rect 147868 -166359 147912 -166315
rect 147968 -166359 148012 -166315
rect 148068 -166359 148112 -166315
rect 148168 -166359 148212 -166315
rect 148268 -166359 148312 -166315
rect 148368 -166359 148412 -166315
rect 148468 -166359 148512 -166315
rect 148568 -166359 148612 -166315
rect 148668 -166359 148712 -166315
rect 148768 -166359 148812 -166315
rect 149268 -166359 149312 -166315
rect 149368 -166359 149412 -166315
rect 149468 -166359 149512 -166315
rect 149568 -166359 149612 -166315
rect 149668 -166359 149712 -166315
rect 149768 -166359 149812 -166315
rect 149868 -166359 149912 -166315
rect 149968 -166359 150012 -166315
rect 150068 -166359 150112 -166315
rect 150168 -166359 150212 -166315
rect 150268 -166359 150312 -166315
rect 150368 -166359 150412 -166315
rect 150468 -166359 150512 -166315
rect 150568 -166359 150612 -166315
rect 150668 -166359 150712 -166315
rect 150768 -166359 150812 -166315
rect 151268 -166359 151312 -166315
rect 151368 -166359 151412 -166315
rect 151468 -166359 151512 -166315
rect 151568 -166359 151612 -166315
rect 151668 -166359 151712 -166315
rect 151768 -166359 151812 -166315
rect 151868 -166359 151912 -166315
rect 151968 -166359 152012 -166315
rect 152068 -166359 152112 -166315
rect 152168 -166359 152212 -166315
rect 152268 -166359 152312 -166315
rect 152368 -166359 152412 -166315
rect 152468 -166359 152512 -166315
rect 152568 -166359 152612 -166315
rect 152668 -166359 152712 -166315
rect 152768 -166359 152812 -166315
rect 145268 -166459 145312 -166415
rect 145368 -166459 145412 -166415
rect 145468 -166459 145512 -166415
rect 145568 -166459 145612 -166415
rect 145668 -166459 145712 -166415
rect 145768 -166459 145812 -166415
rect 145868 -166459 145912 -166415
rect 145968 -166459 146012 -166415
rect 146068 -166459 146112 -166415
rect 146168 -166459 146212 -166415
rect 146268 -166459 146312 -166415
rect 146368 -166459 146412 -166415
rect 146468 -166459 146512 -166415
rect 146568 -166459 146612 -166415
rect 146668 -166459 146712 -166415
rect 146768 -166459 146812 -166415
rect 147268 -166459 147312 -166415
rect 147368 -166459 147412 -166415
rect 147468 -166459 147512 -166415
rect 147568 -166459 147612 -166415
rect 147668 -166459 147712 -166415
rect 147768 -166459 147812 -166415
rect 147868 -166459 147912 -166415
rect 147968 -166459 148012 -166415
rect 148068 -166459 148112 -166415
rect 148168 -166459 148212 -166415
rect 148268 -166459 148312 -166415
rect 148368 -166459 148412 -166415
rect 148468 -166459 148512 -166415
rect 148568 -166459 148612 -166415
rect 148668 -166459 148712 -166415
rect 148768 -166459 148812 -166415
rect 149268 -166459 149312 -166415
rect 149368 -166459 149412 -166415
rect 149468 -166459 149512 -166415
rect 149568 -166459 149612 -166415
rect 149668 -166459 149712 -166415
rect 149768 -166459 149812 -166415
rect 149868 -166459 149912 -166415
rect 149968 -166459 150012 -166415
rect 150068 -166459 150112 -166415
rect 150168 -166459 150212 -166415
rect 150268 -166459 150312 -166415
rect 150368 -166459 150412 -166415
rect 150468 -166459 150512 -166415
rect 150568 -166459 150612 -166415
rect 150668 -166459 150712 -166415
rect 150768 -166459 150812 -166415
rect 151268 -166459 151312 -166415
rect 151368 -166459 151412 -166415
rect 151468 -166459 151512 -166415
rect 151568 -166459 151612 -166415
rect 151668 -166459 151712 -166415
rect 151768 -166459 151812 -166415
rect 151868 -166459 151912 -166415
rect 151968 -166459 152012 -166415
rect 152068 -166459 152112 -166415
rect 152168 -166459 152212 -166415
rect 152268 -166459 152312 -166415
rect 152368 -166459 152412 -166415
rect 152468 -166459 152512 -166415
rect 152568 -166459 152612 -166415
rect 152668 -166459 152712 -166415
rect 152768 -166459 152812 -166415
rect 145268 -166559 145312 -166515
rect 145368 -166559 145412 -166515
rect 145468 -166559 145512 -166515
rect 145568 -166559 145612 -166515
rect 145668 -166559 145712 -166515
rect 145768 -166559 145812 -166515
rect 145868 -166559 145912 -166515
rect 145968 -166559 146012 -166515
rect 146068 -166559 146112 -166515
rect 146168 -166559 146212 -166515
rect 146268 -166559 146312 -166515
rect 146368 -166559 146412 -166515
rect 146468 -166559 146512 -166515
rect 146568 -166559 146612 -166515
rect 146668 -166559 146712 -166515
rect 146768 -166559 146812 -166515
rect 147268 -166559 147312 -166515
rect 147368 -166559 147412 -166515
rect 147468 -166559 147512 -166515
rect 147568 -166559 147612 -166515
rect 147668 -166559 147712 -166515
rect 147768 -166559 147812 -166515
rect 147868 -166559 147912 -166515
rect 147968 -166559 148012 -166515
rect 148068 -166559 148112 -166515
rect 148168 -166559 148212 -166515
rect 148268 -166559 148312 -166515
rect 148368 -166559 148412 -166515
rect 148468 -166559 148512 -166515
rect 148568 -166559 148612 -166515
rect 148668 -166559 148712 -166515
rect 148768 -166559 148812 -166515
rect 149268 -166559 149312 -166515
rect 149368 -166559 149412 -166515
rect 149468 -166559 149512 -166515
rect 149568 -166559 149612 -166515
rect 149668 -166559 149712 -166515
rect 149768 -166559 149812 -166515
rect 149868 -166559 149912 -166515
rect 149968 -166559 150012 -166515
rect 150068 -166559 150112 -166515
rect 150168 -166559 150212 -166515
rect 150268 -166559 150312 -166515
rect 150368 -166559 150412 -166515
rect 150468 -166559 150512 -166515
rect 150568 -166559 150612 -166515
rect 150668 -166559 150712 -166515
rect 150768 -166559 150812 -166515
rect 151268 -166559 151312 -166515
rect 151368 -166559 151412 -166515
rect 151468 -166559 151512 -166515
rect 151568 -166559 151612 -166515
rect 151668 -166559 151712 -166515
rect 151768 -166559 151812 -166515
rect 151868 -166559 151912 -166515
rect 151968 -166559 152012 -166515
rect 152068 -166559 152112 -166515
rect 152168 -166559 152212 -166515
rect 152268 -166559 152312 -166515
rect 152368 -166559 152412 -166515
rect 152468 -166559 152512 -166515
rect 152568 -166559 152612 -166515
rect 152668 -166559 152712 -166515
rect 152768 -166559 152812 -166515
rect 145268 -166659 145312 -166615
rect 145368 -166659 145412 -166615
rect 145468 -166659 145512 -166615
rect 145568 -166659 145612 -166615
rect 145668 -166659 145712 -166615
rect 145768 -166659 145812 -166615
rect 145868 -166659 145912 -166615
rect 145968 -166659 146012 -166615
rect 146068 -166659 146112 -166615
rect 146168 -166659 146212 -166615
rect 146268 -166659 146312 -166615
rect 146368 -166659 146412 -166615
rect 146468 -166659 146512 -166615
rect 146568 -166659 146612 -166615
rect 146668 -166659 146712 -166615
rect 146768 -166659 146812 -166615
rect 147268 -166659 147312 -166615
rect 147368 -166659 147412 -166615
rect 147468 -166659 147512 -166615
rect 147568 -166659 147612 -166615
rect 147668 -166659 147712 -166615
rect 147768 -166659 147812 -166615
rect 147868 -166659 147912 -166615
rect 147968 -166659 148012 -166615
rect 148068 -166659 148112 -166615
rect 148168 -166659 148212 -166615
rect 148268 -166659 148312 -166615
rect 148368 -166659 148412 -166615
rect 148468 -166659 148512 -166615
rect 148568 -166659 148612 -166615
rect 148668 -166659 148712 -166615
rect 148768 -166659 148812 -166615
rect 149268 -166659 149312 -166615
rect 149368 -166659 149412 -166615
rect 149468 -166659 149512 -166615
rect 149568 -166659 149612 -166615
rect 149668 -166659 149712 -166615
rect 149768 -166659 149812 -166615
rect 149868 -166659 149912 -166615
rect 149968 -166659 150012 -166615
rect 150068 -166659 150112 -166615
rect 150168 -166659 150212 -166615
rect 150268 -166659 150312 -166615
rect 150368 -166659 150412 -166615
rect 150468 -166659 150512 -166615
rect 150568 -166659 150612 -166615
rect 150668 -166659 150712 -166615
rect 150768 -166659 150812 -166615
rect 151268 -166659 151312 -166615
rect 151368 -166659 151412 -166615
rect 151468 -166659 151512 -166615
rect 151568 -166659 151612 -166615
rect 151668 -166659 151712 -166615
rect 151768 -166659 151812 -166615
rect 151868 -166659 151912 -166615
rect 151968 -166659 152012 -166615
rect 152068 -166659 152112 -166615
rect 152168 -166659 152212 -166615
rect 152268 -166659 152312 -166615
rect 152368 -166659 152412 -166615
rect 152468 -166659 152512 -166615
rect 152568 -166659 152612 -166615
rect 152668 -166659 152712 -166615
rect 152768 -166659 152812 -166615
rect 145268 -166759 145312 -166715
rect 145368 -166759 145412 -166715
rect 145468 -166759 145512 -166715
rect 145568 -166759 145612 -166715
rect 145668 -166759 145712 -166715
rect 145768 -166759 145812 -166715
rect 145868 -166759 145912 -166715
rect 145968 -166759 146012 -166715
rect 146068 -166759 146112 -166715
rect 146168 -166759 146212 -166715
rect 146268 -166759 146312 -166715
rect 146368 -166759 146412 -166715
rect 146468 -166759 146512 -166715
rect 146568 -166759 146612 -166715
rect 146668 -166759 146712 -166715
rect 146768 -166759 146812 -166715
rect 147268 -166759 147312 -166715
rect 147368 -166759 147412 -166715
rect 147468 -166759 147512 -166715
rect 147568 -166759 147612 -166715
rect 147668 -166759 147712 -166715
rect 147768 -166759 147812 -166715
rect 147868 -166759 147912 -166715
rect 147968 -166759 148012 -166715
rect 148068 -166759 148112 -166715
rect 148168 -166759 148212 -166715
rect 148268 -166759 148312 -166715
rect 148368 -166759 148412 -166715
rect 148468 -166759 148512 -166715
rect 148568 -166759 148612 -166715
rect 148668 -166759 148712 -166715
rect 148768 -166759 148812 -166715
rect 149268 -166759 149312 -166715
rect 149368 -166759 149412 -166715
rect 149468 -166759 149512 -166715
rect 149568 -166759 149612 -166715
rect 149668 -166759 149712 -166715
rect 149768 -166759 149812 -166715
rect 149868 -166759 149912 -166715
rect 149968 -166759 150012 -166715
rect 150068 -166759 150112 -166715
rect 150168 -166759 150212 -166715
rect 150268 -166759 150312 -166715
rect 150368 -166759 150412 -166715
rect 150468 -166759 150512 -166715
rect 150568 -166759 150612 -166715
rect 150668 -166759 150712 -166715
rect 150768 -166759 150812 -166715
rect 151268 -166759 151312 -166715
rect 151368 -166759 151412 -166715
rect 151468 -166759 151512 -166715
rect 151568 -166759 151612 -166715
rect 151668 -166759 151712 -166715
rect 151768 -166759 151812 -166715
rect 151868 -166759 151912 -166715
rect 151968 -166759 152012 -166715
rect 152068 -166759 152112 -166715
rect 152168 -166759 152212 -166715
rect 152268 -166759 152312 -166715
rect 152368 -166759 152412 -166715
rect 152468 -166759 152512 -166715
rect 152568 -166759 152612 -166715
rect 152668 -166759 152712 -166715
rect 152768 -166759 152812 -166715
rect 145268 -166859 145312 -166815
rect 145368 -166859 145412 -166815
rect 145468 -166859 145512 -166815
rect 145568 -166859 145612 -166815
rect 145668 -166859 145712 -166815
rect 145768 -166859 145812 -166815
rect 145868 -166859 145912 -166815
rect 145968 -166859 146012 -166815
rect 146068 -166859 146112 -166815
rect 146168 -166859 146212 -166815
rect 146268 -166859 146312 -166815
rect 146368 -166859 146412 -166815
rect 146468 -166859 146512 -166815
rect 146568 -166859 146612 -166815
rect 146668 -166859 146712 -166815
rect 146768 -166859 146812 -166815
rect 147268 -166859 147312 -166815
rect 147368 -166859 147412 -166815
rect 147468 -166859 147512 -166815
rect 147568 -166859 147612 -166815
rect 147668 -166859 147712 -166815
rect 147768 -166859 147812 -166815
rect 147868 -166859 147912 -166815
rect 147968 -166859 148012 -166815
rect 148068 -166859 148112 -166815
rect 148168 -166859 148212 -166815
rect 148268 -166859 148312 -166815
rect 148368 -166859 148412 -166815
rect 148468 -166859 148512 -166815
rect 148568 -166859 148612 -166815
rect 148668 -166859 148712 -166815
rect 148768 -166859 148812 -166815
rect 149268 -166859 149312 -166815
rect 149368 -166859 149412 -166815
rect 149468 -166859 149512 -166815
rect 149568 -166859 149612 -166815
rect 149668 -166859 149712 -166815
rect 149768 -166859 149812 -166815
rect 149868 -166859 149912 -166815
rect 149968 -166859 150012 -166815
rect 150068 -166859 150112 -166815
rect 150168 -166859 150212 -166815
rect 150268 -166859 150312 -166815
rect 150368 -166859 150412 -166815
rect 150468 -166859 150512 -166815
rect 150568 -166859 150612 -166815
rect 150668 -166859 150712 -166815
rect 150768 -166859 150812 -166815
rect 151268 -166859 151312 -166815
rect 151368 -166859 151412 -166815
rect 151468 -166859 151512 -166815
rect 151568 -166859 151612 -166815
rect 151668 -166859 151712 -166815
rect 151768 -166859 151812 -166815
rect 151868 -166859 151912 -166815
rect 151968 -166859 152012 -166815
rect 152068 -166859 152112 -166815
rect 152168 -166859 152212 -166815
rect 152268 -166859 152312 -166815
rect 152368 -166859 152412 -166815
rect 152468 -166859 152512 -166815
rect 152568 -166859 152612 -166815
rect 152668 -166859 152712 -166815
rect 152768 -166859 152812 -166815
rect 145268 -166959 145312 -166915
rect 145368 -166959 145412 -166915
rect 145468 -166959 145512 -166915
rect 145568 -166959 145612 -166915
rect 145668 -166959 145712 -166915
rect 145768 -166959 145812 -166915
rect 145868 -166959 145912 -166915
rect 145968 -166959 146012 -166915
rect 146068 -166959 146112 -166915
rect 146168 -166959 146212 -166915
rect 146268 -166959 146312 -166915
rect 146368 -166959 146412 -166915
rect 146468 -166959 146512 -166915
rect 146568 -166959 146612 -166915
rect 146668 -166959 146712 -166915
rect 146768 -166959 146812 -166915
rect 147268 -166959 147312 -166915
rect 147368 -166959 147412 -166915
rect 147468 -166959 147512 -166915
rect 147568 -166959 147612 -166915
rect 147668 -166959 147712 -166915
rect 147768 -166959 147812 -166915
rect 147868 -166959 147912 -166915
rect 147968 -166959 148012 -166915
rect 148068 -166959 148112 -166915
rect 148168 -166959 148212 -166915
rect 148268 -166959 148312 -166915
rect 148368 -166959 148412 -166915
rect 148468 -166959 148512 -166915
rect 148568 -166959 148612 -166915
rect 148668 -166959 148712 -166915
rect 148768 -166959 148812 -166915
rect 149268 -166959 149312 -166915
rect 149368 -166959 149412 -166915
rect 149468 -166959 149512 -166915
rect 149568 -166959 149612 -166915
rect 149668 -166959 149712 -166915
rect 149768 -166959 149812 -166915
rect 149868 -166959 149912 -166915
rect 149968 -166959 150012 -166915
rect 150068 -166959 150112 -166915
rect 150168 -166959 150212 -166915
rect 150268 -166959 150312 -166915
rect 150368 -166959 150412 -166915
rect 150468 -166959 150512 -166915
rect 150568 -166959 150612 -166915
rect 150668 -166959 150712 -166915
rect 150768 -166959 150812 -166915
rect 151268 -166959 151312 -166915
rect 151368 -166959 151412 -166915
rect 151468 -166959 151512 -166915
rect 151568 -166959 151612 -166915
rect 151668 -166959 151712 -166915
rect 151768 -166959 151812 -166915
rect 151868 -166959 151912 -166915
rect 151968 -166959 152012 -166915
rect 152068 -166959 152112 -166915
rect 152168 -166959 152212 -166915
rect 152268 -166959 152312 -166915
rect 152368 -166959 152412 -166915
rect 152468 -166959 152512 -166915
rect 152568 -166959 152612 -166915
rect 152668 -166959 152712 -166915
rect 152768 -166959 152812 -166915
rect 145268 -167059 145312 -167015
rect 145368 -167059 145412 -167015
rect 145468 -167059 145512 -167015
rect 145568 -167059 145612 -167015
rect 145668 -167059 145712 -167015
rect 145768 -167059 145812 -167015
rect 145868 -167059 145912 -167015
rect 145968 -167059 146012 -167015
rect 146068 -167059 146112 -167015
rect 146168 -167059 146212 -167015
rect 146268 -167059 146312 -167015
rect 146368 -167059 146412 -167015
rect 146468 -167059 146512 -167015
rect 146568 -167059 146612 -167015
rect 146668 -167059 146712 -167015
rect 146768 -167059 146812 -167015
rect 147268 -167059 147312 -167015
rect 147368 -167059 147412 -167015
rect 147468 -167059 147512 -167015
rect 147568 -167059 147612 -167015
rect 147668 -167059 147712 -167015
rect 147768 -167059 147812 -167015
rect 147868 -167059 147912 -167015
rect 147968 -167059 148012 -167015
rect 148068 -167059 148112 -167015
rect 148168 -167059 148212 -167015
rect 148268 -167059 148312 -167015
rect 148368 -167059 148412 -167015
rect 148468 -167059 148512 -167015
rect 148568 -167059 148612 -167015
rect 148668 -167059 148712 -167015
rect 148768 -167059 148812 -167015
rect 149268 -167059 149312 -167015
rect 149368 -167059 149412 -167015
rect 149468 -167059 149512 -167015
rect 149568 -167059 149612 -167015
rect 149668 -167059 149712 -167015
rect 149768 -167059 149812 -167015
rect 149868 -167059 149912 -167015
rect 149968 -167059 150012 -167015
rect 150068 -167059 150112 -167015
rect 150168 -167059 150212 -167015
rect 150268 -167059 150312 -167015
rect 150368 -167059 150412 -167015
rect 150468 -167059 150512 -167015
rect 150568 -167059 150612 -167015
rect 150668 -167059 150712 -167015
rect 150768 -167059 150812 -167015
rect 151268 -167059 151312 -167015
rect 151368 -167059 151412 -167015
rect 151468 -167059 151512 -167015
rect 151568 -167059 151612 -167015
rect 151668 -167059 151712 -167015
rect 151768 -167059 151812 -167015
rect 151868 -167059 151912 -167015
rect 151968 -167059 152012 -167015
rect 152068 -167059 152112 -167015
rect 152168 -167059 152212 -167015
rect 152268 -167059 152312 -167015
rect 152368 -167059 152412 -167015
rect 152468 -167059 152512 -167015
rect 152568 -167059 152612 -167015
rect 152668 -167059 152712 -167015
rect 152768 -167059 152812 -167015
rect 145268 -167159 145312 -167115
rect 145368 -167159 145412 -167115
rect 145468 -167159 145512 -167115
rect 145568 -167159 145612 -167115
rect 145668 -167159 145712 -167115
rect 145768 -167159 145812 -167115
rect 145868 -167159 145912 -167115
rect 145968 -167159 146012 -167115
rect 146068 -167159 146112 -167115
rect 146168 -167159 146212 -167115
rect 146268 -167159 146312 -167115
rect 146368 -167159 146412 -167115
rect 146468 -167159 146512 -167115
rect 146568 -167159 146612 -167115
rect 146668 -167159 146712 -167115
rect 146768 -167159 146812 -167115
rect 147268 -167159 147312 -167115
rect 147368 -167159 147412 -167115
rect 147468 -167159 147512 -167115
rect 147568 -167159 147612 -167115
rect 147668 -167159 147712 -167115
rect 147768 -167159 147812 -167115
rect 147868 -167159 147912 -167115
rect 147968 -167159 148012 -167115
rect 148068 -167159 148112 -167115
rect 148168 -167159 148212 -167115
rect 148268 -167159 148312 -167115
rect 148368 -167159 148412 -167115
rect 148468 -167159 148512 -167115
rect 148568 -167159 148612 -167115
rect 148668 -167159 148712 -167115
rect 148768 -167159 148812 -167115
rect 149268 -167159 149312 -167115
rect 149368 -167159 149412 -167115
rect 149468 -167159 149512 -167115
rect 149568 -167159 149612 -167115
rect 149668 -167159 149712 -167115
rect 149768 -167159 149812 -167115
rect 149868 -167159 149912 -167115
rect 149968 -167159 150012 -167115
rect 150068 -167159 150112 -167115
rect 150168 -167159 150212 -167115
rect 150268 -167159 150312 -167115
rect 150368 -167159 150412 -167115
rect 150468 -167159 150512 -167115
rect 150568 -167159 150612 -167115
rect 150668 -167159 150712 -167115
rect 150768 -167159 150812 -167115
rect 151268 -167159 151312 -167115
rect 151368 -167159 151412 -167115
rect 151468 -167159 151512 -167115
rect 151568 -167159 151612 -167115
rect 151668 -167159 151712 -167115
rect 151768 -167159 151812 -167115
rect 151868 -167159 151912 -167115
rect 151968 -167159 152012 -167115
rect 152068 -167159 152112 -167115
rect 152168 -167159 152212 -167115
rect 152268 -167159 152312 -167115
rect 152368 -167159 152412 -167115
rect 152468 -167159 152512 -167115
rect 152568 -167159 152612 -167115
rect 152668 -167159 152712 -167115
rect 152768 -167159 152812 -167115
rect 165525 -173033 165569 -172989
rect 165625 -173033 165669 -172989
rect 165725 -173033 165769 -172989
rect 165825 -173033 165869 -172989
rect 165925 -173033 165969 -172989
rect 166025 -173033 166069 -172989
rect 166125 -173033 166169 -172989
rect 166225 -173033 166269 -172989
rect 166325 -173033 166369 -172989
rect 166425 -173033 166469 -172989
rect 166525 -173033 166569 -172989
rect 166625 -173033 166669 -172989
rect 166725 -173033 166769 -172989
rect 166825 -173033 166869 -172989
rect 166925 -173033 166969 -172989
rect 167025 -173033 167069 -172989
rect 167525 -173033 167569 -172989
rect 167625 -173033 167669 -172989
rect 167725 -173033 167769 -172989
rect 167825 -173033 167869 -172989
rect 167925 -173033 167969 -172989
rect 168025 -173033 168069 -172989
rect 168125 -173033 168169 -172989
rect 168225 -173033 168269 -172989
rect 168325 -173033 168369 -172989
rect 168425 -173033 168469 -172989
rect 168525 -173033 168569 -172989
rect 168625 -173033 168669 -172989
rect 168725 -173033 168769 -172989
rect 168825 -173033 168869 -172989
rect 168925 -173033 168969 -172989
rect 169025 -173033 169069 -172989
rect 169525 -173033 169569 -172989
rect 169625 -173033 169669 -172989
rect 169725 -173033 169769 -172989
rect 169825 -173033 169869 -172989
rect 169925 -173033 169969 -172989
rect 170025 -173033 170069 -172989
rect 170125 -173033 170169 -172989
rect 170225 -173033 170269 -172989
rect 170325 -173033 170369 -172989
rect 170425 -173033 170469 -172989
rect 170525 -173033 170569 -172989
rect 170625 -173033 170669 -172989
rect 170725 -173033 170769 -172989
rect 170825 -173033 170869 -172989
rect 170925 -173033 170969 -172989
rect 171025 -173033 171069 -172989
rect 171525 -173033 171569 -172989
rect 171625 -173033 171669 -172989
rect 171725 -173033 171769 -172989
rect 171825 -173033 171869 -172989
rect 171925 -173033 171969 -172989
rect 172025 -173033 172069 -172989
rect 172125 -173033 172169 -172989
rect 172225 -173033 172269 -172989
rect 172325 -173033 172369 -172989
rect 172425 -173033 172469 -172989
rect 172525 -173033 172569 -172989
rect 172625 -173033 172669 -172989
rect 172725 -173033 172769 -172989
rect 172825 -173033 172869 -172989
rect 172925 -173033 172969 -172989
rect 173025 -173033 173069 -172989
rect 81627 -173093 81671 -173049
rect 81727 -173093 81771 -173049
rect 81827 -173093 81871 -173049
rect 81927 -173093 81971 -173049
rect 82027 -173093 82071 -173049
rect 82127 -173093 82171 -173049
rect 82227 -173093 82271 -173049
rect 82327 -173093 82371 -173049
rect 82427 -173093 82471 -173049
rect 82527 -173093 82571 -173049
rect 82627 -173093 82671 -173049
rect 82727 -173093 82771 -173049
rect 82827 -173093 82871 -173049
rect 82927 -173093 82971 -173049
rect 83027 -173093 83071 -173049
rect 83127 -173093 83171 -173049
rect 83627 -173093 83671 -173049
rect 83727 -173093 83771 -173049
rect 83827 -173093 83871 -173049
rect 83927 -173093 83971 -173049
rect 84027 -173093 84071 -173049
rect 84127 -173093 84171 -173049
rect 84227 -173093 84271 -173049
rect 84327 -173093 84371 -173049
rect 84427 -173093 84471 -173049
rect 84527 -173093 84571 -173049
rect 84627 -173093 84671 -173049
rect 84727 -173093 84771 -173049
rect 84827 -173093 84871 -173049
rect 84927 -173093 84971 -173049
rect 85027 -173093 85071 -173049
rect 85127 -173093 85171 -173049
rect 85627 -173093 85671 -173049
rect 85727 -173093 85771 -173049
rect 85827 -173093 85871 -173049
rect 85927 -173093 85971 -173049
rect 86027 -173093 86071 -173049
rect 86127 -173093 86171 -173049
rect 86227 -173093 86271 -173049
rect 86327 -173093 86371 -173049
rect 86427 -173093 86471 -173049
rect 86527 -173093 86571 -173049
rect 86627 -173093 86671 -173049
rect 86727 -173093 86771 -173049
rect 86827 -173093 86871 -173049
rect 86927 -173093 86971 -173049
rect 87027 -173093 87071 -173049
rect 87127 -173093 87171 -173049
rect 87627 -173093 87671 -173049
rect 87727 -173093 87771 -173049
rect 87827 -173093 87871 -173049
rect 87927 -173093 87971 -173049
rect 88027 -173093 88071 -173049
rect 88127 -173093 88171 -173049
rect 88227 -173093 88271 -173049
rect 88327 -173093 88371 -173049
rect 88427 -173093 88471 -173049
rect 88527 -173093 88571 -173049
rect 88627 -173093 88671 -173049
rect 88727 -173093 88771 -173049
rect 88827 -173093 88871 -173049
rect 88927 -173093 88971 -173049
rect 89027 -173093 89071 -173049
rect 89127 -173093 89171 -173049
rect 165525 -173133 165569 -173089
rect 165625 -173133 165669 -173089
rect 165725 -173133 165769 -173089
rect 165825 -173133 165869 -173089
rect 165925 -173133 165969 -173089
rect 166025 -173133 166069 -173089
rect 166125 -173133 166169 -173089
rect 166225 -173133 166269 -173089
rect 166325 -173133 166369 -173089
rect 166425 -173133 166469 -173089
rect 166525 -173133 166569 -173089
rect 166625 -173133 166669 -173089
rect 166725 -173133 166769 -173089
rect 166825 -173133 166869 -173089
rect 166925 -173133 166969 -173089
rect 167025 -173133 167069 -173089
rect 167525 -173133 167569 -173089
rect 167625 -173133 167669 -173089
rect 167725 -173133 167769 -173089
rect 167825 -173133 167869 -173089
rect 167925 -173133 167969 -173089
rect 168025 -173133 168069 -173089
rect 168125 -173133 168169 -173089
rect 168225 -173133 168269 -173089
rect 168325 -173133 168369 -173089
rect 168425 -173133 168469 -173089
rect 168525 -173133 168569 -173089
rect 168625 -173133 168669 -173089
rect 168725 -173133 168769 -173089
rect 168825 -173133 168869 -173089
rect 168925 -173133 168969 -173089
rect 169025 -173133 169069 -173089
rect 169525 -173133 169569 -173089
rect 169625 -173133 169669 -173089
rect 169725 -173133 169769 -173089
rect 169825 -173133 169869 -173089
rect 169925 -173133 169969 -173089
rect 170025 -173133 170069 -173089
rect 170125 -173133 170169 -173089
rect 170225 -173133 170269 -173089
rect 170325 -173133 170369 -173089
rect 170425 -173133 170469 -173089
rect 170525 -173133 170569 -173089
rect 170625 -173133 170669 -173089
rect 170725 -173133 170769 -173089
rect 170825 -173133 170869 -173089
rect 170925 -173133 170969 -173089
rect 171025 -173133 171069 -173089
rect 171525 -173133 171569 -173089
rect 171625 -173133 171669 -173089
rect 171725 -173133 171769 -173089
rect 171825 -173133 171869 -173089
rect 171925 -173133 171969 -173089
rect 172025 -173133 172069 -173089
rect 172125 -173133 172169 -173089
rect 172225 -173133 172269 -173089
rect 172325 -173133 172369 -173089
rect 172425 -173133 172469 -173089
rect 172525 -173133 172569 -173089
rect 172625 -173133 172669 -173089
rect 172725 -173133 172769 -173089
rect 172825 -173133 172869 -173089
rect 172925 -173133 172969 -173089
rect 173025 -173133 173069 -173089
rect 81627 -173193 81671 -173149
rect 81727 -173193 81771 -173149
rect 81827 -173193 81871 -173149
rect 81927 -173193 81971 -173149
rect 82027 -173193 82071 -173149
rect 82127 -173193 82171 -173149
rect 82227 -173193 82271 -173149
rect 82327 -173193 82371 -173149
rect 82427 -173193 82471 -173149
rect 82527 -173193 82571 -173149
rect 82627 -173193 82671 -173149
rect 82727 -173193 82771 -173149
rect 82827 -173193 82871 -173149
rect 82927 -173193 82971 -173149
rect 83027 -173193 83071 -173149
rect 83127 -173193 83171 -173149
rect 83627 -173193 83671 -173149
rect 83727 -173193 83771 -173149
rect 83827 -173193 83871 -173149
rect 83927 -173193 83971 -173149
rect 84027 -173193 84071 -173149
rect 84127 -173193 84171 -173149
rect 84227 -173193 84271 -173149
rect 84327 -173193 84371 -173149
rect 84427 -173193 84471 -173149
rect 84527 -173193 84571 -173149
rect 84627 -173193 84671 -173149
rect 84727 -173193 84771 -173149
rect 84827 -173193 84871 -173149
rect 84927 -173193 84971 -173149
rect 85027 -173193 85071 -173149
rect 85127 -173193 85171 -173149
rect 85627 -173193 85671 -173149
rect 85727 -173193 85771 -173149
rect 85827 -173193 85871 -173149
rect 85927 -173193 85971 -173149
rect 86027 -173193 86071 -173149
rect 86127 -173193 86171 -173149
rect 86227 -173193 86271 -173149
rect 86327 -173193 86371 -173149
rect 86427 -173193 86471 -173149
rect 86527 -173193 86571 -173149
rect 86627 -173193 86671 -173149
rect 86727 -173193 86771 -173149
rect 86827 -173193 86871 -173149
rect 86927 -173193 86971 -173149
rect 87027 -173193 87071 -173149
rect 87127 -173193 87171 -173149
rect 87627 -173193 87671 -173149
rect 87727 -173193 87771 -173149
rect 87827 -173193 87871 -173149
rect 87927 -173193 87971 -173149
rect 88027 -173193 88071 -173149
rect 88127 -173193 88171 -173149
rect 88227 -173193 88271 -173149
rect 88327 -173193 88371 -173149
rect 88427 -173193 88471 -173149
rect 88527 -173193 88571 -173149
rect 88627 -173193 88671 -173149
rect 88727 -173193 88771 -173149
rect 88827 -173193 88871 -173149
rect 88927 -173193 88971 -173149
rect 89027 -173193 89071 -173149
rect 89127 -173193 89171 -173149
rect 165525 -173233 165569 -173189
rect 165625 -173233 165669 -173189
rect 165725 -173233 165769 -173189
rect 165825 -173233 165869 -173189
rect 165925 -173233 165969 -173189
rect 166025 -173233 166069 -173189
rect 166125 -173233 166169 -173189
rect 166225 -173233 166269 -173189
rect 166325 -173233 166369 -173189
rect 166425 -173233 166469 -173189
rect 166525 -173233 166569 -173189
rect 166625 -173233 166669 -173189
rect 166725 -173233 166769 -173189
rect 166825 -173233 166869 -173189
rect 166925 -173233 166969 -173189
rect 167025 -173233 167069 -173189
rect 167525 -173233 167569 -173189
rect 167625 -173233 167669 -173189
rect 167725 -173233 167769 -173189
rect 167825 -173233 167869 -173189
rect 167925 -173233 167969 -173189
rect 168025 -173233 168069 -173189
rect 168125 -173233 168169 -173189
rect 168225 -173233 168269 -173189
rect 168325 -173233 168369 -173189
rect 168425 -173233 168469 -173189
rect 168525 -173233 168569 -173189
rect 168625 -173233 168669 -173189
rect 168725 -173233 168769 -173189
rect 168825 -173233 168869 -173189
rect 168925 -173233 168969 -173189
rect 169025 -173233 169069 -173189
rect 169525 -173233 169569 -173189
rect 169625 -173233 169669 -173189
rect 169725 -173233 169769 -173189
rect 169825 -173233 169869 -173189
rect 169925 -173233 169969 -173189
rect 170025 -173233 170069 -173189
rect 170125 -173233 170169 -173189
rect 170225 -173233 170269 -173189
rect 170325 -173233 170369 -173189
rect 170425 -173233 170469 -173189
rect 170525 -173233 170569 -173189
rect 170625 -173233 170669 -173189
rect 170725 -173233 170769 -173189
rect 170825 -173233 170869 -173189
rect 170925 -173233 170969 -173189
rect 171025 -173233 171069 -173189
rect 171525 -173233 171569 -173189
rect 171625 -173233 171669 -173189
rect 171725 -173233 171769 -173189
rect 171825 -173233 171869 -173189
rect 171925 -173233 171969 -173189
rect 172025 -173233 172069 -173189
rect 172125 -173233 172169 -173189
rect 172225 -173233 172269 -173189
rect 172325 -173233 172369 -173189
rect 172425 -173233 172469 -173189
rect 172525 -173233 172569 -173189
rect 172625 -173233 172669 -173189
rect 172725 -173233 172769 -173189
rect 172825 -173233 172869 -173189
rect 172925 -173233 172969 -173189
rect 173025 -173233 173069 -173189
rect 81627 -173293 81671 -173249
rect 81727 -173293 81771 -173249
rect 81827 -173293 81871 -173249
rect 81927 -173293 81971 -173249
rect 82027 -173293 82071 -173249
rect 82127 -173293 82171 -173249
rect 82227 -173293 82271 -173249
rect 82327 -173293 82371 -173249
rect 82427 -173293 82471 -173249
rect 82527 -173293 82571 -173249
rect 82627 -173293 82671 -173249
rect 82727 -173293 82771 -173249
rect 82827 -173293 82871 -173249
rect 82927 -173293 82971 -173249
rect 83027 -173293 83071 -173249
rect 83127 -173293 83171 -173249
rect 83627 -173293 83671 -173249
rect 83727 -173293 83771 -173249
rect 83827 -173293 83871 -173249
rect 83927 -173293 83971 -173249
rect 84027 -173293 84071 -173249
rect 84127 -173293 84171 -173249
rect 84227 -173293 84271 -173249
rect 84327 -173293 84371 -173249
rect 84427 -173293 84471 -173249
rect 84527 -173293 84571 -173249
rect 84627 -173293 84671 -173249
rect 84727 -173293 84771 -173249
rect 84827 -173293 84871 -173249
rect 84927 -173293 84971 -173249
rect 85027 -173293 85071 -173249
rect 85127 -173293 85171 -173249
rect 85627 -173293 85671 -173249
rect 85727 -173293 85771 -173249
rect 85827 -173293 85871 -173249
rect 85927 -173293 85971 -173249
rect 86027 -173293 86071 -173249
rect 86127 -173293 86171 -173249
rect 86227 -173293 86271 -173249
rect 86327 -173293 86371 -173249
rect 86427 -173293 86471 -173249
rect 86527 -173293 86571 -173249
rect 86627 -173293 86671 -173249
rect 86727 -173293 86771 -173249
rect 86827 -173293 86871 -173249
rect 86927 -173293 86971 -173249
rect 87027 -173293 87071 -173249
rect 87127 -173293 87171 -173249
rect 87627 -173293 87671 -173249
rect 87727 -173293 87771 -173249
rect 87827 -173293 87871 -173249
rect 87927 -173293 87971 -173249
rect 88027 -173293 88071 -173249
rect 88127 -173293 88171 -173249
rect 88227 -173293 88271 -173249
rect 88327 -173293 88371 -173249
rect 88427 -173293 88471 -173249
rect 88527 -173293 88571 -173249
rect 88627 -173293 88671 -173249
rect 88727 -173293 88771 -173249
rect 88827 -173293 88871 -173249
rect 88927 -173293 88971 -173249
rect 89027 -173293 89071 -173249
rect 89127 -173293 89171 -173249
rect 165525 -173333 165569 -173289
rect 165625 -173333 165669 -173289
rect 165725 -173333 165769 -173289
rect 165825 -173333 165869 -173289
rect 165925 -173333 165969 -173289
rect 166025 -173333 166069 -173289
rect 166125 -173333 166169 -173289
rect 166225 -173333 166269 -173289
rect 166325 -173333 166369 -173289
rect 166425 -173333 166469 -173289
rect 166525 -173333 166569 -173289
rect 166625 -173333 166669 -173289
rect 166725 -173333 166769 -173289
rect 166825 -173333 166869 -173289
rect 166925 -173333 166969 -173289
rect 167025 -173333 167069 -173289
rect 167525 -173333 167569 -173289
rect 167625 -173333 167669 -173289
rect 167725 -173333 167769 -173289
rect 167825 -173333 167869 -173289
rect 167925 -173333 167969 -173289
rect 168025 -173333 168069 -173289
rect 168125 -173333 168169 -173289
rect 168225 -173333 168269 -173289
rect 168325 -173333 168369 -173289
rect 168425 -173333 168469 -173289
rect 168525 -173333 168569 -173289
rect 168625 -173333 168669 -173289
rect 168725 -173333 168769 -173289
rect 168825 -173333 168869 -173289
rect 168925 -173333 168969 -173289
rect 169025 -173333 169069 -173289
rect 169525 -173333 169569 -173289
rect 169625 -173333 169669 -173289
rect 169725 -173333 169769 -173289
rect 169825 -173333 169869 -173289
rect 169925 -173333 169969 -173289
rect 170025 -173333 170069 -173289
rect 170125 -173333 170169 -173289
rect 170225 -173333 170269 -173289
rect 170325 -173333 170369 -173289
rect 170425 -173333 170469 -173289
rect 170525 -173333 170569 -173289
rect 170625 -173333 170669 -173289
rect 170725 -173333 170769 -173289
rect 170825 -173333 170869 -173289
rect 170925 -173333 170969 -173289
rect 171025 -173333 171069 -173289
rect 171525 -173333 171569 -173289
rect 171625 -173333 171669 -173289
rect 171725 -173333 171769 -173289
rect 171825 -173333 171869 -173289
rect 171925 -173333 171969 -173289
rect 172025 -173333 172069 -173289
rect 172125 -173333 172169 -173289
rect 172225 -173333 172269 -173289
rect 172325 -173333 172369 -173289
rect 172425 -173333 172469 -173289
rect 172525 -173333 172569 -173289
rect 172625 -173333 172669 -173289
rect 172725 -173333 172769 -173289
rect 172825 -173333 172869 -173289
rect 172925 -173333 172969 -173289
rect 173025 -173333 173069 -173289
rect 81627 -173393 81671 -173349
rect 81727 -173393 81771 -173349
rect 81827 -173393 81871 -173349
rect 81927 -173393 81971 -173349
rect 82027 -173393 82071 -173349
rect 82127 -173393 82171 -173349
rect 82227 -173393 82271 -173349
rect 82327 -173393 82371 -173349
rect 82427 -173393 82471 -173349
rect 82527 -173393 82571 -173349
rect 82627 -173393 82671 -173349
rect 82727 -173393 82771 -173349
rect 82827 -173393 82871 -173349
rect 82927 -173393 82971 -173349
rect 83027 -173393 83071 -173349
rect 83127 -173393 83171 -173349
rect 83627 -173393 83671 -173349
rect 83727 -173393 83771 -173349
rect 83827 -173393 83871 -173349
rect 83927 -173393 83971 -173349
rect 84027 -173393 84071 -173349
rect 84127 -173393 84171 -173349
rect 84227 -173393 84271 -173349
rect 84327 -173393 84371 -173349
rect 84427 -173393 84471 -173349
rect 84527 -173393 84571 -173349
rect 84627 -173393 84671 -173349
rect 84727 -173393 84771 -173349
rect 84827 -173393 84871 -173349
rect 84927 -173393 84971 -173349
rect 85027 -173393 85071 -173349
rect 85127 -173393 85171 -173349
rect 85627 -173393 85671 -173349
rect 85727 -173393 85771 -173349
rect 85827 -173393 85871 -173349
rect 85927 -173393 85971 -173349
rect 86027 -173393 86071 -173349
rect 86127 -173393 86171 -173349
rect 86227 -173393 86271 -173349
rect 86327 -173393 86371 -173349
rect 86427 -173393 86471 -173349
rect 86527 -173393 86571 -173349
rect 86627 -173393 86671 -173349
rect 86727 -173393 86771 -173349
rect 86827 -173393 86871 -173349
rect 86927 -173393 86971 -173349
rect 87027 -173393 87071 -173349
rect 87127 -173393 87171 -173349
rect 87627 -173393 87671 -173349
rect 87727 -173393 87771 -173349
rect 87827 -173393 87871 -173349
rect 87927 -173393 87971 -173349
rect 88027 -173393 88071 -173349
rect 88127 -173393 88171 -173349
rect 88227 -173393 88271 -173349
rect 88327 -173393 88371 -173349
rect 88427 -173393 88471 -173349
rect 88527 -173393 88571 -173349
rect 88627 -173393 88671 -173349
rect 88727 -173393 88771 -173349
rect 88827 -173393 88871 -173349
rect 88927 -173393 88971 -173349
rect 89027 -173393 89071 -173349
rect 89127 -173393 89171 -173349
rect 165525 -173433 165569 -173389
rect 165625 -173433 165669 -173389
rect 165725 -173433 165769 -173389
rect 165825 -173433 165869 -173389
rect 165925 -173433 165969 -173389
rect 166025 -173433 166069 -173389
rect 166125 -173433 166169 -173389
rect 166225 -173433 166269 -173389
rect 166325 -173433 166369 -173389
rect 166425 -173433 166469 -173389
rect 166525 -173433 166569 -173389
rect 166625 -173433 166669 -173389
rect 166725 -173433 166769 -173389
rect 166825 -173433 166869 -173389
rect 166925 -173433 166969 -173389
rect 167025 -173433 167069 -173389
rect 167525 -173433 167569 -173389
rect 167625 -173433 167669 -173389
rect 167725 -173433 167769 -173389
rect 167825 -173433 167869 -173389
rect 167925 -173433 167969 -173389
rect 168025 -173433 168069 -173389
rect 168125 -173433 168169 -173389
rect 168225 -173433 168269 -173389
rect 168325 -173433 168369 -173389
rect 168425 -173433 168469 -173389
rect 168525 -173433 168569 -173389
rect 168625 -173433 168669 -173389
rect 168725 -173433 168769 -173389
rect 168825 -173433 168869 -173389
rect 168925 -173433 168969 -173389
rect 169025 -173433 169069 -173389
rect 169525 -173433 169569 -173389
rect 169625 -173433 169669 -173389
rect 169725 -173433 169769 -173389
rect 169825 -173433 169869 -173389
rect 169925 -173433 169969 -173389
rect 170025 -173433 170069 -173389
rect 170125 -173433 170169 -173389
rect 170225 -173433 170269 -173389
rect 170325 -173433 170369 -173389
rect 170425 -173433 170469 -173389
rect 170525 -173433 170569 -173389
rect 170625 -173433 170669 -173389
rect 170725 -173433 170769 -173389
rect 170825 -173433 170869 -173389
rect 170925 -173433 170969 -173389
rect 171025 -173433 171069 -173389
rect 171525 -173433 171569 -173389
rect 171625 -173433 171669 -173389
rect 171725 -173433 171769 -173389
rect 171825 -173433 171869 -173389
rect 171925 -173433 171969 -173389
rect 172025 -173433 172069 -173389
rect 172125 -173433 172169 -173389
rect 172225 -173433 172269 -173389
rect 172325 -173433 172369 -173389
rect 172425 -173433 172469 -173389
rect 172525 -173433 172569 -173389
rect 172625 -173433 172669 -173389
rect 172725 -173433 172769 -173389
rect 172825 -173433 172869 -173389
rect 172925 -173433 172969 -173389
rect 173025 -173433 173069 -173389
rect 81627 -173493 81671 -173449
rect 81727 -173493 81771 -173449
rect 81827 -173493 81871 -173449
rect 81927 -173493 81971 -173449
rect 82027 -173493 82071 -173449
rect 82127 -173493 82171 -173449
rect 82227 -173493 82271 -173449
rect 82327 -173493 82371 -173449
rect 82427 -173493 82471 -173449
rect 82527 -173493 82571 -173449
rect 82627 -173493 82671 -173449
rect 82727 -173493 82771 -173449
rect 82827 -173493 82871 -173449
rect 82927 -173493 82971 -173449
rect 83027 -173493 83071 -173449
rect 83127 -173493 83171 -173449
rect 83627 -173493 83671 -173449
rect 83727 -173493 83771 -173449
rect 83827 -173493 83871 -173449
rect 83927 -173493 83971 -173449
rect 84027 -173493 84071 -173449
rect 84127 -173493 84171 -173449
rect 84227 -173493 84271 -173449
rect 84327 -173493 84371 -173449
rect 84427 -173493 84471 -173449
rect 84527 -173493 84571 -173449
rect 84627 -173493 84671 -173449
rect 84727 -173493 84771 -173449
rect 84827 -173493 84871 -173449
rect 84927 -173493 84971 -173449
rect 85027 -173493 85071 -173449
rect 85127 -173493 85171 -173449
rect 85627 -173493 85671 -173449
rect 85727 -173493 85771 -173449
rect 85827 -173493 85871 -173449
rect 85927 -173493 85971 -173449
rect 86027 -173493 86071 -173449
rect 86127 -173493 86171 -173449
rect 86227 -173493 86271 -173449
rect 86327 -173493 86371 -173449
rect 86427 -173493 86471 -173449
rect 86527 -173493 86571 -173449
rect 86627 -173493 86671 -173449
rect 86727 -173493 86771 -173449
rect 86827 -173493 86871 -173449
rect 86927 -173493 86971 -173449
rect 87027 -173493 87071 -173449
rect 87127 -173493 87171 -173449
rect 87627 -173493 87671 -173449
rect 87727 -173493 87771 -173449
rect 87827 -173493 87871 -173449
rect 87927 -173493 87971 -173449
rect 88027 -173493 88071 -173449
rect 88127 -173493 88171 -173449
rect 88227 -173493 88271 -173449
rect 88327 -173493 88371 -173449
rect 88427 -173493 88471 -173449
rect 88527 -173493 88571 -173449
rect 88627 -173493 88671 -173449
rect 88727 -173493 88771 -173449
rect 88827 -173493 88871 -173449
rect 88927 -173493 88971 -173449
rect 89027 -173493 89071 -173449
rect 89127 -173493 89171 -173449
rect 165525 -173533 165569 -173489
rect 165625 -173533 165669 -173489
rect 165725 -173533 165769 -173489
rect 165825 -173533 165869 -173489
rect 165925 -173533 165969 -173489
rect 166025 -173533 166069 -173489
rect 166125 -173533 166169 -173489
rect 166225 -173533 166269 -173489
rect 166325 -173533 166369 -173489
rect 166425 -173533 166469 -173489
rect 166525 -173533 166569 -173489
rect 166625 -173533 166669 -173489
rect 166725 -173533 166769 -173489
rect 166825 -173533 166869 -173489
rect 166925 -173533 166969 -173489
rect 167025 -173533 167069 -173489
rect 167525 -173533 167569 -173489
rect 167625 -173533 167669 -173489
rect 167725 -173533 167769 -173489
rect 167825 -173533 167869 -173489
rect 167925 -173533 167969 -173489
rect 168025 -173533 168069 -173489
rect 168125 -173533 168169 -173489
rect 168225 -173533 168269 -173489
rect 168325 -173533 168369 -173489
rect 168425 -173533 168469 -173489
rect 168525 -173533 168569 -173489
rect 168625 -173533 168669 -173489
rect 168725 -173533 168769 -173489
rect 168825 -173533 168869 -173489
rect 168925 -173533 168969 -173489
rect 169025 -173533 169069 -173489
rect 169525 -173533 169569 -173489
rect 169625 -173533 169669 -173489
rect 169725 -173533 169769 -173489
rect 169825 -173533 169869 -173489
rect 169925 -173533 169969 -173489
rect 170025 -173533 170069 -173489
rect 170125 -173533 170169 -173489
rect 170225 -173533 170269 -173489
rect 170325 -173533 170369 -173489
rect 170425 -173533 170469 -173489
rect 170525 -173533 170569 -173489
rect 170625 -173533 170669 -173489
rect 170725 -173533 170769 -173489
rect 170825 -173533 170869 -173489
rect 170925 -173533 170969 -173489
rect 171025 -173533 171069 -173489
rect 171525 -173533 171569 -173489
rect 171625 -173533 171669 -173489
rect 171725 -173533 171769 -173489
rect 171825 -173533 171869 -173489
rect 171925 -173533 171969 -173489
rect 172025 -173533 172069 -173489
rect 172125 -173533 172169 -173489
rect 172225 -173533 172269 -173489
rect 172325 -173533 172369 -173489
rect 172425 -173533 172469 -173489
rect 172525 -173533 172569 -173489
rect 172625 -173533 172669 -173489
rect 172725 -173533 172769 -173489
rect 172825 -173533 172869 -173489
rect 172925 -173533 172969 -173489
rect 173025 -173533 173069 -173489
rect 81627 -173593 81671 -173549
rect 81727 -173593 81771 -173549
rect 81827 -173593 81871 -173549
rect 81927 -173593 81971 -173549
rect 82027 -173593 82071 -173549
rect 82127 -173593 82171 -173549
rect 82227 -173593 82271 -173549
rect 82327 -173593 82371 -173549
rect 82427 -173593 82471 -173549
rect 82527 -173593 82571 -173549
rect 82627 -173593 82671 -173549
rect 82727 -173593 82771 -173549
rect 82827 -173593 82871 -173549
rect 82927 -173593 82971 -173549
rect 83027 -173593 83071 -173549
rect 83127 -173593 83171 -173549
rect 83627 -173593 83671 -173549
rect 83727 -173593 83771 -173549
rect 83827 -173593 83871 -173549
rect 83927 -173593 83971 -173549
rect 84027 -173593 84071 -173549
rect 84127 -173593 84171 -173549
rect 84227 -173593 84271 -173549
rect 84327 -173593 84371 -173549
rect 84427 -173593 84471 -173549
rect 84527 -173593 84571 -173549
rect 84627 -173593 84671 -173549
rect 84727 -173593 84771 -173549
rect 84827 -173593 84871 -173549
rect 84927 -173593 84971 -173549
rect 85027 -173593 85071 -173549
rect 85127 -173593 85171 -173549
rect 85627 -173593 85671 -173549
rect 85727 -173593 85771 -173549
rect 85827 -173593 85871 -173549
rect 85927 -173593 85971 -173549
rect 86027 -173593 86071 -173549
rect 86127 -173593 86171 -173549
rect 86227 -173593 86271 -173549
rect 86327 -173593 86371 -173549
rect 86427 -173593 86471 -173549
rect 86527 -173593 86571 -173549
rect 86627 -173593 86671 -173549
rect 86727 -173593 86771 -173549
rect 86827 -173593 86871 -173549
rect 86927 -173593 86971 -173549
rect 87027 -173593 87071 -173549
rect 87127 -173593 87171 -173549
rect 87627 -173593 87671 -173549
rect 87727 -173593 87771 -173549
rect 87827 -173593 87871 -173549
rect 87927 -173593 87971 -173549
rect 88027 -173593 88071 -173549
rect 88127 -173593 88171 -173549
rect 88227 -173593 88271 -173549
rect 88327 -173593 88371 -173549
rect 88427 -173593 88471 -173549
rect 88527 -173593 88571 -173549
rect 88627 -173593 88671 -173549
rect 88727 -173593 88771 -173549
rect 88827 -173593 88871 -173549
rect 88927 -173593 88971 -173549
rect 89027 -173593 89071 -173549
rect 89127 -173593 89171 -173549
rect 165525 -173633 165569 -173589
rect 165625 -173633 165669 -173589
rect 165725 -173633 165769 -173589
rect 165825 -173633 165869 -173589
rect 165925 -173633 165969 -173589
rect 166025 -173633 166069 -173589
rect 166125 -173633 166169 -173589
rect 166225 -173633 166269 -173589
rect 166325 -173633 166369 -173589
rect 166425 -173633 166469 -173589
rect 166525 -173633 166569 -173589
rect 166625 -173633 166669 -173589
rect 166725 -173633 166769 -173589
rect 166825 -173633 166869 -173589
rect 166925 -173633 166969 -173589
rect 167025 -173633 167069 -173589
rect 167525 -173633 167569 -173589
rect 167625 -173633 167669 -173589
rect 167725 -173633 167769 -173589
rect 167825 -173633 167869 -173589
rect 167925 -173633 167969 -173589
rect 168025 -173633 168069 -173589
rect 168125 -173633 168169 -173589
rect 168225 -173633 168269 -173589
rect 168325 -173633 168369 -173589
rect 168425 -173633 168469 -173589
rect 168525 -173633 168569 -173589
rect 168625 -173633 168669 -173589
rect 168725 -173633 168769 -173589
rect 168825 -173633 168869 -173589
rect 168925 -173633 168969 -173589
rect 169025 -173633 169069 -173589
rect 169525 -173633 169569 -173589
rect 169625 -173633 169669 -173589
rect 169725 -173633 169769 -173589
rect 169825 -173633 169869 -173589
rect 169925 -173633 169969 -173589
rect 170025 -173633 170069 -173589
rect 170125 -173633 170169 -173589
rect 170225 -173633 170269 -173589
rect 170325 -173633 170369 -173589
rect 170425 -173633 170469 -173589
rect 170525 -173633 170569 -173589
rect 170625 -173633 170669 -173589
rect 170725 -173633 170769 -173589
rect 170825 -173633 170869 -173589
rect 170925 -173633 170969 -173589
rect 171025 -173633 171069 -173589
rect 171525 -173633 171569 -173589
rect 171625 -173633 171669 -173589
rect 171725 -173633 171769 -173589
rect 171825 -173633 171869 -173589
rect 171925 -173633 171969 -173589
rect 172025 -173633 172069 -173589
rect 172125 -173633 172169 -173589
rect 172225 -173633 172269 -173589
rect 172325 -173633 172369 -173589
rect 172425 -173633 172469 -173589
rect 172525 -173633 172569 -173589
rect 172625 -173633 172669 -173589
rect 172725 -173633 172769 -173589
rect 172825 -173633 172869 -173589
rect 172925 -173633 172969 -173589
rect 173025 -173633 173069 -173589
rect 81627 -173693 81671 -173649
rect 81727 -173693 81771 -173649
rect 81827 -173693 81871 -173649
rect 81927 -173693 81971 -173649
rect 82027 -173693 82071 -173649
rect 82127 -173693 82171 -173649
rect 82227 -173693 82271 -173649
rect 82327 -173693 82371 -173649
rect 82427 -173693 82471 -173649
rect 82527 -173693 82571 -173649
rect 82627 -173693 82671 -173649
rect 82727 -173693 82771 -173649
rect 82827 -173693 82871 -173649
rect 82927 -173693 82971 -173649
rect 83027 -173693 83071 -173649
rect 83127 -173693 83171 -173649
rect 83627 -173693 83671 -173649
rect 83727 -173693 83771 -173649
rect 83827 -173693 83871 -173649
rect 83927 -173693 83971 -173649
rect 84027 -173693 84071 -173649
rect 84127 -173693 84171 -173649
rect 84227 -173693 84271 -173649
rect 84327 -173693 84371 -173649
rect 84427 -173693 84471 -173649
rect 84527 -173693 84571 -173649
rect 84627 -173693 84671 -173649
rect 84727 -173693 84771 -173649
rect 84827 -173693 84871 -173649
rect 84927 -173693 84971 -173649
rect 85027 -173693 85071 -173649
rect 85127 -173693 85171 -173649
rect 85627 -173693 85671 -173649
rect 85727 -173693 85771 -173649
rect 85827 -173693 85871 -173649
rect 85927 -173693 85971 -173649
rect 86027 -173693 86071 -173649
rect 86127 -173693 86171 -173649
rect 86227 -173693 86271 -173649
rect 86327 -173693 86371 -173649
rect 86427 -173693 86471 -173649
rect 86527 -173693 86571 -173649
rect 86627 -173693 86671 -173649
rect 86727 -173693 86771 -173649
rect 86827 -173693 86871 -173649
rect 86927 -173693 86971 -173649
rect 87027 -173693 87071 -173649
rect 87127 -173693 87171 -173649
rect 87627 -173693 87671 -173649
rect 87727 -173693 87771 -173649
rect 87827 -173693 87871 -173649
rect 87927 -173693 87971 -173649
rect 88027 -173693 88071 -173649
rect 88127 -173693 88171 -173649
rect 88227 -173693 88271 -173649
rect 88327 -173693 88371 -173649
rect 88427 -173693 88471 -173649
rect 88527 -173693 88571 -173649
rect 88627 -173693 88671 -173649
rect 88727 -173693 88771 -173649
rect 88827 -173693 88871 -173649
rect 88927 -173693 88971 -173649
rect 89027 -173693 89071 -173649
rect 89127 -173693 89171 -173649
rect 165525 -173733 165569 -173689
rect 165625 -173733 165669 -173689
rect 165725 -173733 165769 -173689
rect 165825 -173733 165869 -173689
rect 165925 -173733 165969 -173689
rect 166025 -173733 166069 -173689
rect 166125 -173733 166169 -173689
rect 166225 -173733 166269 -173689
rect 166325 -173733 166369 -173689
rect 166425 -173733 166469 -173689
rect 166525 -173733 166569 -173689
rect 166625 -173733 166669 -173689
rect 166725 -173733 166769 -173689
rect 166825 -173733 166869 -173689
rect 166925 -173733 166969 -173689
rect 167025 -173733 167069 -173689
rect 167525 -173733 167569 -173689
rect 167625 -173733 167669 -173689
rect 167725 -173733 167769 -173689
rect 167825 -173733 167869 -173689
rect 167925 -173733 167969 -173689
rect 168025 -173733 168069 -173689
rect 168125 -173733 168169 -173689
rect 168225 -173733 168269 -173689
rect 168325 -173733 168369 -173689
rect 168425 -173733 168469 -173689
rect 168525 -173733 168569 -173689
rect 168625 -173733 168669 -173689
rect 168725 -173733 168769 -173689
rect 168825 -173733 168869 -173689
rect 168925 -173733 168969 -173689
rect 169025 -173733 169069 -173689
rect 169525 -173733 169569 -173689
rect 169625 -173733 169669 -173689
rect 169725 -173733 169769 -173689
rect 169825 -173733 169869 -173689
rect 169925 -173733 169969 -173689
rect 170025 -173733 170069 -173689
rect 170125 -173733 170169 -173689
rect 170225 -173733 170269 -173689
rect 170325 -173733 170369 -173689
rect 170425 -173733 170469 -173689
rect 170525 -173733 170569 -173689
rect 170625 -173733 170669 -173689
rect 170725 -173733 170769 -173689
rect 170825 -173733 170869 -173689
rect 170925 -173733 170969 -173689
rect 171025 -173733 171069 -173689
rect 171525 -173733 171569 -173689
rect 171625 -173733 171669 -173689
rect 171725 -173733 171769 -173689
rect 171825 -173733 171869 -173689
rect 171925 -173733 171969 -173689
rect 172025 -173733 172069 -173689
rect 172125 -173733 172169 -173689
rect 172225 -173733 172269 -173689
rect 172325 -173733 172369 -173689
rect 172425 -173733 172469 -173689
rect 172525 -173733 172569 -173689
rect 172625 -173733 172669 -173689
rect 172725 -173733 172769 -173689
rect 172825 -173733 172869 -173689
rect 172925 -173733 172969 -173689
rect 173025 -173733 173069 -173689
rect 81627 -173793 81671 -173749
rect 81727 -173793 81771 -173749
rect 81827 -173793 81871 -173749
rect 81927 -173793 81971 -173749
rect 82027 -173793 82071 -173749
rect 82127 -173793 82171 -173749
rect 82227 -173793 82271 -173749
rect 82327 -173793 82371 -173749
rect 82427 -173793 82471 -173749
rect 82527 -173793 82571 -173749
rect 82627 -173793 82671 -173749
rect 82727 -173793 82771 -173749
rect 82827 -173793 82871 -173749
rect 82927 -173793 82971 -173749
rect 83027 -173793 83071 -173749
rect 83127 -173793 83171 -173749
rect 83627 -173793 83671 -173749
rect 83727 -173793 83771 -173749
rect 83827 -173793 83871 -173749
rect 83927 -173793 83971 -173749
rect 84027 -173793 84071 -173749
rect 84127 -173793 84171 -173749
rect 84227 -173793 84271 -173749
rect 84327 -173793 84371 -173749
rect 84427 -173793 84471 -173749
rect 84527 -173793 84571 -173749
rect 84627 -173793 84671 -173749
rect 84727 -173793 84771 -173749
rect 84827 -173793 84871 -173749
rect 84927 -173793 84971 -173749
rect 85027 -173793 85071 -173749
rect 85127 -173793 85171 -173749
rect 85627 -173793 85671 -173749
rect 85727 -173793 85771 -173749
rect 85827 -173793 85871 -173749
rect 85927 -173793 85971 -173749
rect 86027 -173793 86071 -173749
rect 86127 -173793 86171 -173749
rect 86227 -173793 86271 -173749
rect 86327 -173793 86371 -173749
rect 86427 -173793 86471 -173749
rect 86527 -173793 86571 -173749
rect 86627 -173793 86671 -173749
rect 86727 -173793 86771 -173749
rect 86827 -173793 86871 -173749
rect 86927 -173793 86971 -173749
rect 87027 -173793 87071 -173749
rect 87127 -173793 87171 -173749
rect 87627 -173793 87671 -173749
rect 87727 -173793 87771 -173749
rect 87827 -173793 87871 -173749
rect 87927 -173793 87971 -173749
rect 88027 -173793 88071 -173749
rect 88127 -173793 88171 -173749
rect 88227 -173793 88271 -173749
rect 88327 -173793 88371 -173749
rect 88427 -173793 88471 -173749
rect 88527 -173793 88571 -173749
rect 88627 -173793 88671 -173749
rect 88727 -173793 88771 -173749
rect 88827 -173793 88871 -173749
rect 88927 -173793 88971 -173749
rect 89027 -173793 89071 -173749
rect 89127 -173793 89171 -173749
rect 165525 -173833 165569 -173789
rect 165625 -173833 165669 -173789
rect 165725 -173833 165769 -173789
rect 165825 -173833 165869 -173789
rect 165925 -173833 165969 -173789
rect 166025 -173833 166069 -173789
rect 166125 -173833 166169 -173789
rect 166225 -173833 166269 -173789
rect 166325 -173833 166369 -173789
rect 166425 -173833 166469 -173789
rect 166525 -173833 166569 -173789
rect 166625 -173833 166669 -173789
rect 166725 -173833 166769 -173789
rect 166825 -173833 166869 -173789
rect 166925 -173833 166969 -173789
rect 167025 -173833 167069 -173789
rect 167525 -173833 167569 -173789
rect 167625 -173833 167669 -173789
rect 167725 -173833 167769 -173789
rect 167825 -173833 167869 -173789
rect 167925 -173833 167969 -173789
rect 168025 -173833 168069 -173789
rect 168125 -173833 168169 -173789
rect 168225 -173833 168269 -173789
rect 168325 -173833 168369 -173789
rect 168425 -173833 168469 -173789
rect 168525 -173833 168569 -173789
rect 168625 -173833 168669 -173789
rect 168725 -173833 168769 -173789
rect 168825 -173833 168869 -173789
rect 168925 -173833 168969 -173789
rect 169025 -173833 169069 -173789
rect 169525 -173833 169569 -173789
rect 169625 -173833 169669 -173789
rect 169725 -173833 169769 -173789
rect 169825 -173833 169869 -173789
rect 169925 -173833 169969 -173789
rect 170025 -173833 170069 -173789
rect 170125 -173833 170169 -173789
rect 170225 -173833 170269 -173789
rect 170325 -173833 170369 -173789
rect 170425 -173833 170469 -173789
rect 170525 -173833 170569 -173789
rect 170625 -173833 170669 -173789
rect 170725 -173833 170769 -173789
rect 170825 -173833 170869 -173789
rect 170925 -173833 170969 -173789
rect 171025 -173833 171069 -173789
rect 171525 -173833 171569 -173789
rect 171625 -173833 171669 -173789
rect 171725 -173833 171769 -173789
rect 171825 -173833 171869 -173789
rect 171925 -173833 171969 -173789
rect 172025 -173833 172069 -173789
rect 172125 -173833 172169 -173789
rect 172225 -173833 172269 -173789
rect 172325 -173833 172369 -173789
rect 172425 -173833 172469 -173789
rect 172525 -173833 172569 -173789
rect 172625 -173833 172669 -173789
rect 172725 -173833 172769 -173789
rect 172825 -173833 172869 -173789
rect 172925 -173833 172969 -173789
rect 173025 -173833 173069 -173789
rect 81627 -173893 81671 -173849
rect 81727 -173893 81771 -173849
rect 81827 -173893 81871 -173849
rect 81927 -173893 81971 -173849
rect 82027 -173893 82071 -173849
rect 82127 -173893 82171 -173849
rect 82227 -173893 82271 -173849
rect 82327 -173893 82371 -173849
rect 82427 -173893 82471 -173849
rect 82527 -173893 82571 -173849
rect 82627 -173893 82671 -173849
rect 82727 -173893 82771 -173849
rect 82827 -173893 82871 -173849
rect 82927 -173893 82971 -173849
rect 83027 -173893 83071 -173849
rect 83127 -173893 83171 -173849
rect 83627 -173893 83671 -173849
rect 83727 -173893 83771 -173849
rect 83827 -173893 83871 -173849
rect 83927 -173893 83971 -173849
rect 84027 -173893 84071 -173849
rect 84127 -173893 84171 -173849
rect 84227 -173893 84271 -173849
rect 84327 -173893 84371 -173849
rect 84427 -173893 84471 -173849
rect 84527 -173893 84571 -173849
rect 84627 -173893 84671 -173849
rect 84727 -173893 84771 -173849
rect 84827 -173893 84871 -173849
rect 84927 -173893 84971 -173849
rect 85027 -173893 85071 -173849
rect 85127 -173893 85171 -173849
rect 85627 -173893 85671 -173849
rect 85727 -173893 85771 -173849
rect 85827 -173893 85871 -173849
rect 85927 -173893 85971 -173849
rect 86027 -173893 86071 -173849
rect 86127 -173893 86171 -173849
rect 86227 -173893 86271 -173849
rect 86327 -173893 86371 -173849
rect 86427 -173893 86471 -173849
rect 86527 -173893 86571 -173849
rect 86627 -173893 86671 -173849
rect 86727 -173893 86771 -173849
rect 86827 -173893 86871 -173849
rect 86927 -173893 86971 -173849
rect 87027 -173893 87071 -173849
rect 87127 -173893 87171 -173849
rect 87627 -173893 87671 -173849
rect 87727 -173893 87771 -173849
rect 87827 -173893 87871 -173849
rect 87927 -173893 87971 -173849
rect 88027 -173893 88071 -173849
rect 88127 -173893 88171 -173849
rect 88227 -173893 88271 -173849
rect 88327 -173893 88371 -173849
rect 88427 -173893 88471 -173849
rect 88527 -173893 88571 -173849
rect 88627 -173893 88671 -173849
rect 88727 -173893 88771 -173849
rect 88827 -173893 88871 -173849
rect 88927 -173893 88971 -173849
rect 89027 -173893 89071 -173849
rect 89127 -173893 89171 -173849
rect 165525 -173933 165569 -173889
rect 165625 -173933 165669 -173889
rect 165725 -173933 165769 -173889
rect 165825 -173933 165869 -173889
rect 165925 -173933 165969 -173889
rect 166025 -173933 166069 -173889
rect 166125 -173933 166169 -173889
rect 166225 -173933 166269 -173889
rect 166325 -173933 166369 -173889
rect 166425 -173933 166469 -173889
rect 166525 -173933 166569 -173889
rect 166625 -173933 166669 -173889
rect 166725 -173933 166769 -173889
rect 166825 -173933 166869 -173889
rect 166925 -173933 166969 -173889
rect 167025 -173933 167069 -173889
rect 167525 -173933 167569 -173889
rect 167625 -173933 167669 -173889
rect 167725 -173933 167769 -173889
rect 167825 -173933 167869 -173889
rect 167925 -173933 167969 -173889
rect 168025 -173933 168069 -173889
rect 168125 -173933 168169 -173889
rect 168225 -173933 168269 -173889
rect 168325 -173933 168369 -173889
rect 168425 -173933 168469 -173889
rect 168525 -173933 168569 -173889
rect 168625 -173933 168669 -173889
rect 168725 -173933 168769 -173889
rect 168825 -173933 168869 -173889
rect 168925 -173933 168969 -173889
rect 169025 -173933 169069 -173889
rect 169525 -173933 169569 -173889
rect 169625 -173933 169669 -173889
rect 169725 -173933 169769 -173889
rect 169825 -173933 169869 -173889
rect 169925 -173933 169969 -173889
rect 170025 -173933 170069 -173889
rect 170125 -173933 170169 -173889
rect 170225 -173933 170269 -173889
rect 170325 -173933 170369 -173889
rect 170425 -173933 170469 -173889
rect 170525 -173933 170569 -173889
rect 170625 -173933 170669 -173889
rect 170725 -173933 170769 -173889
rect 170825 -173933 170869 -173889
rect 170925 -173933 170969 -173889
rect 171025 -173933 171069 -173889
rect 171525 -173933 171569 -173889
rect 171625 -173933 171669 -173889
rect 171725 -173933 171769 -173889
rect 171825 -173933 171869 -173889
rect 171925 -173933 171969 -173889
rect 172025 -173933 172069 -173889
rect 172125 -173933 172169 -173889
rect 172225 -173933 172269 -173889
rect 172325 -173933 172369 -173889
rect 172425 -173933 172469 -173889
rect 172525 -173933 172569 -173889
rect 172625 -173933 172669 -173889
rect 172725 -173933 172769 -173889
rect 172825 -173933 172869 -173889
rect 172925 -173933 172969 -173889
rect 173025 -173933 173069 -173889
rect 81627 -173993 81671 -173949
rect 81727 -173993 81771 -173949
rect 81827 -173993 81871 -173949
rect 81927 -173993 81971 -173949
rect 82027 -173993 82071 -173949
rect 82127 -173993 82171 -173949
rect 82227 -173993 82271 -173949
rect 82327 -173993 82371 -173949
rect 82427 -173993 82471 -173949
rect 82527 -173993 82571 -173949
rect 82627 -173993 82671 -173949
rect 82727 -173993 82771 -173949
rect 82827 -173993 82871 -173949
rect 82927 -173993 82971 -173949
rect 83027 -173993 83071 -173949
rect 83127 -173993 83171 -173949
rect 83627 -173993 83671 -173949
rect 83727 -173993 83771 -173949
rect 83827 -173993 83871 -173949
rect 83927 -173993 83971 -173949
rect 84027 -173993 84071 -173949
rect 84127 -173993 84171 -173949
rect 84227 -173993 84271 -173949
rect 84327 -173993 84371 -173949
rect 84427 -173993 84471 -173949
rect 84527 -173993 84571 -173949
rect 84627 -173993 84671 -173949
rect 84727 -173993 84771 -173949
rect 84827 -173993 84871 -173949
rect 84927 -173993 84971 -173949
rect 85027 -173993 85071 -173949
rect 85127 -173993 85171 -173949
rect 85627 -173993 85671 -173949
rect 85727 -173993 85771 -173949
rect 85827 -173993 85871 -173949
rect 85927 -173993 85971 -173949
rect 86027 -173993 86071 -173949
rect 86127 -173993 86171 -173949
rect 86227 -173993 86271 -173949
rect 86327 -173993 86371 -173949
rect 86427 -173993 86471 -173949
rect 86527 -173993 86571 -173949
rect 86627 -173993 86671 -173949
rect 86727 -173993 86771 -173949
rect 86827 -173993 86871 -173949
rect 86927 -173993 86971 -173949
rect 87027 -173993 87071 -173949
rect 87127 -173993 87171 -173949
rect 87627 -173993 87671 -173949
rect 87727 -173993 87771 -173949
rect 87827 -173993 87871 -173949
rect 87927 -173993 87971 -173949
rect 88027 -173993 88071 -173949
rect 88127 -173993 88171 -173949
rect 88227 -173993 88271 -173949
rect 88327 -173993 88371 -173949
rect 88427 -173993 88471 -173949
rect 88527 -173993 88571 -173949
rect 88627 -173993 88671 -173949
rect 88727 -173993 88771 -173949
rect 88827 -173993 88871 -173949
rect 88927 -173993 88971 -173949
rect 89027 -173993 89071 -173949
rect 89127 -173993 89171 -173949
rect 165525 -174033 165569 -173989
rect 165625 -174033 165669 -173989
rect 165725 -174033 165769 -173989
rect 165825 -174033 165869 -173989
rect 165925 -174033 165969 -173989
rect 166025 -174033 166069 -173989
rect 166125 -174033 166169 -173989
rect 166225 -174033 166269 -173989
rect 166325 -174033 166369 -173989
rect 166425 -174033 166469 -173989
rect 166525 -174033 166569 -173989
rect 166625 -174033 166669 -173989
rect 166725 -174033 166769 -173989
rect 166825 -174033 166869 -173989
rect 166925 -174033 166969 -173989
rect 167025 -174033 167069 -173989
rect 167525 -174033 167569 -173989
rect 167625 -174033 167669 -173989
rect 167725 -174033 167769 -173989
rect 167825 -174033 167869 -173989
rect 167925 -174033 167969 -173989
rect 168025 -174033 168069 -173989
rect 168125 -174033 168169 -173989
rect 168225 -174033 168269 -173989
rect 168325 -174033 168369 -173989
rect 168425 -174033 168469 -173989
rect 168525 -174033 168569 -173989
rect 168625 -174033 168669 -173989
rect 168725 -174033 168769 -173989
rect 168825 -174033 168869 -173989
rect 168925 -174033 168969 -173989
rect 169025 -174033 169069 -173989
rect 169525 -174033 169569 -173989
rect 169625 -174033 169669 -173989
rect 169725 -174033 169769 -173989
rect 169825 -174033 169869 -173989
rect 169925 -174033 169969 -173989
rect 170025 -174033 170069 -173989
rect 170125 -174033 170169 -173989
rect 170225 -174033 170269 -173989
rect 170325 -174033 170369 -173989
rect 170425 -174033 170469 -173989
rect 170525 -174033 170569 -173989
rect 170625 -174033 170669 -173989
rect 170725 -174033 170769 -173989
rect 170825 -174033 170869 -173989
rect 170925 -174033 170969 -173989
rect 171025 -174033 171069 -173989
rect 171525 -174033 171569 -173989
rect 171625 -174033 171669 -173989
rect 171725 -174033 171769 -173989
rect 171825 -174033 171869 -173989
rect 171925 -174033 171969 -173989
rect 172025 -174033 172069 -173989
rect 172125 -174033 172169 -173989
rect 172225 -174033 172269 -173989
rect 172325 -174033 172369 -173989
rect 172425 -174033 172469 -173989
rect 172525 -174033 172569 -173989
rect 172625 -174033 172669 -173989
rect 172725 -174033 172769 -173989
rect 172825 -174033 172869 -173989
rect 172925 -174033 172969 -173989
rect 173025 -174033 173069 -173989
rect 81627 -174093 81671 -174049
rect 81727 -174093 81771 -174049
rect 81827 -174093 81871 -174049
rect 81927 -174093 81971 -174049
rect 82027 -174093 82071 -174049
rect 82127 -174093 82171 -174049
rect 82227 -174093 82271 -174049
rect 82327 -174093 82371 -174049
rect 82427 -174093 82471 -174049
rect 82527 -174093 82571 -174049
rect 82627 -174093 82671 -174049
rect 82727 -174093 82771 -174049
rect 82827 -174093 82871 -174049
rect 82927 -174093 82971 -174049
rect 83027 -174093 83071 -174049
rect 83127 -174093 83171 -174049
rect 83627 -174093 83671 -174049
rect 83727 -174093 83771 -174049
rect 83827 -174093 83871 -174049
rect 83927 -174093 83971 -174049
rect 84027 -174093 84071 -174049
rect 84127 -174093 84171 -174049
rect 84227 -174093 84271 -174049
rect 84327 -174093 84371 -174049
rect 84427 -174093 84471 -174049
rect 84527 -174093 84571 -174049
rect 84627 -174093 84671 -174049
rect 84727 -174093 84771 -174049
rect 84827 -174093 84871 -174049
rect 84927 -174093 84971 -174049
rect 85027 -174093 85071 -174049
rect 85127 -174093 85171 -174049
rect 85627 -174093 85671 -174049
rect 85727 -174093 85771 -174049
rect 85827 -174093 85871 -174049
rect 85927 -174093 85971 -174049
rect 86027 -174093 86071 -174049
rect 86127 -174093 86171 -174049
rect 86227 -174093 86271 -174049
rect 86327 -174093 86371 -174049
rect 86427 -174093 86471 -174049
rect 86527 -174093 86571 -174049
rect 86627 -174093 86671 -174049
rect 86727 -174093 86771 -174049
rect 86827 -174093 86871 -174049
rect 86927 -174093 86971 -174049
rect 87027 -174093 87071 -174049
rect 87127 -174093 87171 -174049
rect 87627 -174093 87671 -174049
rect 87727 -174093 87771 -174049
rect 87827 -174093 87871 -174049
rect 87927 -174093 87971 -174049
rect 88027 -174093 88071 -174049
rect 88127 -174093 88171 -174049
rect 88227 -174093 88271 -174049
rect 88327 -174093 88371 -174049
rect 88427 -174093 88471 -174049
rect 88527 -174093 88571 -174049
rect 88627 -174093 88671 -174049
rect 88727 -174093 88771 -174049
rect 88827 -174093 88871 -174049
rect 88927 -174093 88971 -174049
rect 89027 -174093 89071 -174049
rect 89127 -174093 89171 -174049
rect 165525 -174133 165569 -174089
rect 165625 -174133 165669 -174089
rect 165725 -174133 165769 -174089
rect 165825 -174133 165869 -174089
rect 165925 -174133 165969 -174089
rect 166025 -174133 166069 -174089
rect 166125 -174133 166169 -174089
rect 166225 -174133 166269 -174089
rect 166325 -174133 166369 -174089
rect 166425 -174133 166469 -174089
rect 166525 -174133 166569 -174089
rect 166625 -174133 166669 -174089
rect 166725 -174133 166769 -174089
rect 166825 -174133 166869 -174089
rect 166925 -174133 166969 -174089
rect 167025 -174133 167069 -174089
rect 167525 -174133 167569 -174089
rect 167625 -174133 167669 -174089
rect 167725 -174133 167769 -174089
rect 167825 -174133 167869 -174089
rect 167925 -174133 167969 -174089
rect 168025 -174133 168069 -174089
rect 168125 -174133 168169 -174089
rect 168225 -174133 168269 -174089
rect 168325 -174133 168369 -174089
rect 168425 -174133 168469 -174089
rect 168525 -174133 168569 -174089
rect 168625 -174133 168669 -174089
rect 168725 -174133 168769 -174089
rect 168825 -174133 168869 -174089
rect 168925 -174133 168969 -174089
rect 169025 -174133 169069 -174089
rect 169525 -174133 169569 -174089
rect 169625 -174133 169669 -174089
rect 169725 -174133 169769 -174089
rect 169825 -174133 169869 -174089
rect 169925 -174133 169969 -174089
rect 170025 -174133 170069 -174089
rect 170125 -174133 170169 -174089
rect 170225 -174133 170269 -174089
rect 170325 -174133 170369 -174089
rect 170425 -174133 170469 -174089
rect 170525 -174133 170569 -174089
rect 170625 -174133 170669 -174089
rect 170725 -174133 170769 -174089
rect 170825 -174133 170869 -174089
rect 170925 -174133 170969 -174089
rect 171025 -174133 171069 -174089
rect 171525 -174133 171569 -174089
rect 171625 -174133 171669 -174089
rect 171725 -174133 171769 -174089
rect 171825 -174133 171869 -174089
rect 171925 -174133 171969 -174089
rect 172025 -174133 172069 -174089
rect 172125 -174133 172169 -174089
rect 172225 -174133 172269 -174089
rect 172325 -174133 172369 -174089
rect 172425 -174133 172469 -174089
rect 172525 -174133 172569 -174089
rect 172625 -174133 172669 -174089
rect 172725 -174133 172769 -174089
rect 172825 -174133 172869 -174089
rect 172925 -174133 172969 -174089
rect 173025 -174133 173069 -174089
rect 81627 -174193 81671 -174149
rect 81727 -174193 81771 -174149
rect 81827 -174193 81871 -174149
rect 81927 -174193 81971 -174149
rect 82027 -174193 82071 -174149
rect 82127 -174193 82171 -174149
rect 82227 -174193 82271 -174149
rect 82327 -174193 82371 -174149
rect 82427 -174193 82471 -174149
rect 82527 -174193 82571 -174149
rect 82627 -174193 82671 -174149
rect 82727 -174193 82771 -174149
rect 82827 -174193 82871 -174149
rect 82927 -174193 82971 -174149
rect 83027 -174193 83071 -174149
rect 83127 -174193 83171 -174149
rect 83627 -174193 83671 -174149
rect 83727 -174193 83771 -174149
rect 83827 -174193 83871 -174149
rect 83927 -174193 83971 -174149
rect 84027 -174193 84071 -174149
rect 84127 -174193 84171 -174149
rect 84227 -174193 84271 -174149
rect 84327 -174193 84371 -174149
rect 84427 -174193 84471 -174149
rect 84527 -174193 84571 -174149
rect 84627 -174193 84671 -174149
rect 84727 -174193 84771 -174149
rect 84827 -174193 84871 -174149
rect 84927 -174193 84971 -174149
rect 85027 -174193 85071 -174149
rect 85127 -174193 85171 -174149
rect 85627 -174193 85671 -174149
rect 85727 -174193 85771 -174149
rect 85827 -174193 85871 -174149
rect 85927 -174193 85971 -174149
rect 86027 -174193 86071 -174149
rect 86127 -174193 86171 -174149
rect 86227 -174193 86271 -174149
rect 86327 -174193 86371 -174149
rect 86427 -174193 86471 -174149
rect 86527 -174193 86571 -174149
rect 86627 -174193 86671 -174149
rect 86727 -174193 86771 -174149
rect 86827 -174193 86871 -174149
rect 86927 -174193 86971 -174149
rect 87027 -174193 87071 -174149
rect 87127 -174193 87171 -174149
rect 87627 -174193 87671 -174149
rect 87727 -174193 87771 -174149
rect 87827 -174193 87871 -174149
rect 87927 -174193 87971 -174149
rect 88027 -174193 88071 -174149
rect 88127 -174193 88171 -174149
rect 88227 -174193 88271 -174149
rect 88327 -174193 88371 -174149
rect 88427 -174193 88471 -174149
rect 88527 -174193 88571 -174149
rect 88627 -174193 88671 -174149
rect 88727 -174193 88771 -174149
rect 88827 -174193 88871 -174149
rect 88927 -174193 88971 -174149
rect 89027 -174193 89071 -174149
rect 89127 -174193 89171 -174149
rect 165525 -174233 165569 -174189
rect 165625 -174233 165669 -174189
rect 165725 -174233 165769 -174189
rect 165825 -174233 165869 -174189
rect 165925 -174233 165969 -174189
rect 166025 -174233 166069 -174189
rect 166125 -174233 166169 -174189
rect 166225 -174233 166269 -174189
rect 166325 -174233 166369 -174189
rect 166425 -174233 166469 -174189
rect 166525 -174233 166569 -174189
rect 166625 -174233 166669 -174189
rect 166725 -174233 166769 -174189
rect 166825 -174233 166869 -174189
rect 166925 -174233 166969 -174189
rect 167025 -174233 167069 -174189
rect 167525 -174233 167569 -174189
rect 167625 -174233 167669 -174189
rect 167725 -174233 167769 -174189
rect 167825 -174233 167869 -174189
rect 167925 -174233 167969 -174189
rect 168025 -174233 168069 -174189
rect 168125 -174233 168169 -174189
rect 168225 -174233 168269 -174189
rect 168325 -174233 168369 -174189
rect 168425 -174233 168469 -174189
rect 168525 -174233 168569 -174189
rect 168625 -174233 168669 -174189
rect 168725 -174233 168769 -174189
rect 168825 -174233 168869 -174189
rect 168925 -174233 168969 -174189
rect 169025 -174233 169069 -174189
rect 169525 -174233 169569 -174189
rect 169625 -174233 169669 -174189
rect 169725 -174233 169769 -174189
rect 169825 -174233 169869 -174189
rect 169925 -174233 169969 -174189
rect 170025 -174233 170069 -174189
rect 170125 -174233 170169 -174189
rect 170225 -174233 170269 -174189
rect 170325 -174233 170369 -174189
rect 170425 -174233 170469 -174189
rect 170525 -174233 170569 -174189
rect 170625 -174233 170669 -174189
rect 170725 -174233 170769 -174189
rect 170825 -174233 170869 -174189
rect 170925 -174233 170969 -174189
rect 171025 -174233 171069 -174189
rect 171525 -174233 171569 -174189
rect 171625 -174233 171669 -174189
rect 171725 -174233 171769 -174189
rect 171825 -174233 171869 -174189
rect 171925 -174233 171969 -174189
rect 172025 -174233 172069 -174189
rect 172125 -174233 172169 -174189
rect 172225 -174233 172269 -174189
rect 172325 -174233 172369 -174189
rect 172425 -174233 172469 -174189
rect 172525 -174233 172569 -174189
rect 172625 -174233 172669 -174189
rect 172725 -174233 172769 -174189
rect 172825 -174233 172869 -174189
rect 172925 -174233 172969 -174189
rect 173025 -174233 173069 -174189
rect 81627 -174293 81671 -174249
rect 81727 -174293 81771 -174249
rect 81827 -174293 81871 -174249
rect 81927 -174293 81971 -174249
rect 82027 -174293 82071 -174249
rect 82127 -174293 82171 -174249
rect 82227 -174293 82271 -174249
rect 82327 -174293 82371 -174249
rect 82427 -174293 82471 -174249
rect 82527 -174293 82571 -174249
rect 82627 -174293 82671 -174249
rect 82727 -174293 82771 -174249
rect 82827 -174293 82871 -174249
rect 82927 -174293 82971 -174249
rect 83027 -174293 83071 -174249
rect 83127 -174293 83171 -174249
rect 83627 -174293 83671 -174249
rect 83727 -174293 83771 -174249
rect 83827 -174293 83871 -174249
rect 83927 -174293 83971 -174249
rect 84027 -174293 84071 -174249
rect 84127 -174293 84171 -174249
rect 84227 -174293 84271 -174249
rect 84327 -174293 84371 -174249
rect 84427 -174293 84471 -174249
rect 84527 -174293 84571 -174249
rect 84627 -174293 84671 -174249
rect 84727 -174293 84771 -174249
rect 84827 -174293 84871 -174249
rect 84927 -174293 84971 -174249
rect 85027 -174293 85071 -174249
rect 85127 -174293 85171 -174249
rect 85627 -174293 85671 -174249
rect 85727 -174293 85771 -174249
rect 85827 -174293 85871 -174249
rect 85927 -174293 85971 -174249
rect 86027 -174293 86071 -174249
rect 86127 -174293 86171 -174249
rect 86227 -174293 86271 -174249
rect 86327 -174293 86371 -174249
rect 86427 -174293 86471 -174249
rect 86527 -174293 86571 -174249
rect 86627 -174293 86671 -174249
rect 86727 -174293 86771 -174249
rect 86827 -174293 86871 -174249
rect 86927 -174293 86971 -174249
rect 87027 -174293 87071 -174249
rect 87127 -174293 87171 -174249
rect 87627 -174293 87671 -174249
rect 87727 -174293 87771 -174249
rect 87827 -174293 87871 -174249
rect 87927 -174293 87971 -174249
rect 88027 -174293 88071 -174249
rect 88127 -174293 88171 -174249
rect 88227 -174293 88271 -174249
rect 88327 -174293 88371 -174249
rect 88427 -174293 88471 -174249
rect 88527 -174293 88571 -174249
rect 88627 -174293 88671 -174249
rect 88727 -174293 88771 -174249
rect 88827 -174293 88871 -174249
rect 88927 -174293 88971 -174249
rect 89027 -174293 89071 -174249
rect 89127 -174293 89171 -174249
rect 165525 -174333 165569 -174289
rect 165625 -174333 165669 -174289
rect 165725 -174333 165769 -174289
rect 165825 -174333 165869 -174289
rect 165925 -174333 165969 -174289
rect 166025 -174333 166069 -174289
rect 166125 -174333 166169 -174289
rect 166225 -174333 166269 -174289
rect 166325 -174333 166369 -174289
rect 166425 -174333 166469 -174289
rect 166525 -174333 166569 -174289
rect 166625 -174333 166669 -174289
rect 166725 -174333 166769 -174289
rect 166825 -174333 166869 -174289
rect 166925 -174333 166969 -174289
rect 167025 -174333 167069 -174289
rect 167525 -174333 167569 -174289
rect 167625 -174333 167669 -174289
rect 167725 -174333 167769 -174289
rect 167825 -174333 167869 -174289
rect 167925 -174333 167969 -174289
rect 168025 -174333 168069 -174289
rect 168125 -174333 168169 -174289
rect 168225 -174333 168269 -174289
rect 168325 -174333 168369 -174289
rect 168425 -174333 168469 -174289
rect 168525 -174333 168569 -174289
rect 168625 -174333 168669 -174289
rect 168725 -174333 168769 -174289
rect 168825 -174333 168869 -174289
rect 168925 -174333 168969 -174289
rect 169025 -174333 169069 -174289
rect 169525 -174333 169569 -174289
rect 169625 -174333 169669 -174289
rect 169725 -174333 169769 -174289
rect 169825 -174333 169869 -174289
rect 169925 -174333 169969 -174289
rect 170025 -174333 170069 -174289
rect 170125 -174333 170169 -174289
rect 170225 -174333 170269 -174289
rect 170325 -174333 170369 -174289
rect 170425 -174333 170469 -174289
rect 170525 -174333 170569 -174289
rect 170625 -174333 170669 -174289
rect 170725 -174333 170769 -174289
rect 170825 -174333 170869 -174289
rect 170925 -174333 170969 -174289
rect 171025 -174333 171069 -174289
rect 171525 -174333 171569 -174289
rect 171625 -174333 171669 -174289
rect 171725 -174333 171769 -174289
rect 171825 -174333 171869 -174289
rect 171925 -174333 171969 -174289
rect 172025 -174333 172069 -174289
rect 172125 -174333 172169 -174289
rect 172225 -174333 172269 -174289
rect 172325 -174333 172369 -174289
rect 172425 -174333 172469 -174289
rect 172525 -174333 172569 -174289
rect 172625 -174333 172669 -174289
rect 172725 -174333 172769 -174289
rect 172825 -174333 172869 -174289
rect 172925 -174333 172969 -174289
rect 173025 -174333 173069 -174289
rect 81627 -174393 81671 -174349
rect 81727 -174393 81771 -174349
rect 81827 -174393 81871 -174349
rect 81927 -174393 81971 -174349
rect 82027 -174393 82071 -174349
rect 82127 -174393 82171 -174349
rect 82227 -174393 82271 -174349
rect 82327 -174393 82371 -174349
rect 82427 -174393 82471 -174349
rect 82527 -174393 82571 -174349
rect 82627 -174393 82671 -174349
rect 82727 -174393 82771 -174349
rect 82827 -174393 82871 -174349
rect 82927 -174393 82971 -174349
rect 83027 -174393 83071 -174349
rect 83127 -174393 83171 -174349
rect 83627 -174393 83671 -174349
rect 83727 -174393 83771 -174349
rect 83827 -174393 83871 -174349
rect 83927 -174393 83971 -174349
rect 84027 -174393 84071 -174349
rect 84127 -174393 84171 -174349
rect 84227 -174393 84271 -174349
rect 84327 -174393 84371 -174349
rect 84427 -174393 84471 -174349
rect 84527 -174393 84571 -174349
rect 84627 -174393 84671 -174349
rect 84727 -174393 84771 -174349
rect 84827 -174393 84871 -174349
rect 84927 -174393 84971 -174349
rect 85027 -174393 85071 -174349
rect 85127 -174393 85171 -174349
rect 85627 -174393 85671 -174349
rect 85727 -174393 85771 -174349
rect 85827 -174393 85871 -174349
rect 85927 -174393 85971 -174349
rect 86027 -174393 86071 -174349
rect 86127 -174393 86171 -174349
rect 86227 -174393 86271 -174349
rect 86327 -174393 86371 -174349
rect 86427 -174393 86471 -174349
rect 86527 -174393 86571 -174349
rect 86627 -174393 86671 -174349
rect 86727 -174393 86771 -174349
rect 86827 -174393 86871 -174349
rect 86927 -174393 86971 -174349
rect 87027 -174393 87071 -174349
rect 87127 -174393 87171 -174349
rect 87627 -174393 87671 -174349
rect 87727 -174393 87771 -174349
rect 87827 -174393 87871 -174349
rect 87927 -174393 87971 -174349
rect 88027 -174393 88071 -174349
rect 88127 -174393 88171 -174349
rect 88227 -174393 88271 -174349
rect 88327 -174393 88371 -174349
rect 88427 -174393 88471 -174349
rect 88527 -174393 88571 -174349
rect 88627 -174393 88671 -174349
rect 88727 -174393 88771 -174349
rect 88827 -174393 88871 -174349
rect 88927 -174393 88971 -174349
rect 89027 -174393 89071 -174349
rect 89127 -174393 89171 -174349
rect 165525 -174433 165569 -174389
rect 165625 -174433 165669 -174389
rect 165725 -174433 165769 -174389
rect 165825 -174433 165869 -174389
rect 165925 -174433 165969 -174389
rect 166025 -174433 166069 -174389
rect 166125 -174433 166169 -174389
rect 166225 -174433 166269 -174389
rect 166325 -174433 166369 -174389
rect 166425 -174433 166469 -174389
rect 166525 -174433 166569 -174389
rect 166625 -174433 166669 -174389
rect 166725 -174433 166769 -174389
rect 166825 -174433 166869 -174389
rect 166925 -174433 166969 -174389
rect 167025 -174433 167069 -174389
rect 167525 -174433 167569 -174389
rect 167625 -174433 167669 -174389
rect 167725 -174433 167769 -174389
rect 167825 -174433 167869 -174389
rect 167925 -174433 167969 -174389
rect 168025 -174433 168069 -174389
rect 168125 -174433 168169 -174389
rect 168225 -174433 168269 -174389
rect 168325 -174433 168369 -174389
rect 168425 -174433 168469 -174389
rect 168525 -174433 168569 -174389
rect 168625 -174433 168669 -174389
rect 168725 -174433 168769 -174389
rect 168825 -174433 168869 -174389
rect 168925 -174433 168969 -174389
rect 169025 -174433 169069 -174389
rect 169525 -174433 169569 -174389
rect 169625 -174433 169669 -174389
rect 169725 -174433 169769 -174389
rect 169825 -174433 169869 -174389
rect 169925 -174433 169969 -174389
rect 170025 -174433 170069 -174389
rect 170125 -174433 170169 -174389
rect 170225 -174433 170269 -174389
rect 170325 -174433 170369 -174389
rect 170425 -174433 170469 -174389
rect 170525 -174433 170569 -174389
rect 170625 -174433 170669 -174389
rect 170725 -174433 170769 -174389
rect 170825 -174433 170869 -174389
rect 170925 -174433 170969 -174389
rect 171025 -174433 171069 -174389
rect 171525 -174433 171569 -174389
rect 171625 -174433 171669 -174389
rect 171725 -174433 171769 -174389
rect 171825 -174433 171869 -174389
rect 171925 -174433 171969 -174389
rect 172025 -174433 172069 -174389
rect 172125 -174433 172169 -174389
rect 172225 -174433 172269 -174389
rect 172325 -174433 172369 -174389
rect 172425 -174433 172469 -174389
rect 172525 -174433 172569 -174389
rect 172625 -174433 172669 -174389
rect 172725 -174433 172769 -174389
rect 172825 -174433 172869 -174389
rect 172925 -174433 172969 -174389
rect 173025 -174433 173069 -174389
rect 81627 -174493 81671 -174449
rect 81727 -174493 81771 -174449
rect 81827 -174493 81871 -174449
rect 81927 -174493 81971 -174449
rect 82027 -174493 82071 -174449
rect 82127 -174493 82171 -174449
rect 82227 -174493 82271 -174449
rect 82327 -174493 82371 -174449
rect 82427 -174493 82471 -174449
rect 82527 -174493 82571 -174449
rect 82627 -174493 82671 -174449
rect 82727 -174493 82771 -174449
rect 82827 -174493 82871 -174449
rect 82927 -174493 82971 -174449
rect 83027 -174493 83071 -174449
rect 83127 -174493 83171 -174449
rect 83627 -174493 83671 -174449
rect 83727 -174493 83771 -174449
rect 83827 -174493 83871 -174449
rect 83927 -174493 83971 -174449
rect 84027 -174493 84071 -174449
rect 84127 -174493 84171 -174449
rect 84227 -174493 84271 -174449
rect 84327 -174493 84371 -174449
rect 84427 -174493 84471 -174449
rect 84527 -174493 84571 -174449
rect 84627 -174493 84671 -174449
rect 84727 -174493 84771 -174449
rect 84827 -174493 84871 -174449
rect 84927 -174493 84971 -174449
rect 85027 -174493 85071 -174449
rect 85127 -174493 85171 -174449
rect 85627 -174493 85671 -174449
rect 85727 -174493 85771 -174449
rect 85827 -174493 85871 -174449
rect 85927 -174493 85971 -174449
rect 86027 -174493 86071 -174449
rect 86127 -174493 86171 -174449
rect 86227 -174493 86271 -174449
rect 86327 -174493 86371 -174449
rect 86427 -174493 86471 -174449
rect 86527 -174493 86571 -174449
rect 86627 -174493 86671 -174449
rect 86727 -174493 86771 -174449
rect 86827 -174493 86871 -174449
rect 86927 -174493 86971 -174449
rect 87027 -174493 87071 -174449
rect 87127 -174493 87171 -174449
rect 87627 -174493 87671 -174449
rect 87727 -174493 87771 -174449
rect 87827 -174493 87871 -174449
rect 87927 -174493 87971 -174449
rect 88027 -174493 88071 -174449
rect 88127 -174493 88171 -174449
rect 88227 -174493 88271 -174449
rect 88327 -174493 88371 -174449
rect 88427 -174493 88471 -174449
rect 88527 -174493 88571 -174449
rect 88627 -174493 88671 -174449
rect 88727 -174493 88771 -174449
rect 88827 -174493 88871 -174449
rect 88927 -174493 88971 -174449
rect 89027 -174493 89071 -174449
rect 89127 -174493 89171 -174449
rect 165525 -174533 165569 -174489
rect 165625 -174533 165669 -174489
rect 165725 -174533 165769 -174489
rect 165825 -174533 165869 -174489
rect 165925 -174533 165969 -174489
rect 166025 -174533 166069 -174489
rect 166125 -174533 166169 -174489
rect 166225 -174533 166269 -174489
rect 166325 -174533 166369 -174489
rect 166425 -174533 166469 -174489
rect 166525 -174533 166569 -174489
rect 166625 -174533 166669 -174489
rect 166725 -174533 166769 -174489
rect 166825 -174533 166869 -174489
rect 166925 -174533 166969 -174489
rect 167025 -174533 167069 -174489
rect 167525 -174533 167569 -174489
rect 167625 -174533 167669 -174489
rect 167725 -174533 167769 -174489
rect 167825 -174533 167869 -174489
rect 167925 -174533 167969 -174489
rect 168025 -174533 168069 -174489
rect 168125 -174533 168169 -174489
rect 168225 -174533 168269 -174489
rect 168325 -174533 168369 -174489
rect 168425 -174533 168469 -174489
rect 168525 -174533 168569 -174489
rect 168625 -174533 168669 -174489
rect 168725 -174533 168769 -174489
rect 168825 -174533 168869 -174489
rect 168925 -174533 168969 -174489
rect 169025 -174533 169069 -174489
rect 169525 -174533 169569 -174489
rect 169625 -174533 169669 -174489
rect 169725 -174533 169769 -174489
rect 169825 -174533 169869 -174489
rect 169925 -174533 169969 -174489
rect 170025 -174533 170069 -174489
rect 170125 -174533 170169 -174489
rect 170225 -174533 170269 -174489
rect 170325 -174533 170369 -174489
rect 170425 -174533 170469 -174489
rect 170525 -174533 170569 -174489
rect 170625 -174533 170669 -174489
rect 170725 -174533 170769 -174489
rect 170825 -174533 170869 -174489
rect 170925 -174533 170969 -174489
rect 171025 -174533 171069 -174489
rect 171525 -174533 171569 -174489
rect 171625 -174533 171669 -174489
rect 171725 -174533 171769 -174489
rect 171825 -174533 171869 -174489
rect 171925 -174533 171969 -174489
rect 172025 -174533 172069 -174489
rect 172125 -174533 172169 -174489
rect 172225 -174533 172269 -174489
rect 172325 -174533 172369 -174489
rect 172425 -174533 172469 -174489
rect 172525 -174533 172569 -174489
rect 172625 -174533 172669 -174489
rect 172725 -174533 172769 -174489
rect 172825 -174533 172869 -174489
rect 172925 -174533 172969 -174489
rect 173025 -174533 173069 -174489
rect 81627 -174593 81671 -174549
rect 81727 -174593 81771 -174549
rect 81827 -174593 81871 -174549
rect 81927 -174593 81971 -174549
rect 82027 -174593 82071 -174549
rect 82127 -174593 82171 -174549
rect 82227 -174593 82271 -174549
rect 82327 -174593 82371 -174549
rect 82427 -174593 82471 -174549
rect 82527 -174593 82571 -174549
rect 82627 -174593 82671 -174549
rect 82727 -174593 82771 -174549
rect 82827 -174593 82871 -174549
rect 82927 -174593 82971 -174549
rect 83027 -174593 83071 -174549
rect 83127 -174593 83171 -174549
rect 83627 -174593 83671 -174549
rect 83727 -174593 83771 -174549
rect 83827 -174593 83871 -174549
rect 83927 -174593 83971 -174549
rect 84027 -174593 84071 -174549
rect 84127 -174593 84171 -174549
rect 84227 -174593 84271 -174549
rect 84327 -174593 84371 -174549
rect 84427 -174593 84471 -174549
rect 84527 -174593 84571 -174549
rect 84627 -174593 84671 -174549
rect 84727 -174593 84771 -174549
rect 84827 -174593 84871 -174549
rect 84927 -174593 84971 -174549
rect 85027 -174593 85071 -174549
rect 85127 -174593 85171 -174549
rect 85627 -174593 85671 -174549
rect 85727 -174593 85771 -174549
rect 85827 -174593 85871 -174549
rect 85927 -174593 85971 -174549
rect 86027 -174593 86071 -174549
rect 86127 -174593 86171 -174549
rect 86227 -174593 86271 -174549
rect 86327 -174593 86371 -174549
rect 86427 -174593 86471 -174549
rect 86527 -174593 86571 -174549
rect 86627 -174593 86671 -174549
rect 86727 -174593 86771 -174549
rect 86827 -174593 86871 -174549
rect 86927 -174593 86971 -174549
rect 87027 -174593 87071 -174549
rect 87127 -174593 87171 -174549
rect 87627 -174593 87671 -174549
rect 87727 -174593 87771 -174549
rect 87827 -174593 87871 -174549
rect 87927 -174593 87971 -174549
rect 88027 -174593 88071 -174549
rect 88127 -174593 88171 -174549
rect 88227 -174593 88271 -174549
rect 88327 -174593 88371 -174549
rect 88427 -174593 88471 -174549
rect 88527 -174593 88571 -174549
rect 88627 -174593 88671 -174549
rect 88727 -174593 88771 -174549
rect 88827 -174593 88871 -174549
rect 88927 -174593 88971 -174549
rect 89027 -174593 89071 -174549
rect 89127 -174593 89171 -174549
<< metal2 >>
rect 178461 9674 181332 10636
rect 178461 9144 179458 9674
rect 180057 9144 181332 9674
rect -105430 3555 -18301 5041
rect -105430 3511 -27407 3555
rect -27363 3511 -27307 3555
rect -27263 3511 -27207 3555
rect -27163 3511 -27107 3555
rect -27063 3511 -27007 3555
rect -26963 3511 -26907 3555
rect -26863 3511 -26807 3555
rect -26763 3511 -26707 3555
rect -26663 3511 -26607 3555
rect -26563 3511 -26507 3555
rect -26463 3511 -26407 3555
rect -26363 3511 -26307 3555
rect -26263 3511 -26207 3555
rect -26163 3511 -26107 3555
rect -26063 3511 -26007 3555
rect -25963 3511 -25907 3555
rect -25863 3511 -25407 3555
rect -25363 3511 -25307 3555
rect -25263 3511 -25207 3555
rect -25163 3511 -25107 3555
rect -25063 3511 -25007 3555
rect -24963 3511 -24907 3555
rect -24863 3511 -24807 3555
rect -24763 3511 -24707 3555
rect -24663 3511 -24607 3555
rect -24563 3511 -24507 3555
rect -24463 3511 -24407 3555
rect -24363 3511 -24307 3555
rect -24263 3511 -24207 3555
rect -24163 3511 -24107 3555
rect -24063 3511 -24007 3555
rect -23963 3511 -23907 3555
rect -23863 3511 -23407 3555
rect -23363 3511 -23307 3555
rect -23263 3511 -23207 3555
rect -23163 3511 -23107 3555
rect -23063 3511 -23007 3555
rect -22963 3511 -22907 3555
rect -22863 3511 -22807 3555
rect -22763 3511 -22707 3555
rect -22663 3511 -22607 3555
rect -22563 3511 -22507 3555
rect -22463 3511 -22407 3555
rect -22363 3511 -22307 3555
rect -22263 3511 -22207 3555
rect -22163 3511 -22107 3555
rect -22063 3511 -22007 3555
rect -21963 3511 -21907 3555
rect -21863 3511 -21407 3555
rect -21363 3511 -21307 3555
rect -21263 3511 -21207 3555
rect -21163 3511 -21107 3555
rect -21063 3511 -21007 3555
rect -20963 3511 -20907 3555
rect -20863 3511 -20807 3555
rect -20763 3511 -20707 3555
rect -20663 3511 -20607 3555
rect -20563 3511 -20507 3555
rect -20463 3511 -20407 3555
rect -20363 3511 -20307 3555
rect -20263 3511 -20207 3555
rect -20163 3511 -20107 3555
rect -20063 3511 -20007 3555
rect -19963 3511 -19907 3555
rect -19863 3511 -18301 3555
rect -105430 3455 -18301 3511
rect -105430 3411 -27407 3455
rect -27363 3411 -27307 3455
rect -27263 3411 -27207 3455
rect -27163 3411 -27107 3455
rect -27063 3411 -27007 3455
rect -26963 3411 -26907 3455
rect -26863 3411 -26807 3455
rect -26763 3411 -26707 3455
rect -26663 3411 -26607 3455
rect -26563 3411 -26507 3455
rect -26463 3411 -26407 3455
rect -26363 3411 -26307 3455
rect -26263 3411 -26207 3455
rect -26163 3411 -26107 3455
rect -26063 3411 -26007 3455
rect -25963 3411 -25907 3455
rect -25863 3411 -25407 3455
rect -25363 3411 -25307 3455
rect -25263 3411 -25207 3455
rect -25163 3411 -25107 3455
rect -25063 3411 -25007 3455
rect -24963 3411 -24907 3455
rect -24863 3411 -24807 3455
rect -24763 3411 -24707 3455
rect -24663 3411 -24607 3455
rect -24563 3411 -24507 3455
rect -24463 3411 -24407 3455
rect -24363 3411 -24307 3455
rect -24263 3411 -24207 3455
rect -24163 3411 -24107 3455
rect -24063 3411 -24007 3455
rect -23963 3411 -23907 3455
rect -23863 3411 -23407 3455
rect -23363 3411 -23307 3455
rect -23263 3411 -23207 3455
rect -23163 3411 -23107 3455
rect -23063 3411 -23007 3455
rect -22963 3411 -22907 3455
rect -22863 3411 -22807 3455
rect -22763 3411 -22707 3455
rect -22663 3411 -22607 3455
rect -22563 3411 -22507 3455
rect -22463 3411 -22407 3455
rect -22363 3411 -22307 3455
rect -22263 3411 -22207 3455
rect -22163 3411 -22107 3455
rect -22063 3411 -22007 3455
rect -21963 3411 -21907 3455
rect -21863 3411 -21407 3455
rect -21363 3411 -21307 3455
rect -21263 3411 -21207 3455
rect -21163 3411 -21107 3455
rect -21063 3411 -21007 3455
rect -20963 3411 -20907 3455
rect -20863 3411 -20807 3455
rect -20763 3411 -20707 3455
rect -20663 3411 -20607 3455
rect -20563 3411 -20507 3455
rect -20463 3411 -20407 3455
rect -20363 3411 -20307 3455
rect -20263 3411 -20207 3455
rect -20163 3411 -20107 3455
rect -20063 3411 -20007 3455
rect -19963 3411 -19907 3455
rect -19863 3411 -18301 3455
rect -105430 3355 -18301 3411
rect -105430 3311 -27407 3355
rect -27363 3311 -27307 3355
rect -27263 3311 -27207 3355
rect -27163 3311 -27107 3355
rect -27063 3311 -27007 3355
rect -26963 3311 -26907 3355
rect -26863 3311 -26807 3355
rect -26763 3311 -26707 3355
rect -26663 3311 -26607 3355
rect -26563 3311 -26507 3355
rect -26463 3311 -26407 3355
rect -26363 3311 -26307 3355
rect -26263 3311 -26207 3355
rect -26163 3311 -26107 3355
rect -26063 3311 -26007 3355
rect -25963 3311 -25907 3355
rect -25863 3311 -25407 3355
rect -25363 3311 -25307 3355
rect -25263 3311 -25207 3355
rect -25163 3311 -25107 3355
rect -25063 3311 -25007 3355
rect -24963 3311 -24907 3355
rect -24863 3311 -24807 3355
rect -24763 3311 -24707 3355
rect -24663 3311 -24607 3355
rect -24563 3311 -24507 3355
rect -24463 3311 -24407 3355
rect -24363 3311 -24307 3355
rect -24263 3311 -24207 3355
rect -24163 3311 -24107 3355
rect -24063 3311 -24007 3355
rect -23963 3311 -23907 3355
rect -23863 3311 -23407 3355
rect -23363 3311 -23307 3355
rect -23263 3311 -23207 3355
rect -23163 3311 -23107 3355
rect -23063 3311 -23007 3355
rect -22963 3311 -22907 3355
rect -22863 3311 -22807 3355
rect -22763 3311 -22707 3355
rect -22663 3311 -22607 3355
rect -22563 3311 -22507 3355
rect -22463 3311 -22407 3355
rect -22363 3311 -22307 3355
rect -22263 3311 -22207 3355
rect -22163 3311 -22107 3355
rect -22063 3311 -22007 3355
rect -21963 3311 -21907 3355
rect -21863 3311 -21407 3355
rect -21363 3311 -21307 3355
rect -21263 3311 -21207 3355
rect -21163 3311 -21107 3355
rect -21063 3311 -21007 3355
rect -20963 3311 -20907 3355
rect -20863 3311 -20807 3355
rect -20763 3311 -20707 3355
rect -20663 3311 -20607 3355
rect -20563 3311 -20507 3355
rect -20463 3311 -20407 3355
rect -20363 3311 -20307 3355
rect -20263 3311 -20207 3355
rect -20163 3311 -20107 3355
rect -20063 3311 -20007 3355
rect -19963 3311 -19907 3355
rect -19863 3311 -18301 3355
rect -105430 3255 -18301 3311
rect -105430 3211 -27407 3255
rect -27363 3211 -27307 3255
rect -27263 3211 -27207 3255
rect -27163 3211 -27107 3255
rect -27063 3211 -27007 3255
rect -26963 3211 -26907 3255
rect -26863 3211 -26807 3255
rect -26763 3211 -26707 3255
rect -26663 3211 -26607 3255
rect -26563 3211 -26507 3255
rect -26463 3211 -26407 3255
rect -26363 3211 -26307 3255
rect -26263 3211 -26207 3255
rect -26163 3211 -26107 3255
rect -26063 3211 -26007 3255
rect -25963 3211 -25907 3255
rect -25863 3211 -25407 3255
rect -25363 3211 -25307 3255
rect -25263 3211 -25207 3255
rect -25163 3211 -25107 3255
rect -25063 3211 -25007 3255
rect -24963 3211 -24907 3255
rect -24863 3211 -24807 3255
rect -24763 3211 -24707 3255
rect -24663 3211 -24607 3255
rect -24563 3211 -24507 3255
rect -24463 3211 -24407 3255
rect -24363 3211 -24307 3255
rect -24263 3211 -24207 3255
rect -24163 3211 -24107 3255
rect -24063 3211 -24007 3255
rect -23963 3211 -23907 3255
rect -23863 3211 -23407 3255
rect -23363 3211 -23307 3255
rect -23263 3211 -23207 3255
rect -23163 3211 -23107 3255
rect -23063 3211 -23007 3255
rect -22963 3211 -22907 3255
rect -22863 3211 -22807 3255
rect -22763 3211 -22707 3255
rect -22663 3211 -22607 3255
rect -22563 3211 -22507 3255
rect -22463 3211 -22407 3255
rect -22363 3211 -22307 3255
rect -22263 3211 -22207 3255
rect -22163 3211 -22107 3255
rect -22063 3211 -22007 3255
rect -21963 3211 -21907 3255
rect -21863 3211 -21407 3255
rect -21363 3211 -21307 3255
rect -21263 3211 -21207 3255
rect -21163 3211 -21107 3255
rect -21063 3211 -21007 3255
rect -20963 3211 -20907 3255
rect -20863 3211 -20807 3255
rect -20763 3211 -20707 3255
rect -20663 3211 -20607 3255
rect -20563 3211 -20507 3255
rect -20463 3211 -20407 3255
rect -20363 3211 -20307 3255
rect -20263 3211 -20207 3255
rect -20163 3211 -20107 3255
rect -20063 3211 -20007 3255
rect -19963 3211 -19907 3255
rect -19863 3211 -18301 3255
rect -105430 3155 -18301 3211
rect -105430 3111 -27407 3155
rect -27363 3111 -27307 3155
rect -27263 3111 -27207 3155
rect -27163 3111 -27107 3155
rect -27063 3111 -27007 3155
rect -26963 3111 -26907 3155
rect -26863 3111 -26807 3155
rect -26763 3111 -26707 3155
rect -26663 3111 -26607 3155
rect -26563 3111 -26507 3155
rect -26463 3111 -26407 3155
rect -26363 3111 -26307 3155
rect -26263 3111 -26207 3155
rect -26163 3111 -26107 3155
rect -26063 3111 -26007 3155
rect -25963 3111 -25907 3155
rect -25863 3111 -25407 3155
rect -25363 3111 -25307 3155
rect -25263 3111 -25207 3155
rect -25163 3111 -25107 3155
rect -25063 3111 -25007 3155
rect -24963 3111 -24907 3155
rect -24863 3111 -24807 3155
rect -24763 3111 -24707 3155
rect -24663 3111 -24607 3155
rect -24563 3111 -24507 3155
rect -24463 3111 -24407 3155
rect -24363 3111 -24307 3155
rect -24263 3111 -24207 3155
rect -24163 3111 -24107 3155
rect -24063 3111 -24007 3155
rect -23963 3111 -23907 3155
rect -23863 3111 -23407 3155
rect -23363 3111 -23307 3155
rect -23263 3111 -23207 3155
rect -23163 3111 -23107 3155
rect -23063 3111 -23007 3155
rect -22963 3111 -22907 3155
rect -22863 3111 -22807 3155
rect -22763 3111 -22707 3155
rect -22663 3111 -22607 3155
rect -22563 3111 -22507 3155
rect -22463 3111 -22407 3155
rect -22363 3111 -22307 3155
rect -22263 3111 -22207 3155
rect -22163 3111 -22107 3155
rect -22063 3111 -22007 3155
rect -21963 3111 -21907 3155
rect -21863 3111 -21407 3155
rect -21363 3111 -21307 3155
rect -21263 3111 -21207 3155
rect -21163 3111 -21107 3155
rect -21063 3111 -21007 3155
rect -20963 3111 -20907 3155
rect -20863 3111 -20807 3155
rect -20763 3111 -20707 3155
rect -20663 3111 -20607 3155
rect -20563 3111 -20507 3155
rect -20463 3111 -20407 3155
rect -20363 3111 -20307 3155
rect -20263 3111 -20207 3155
rect -20163 3111 -20107 3155
rect -20063 3111 -20007 3155
rect -19963 3111 -19907 3155
rect -19863 3111 -18301 3155
rect -105430 3055 -18301 3111
rect -105430 3011 -27407 3055
rect -27363 3011 -27307 3055
rect -27263 3011 -27207 3055
rect -27163 3011 -27107 3055
rect -27063 3011 -27007 3055
rect -26963 3011 -26907 3055
rect -26863 3011 -26807 3055
rect -26763 3011 -26707 3055
rect -26663 3011 -26607 3055
rect -26563 3011 -26507 3055
rect -26463 3011 -26407 3055
rect -26363 3011 -26307 3055
rect -26263 3011 -26207 3055
rect -26163 3011 -26107 3055
rect -26063 3011 -26007 3055
rect -25963 3011 -25907 3055
rect -25863 3011 -25407 3055
rect -25363 3011 -25307 3055
rect -25263 3011 -25207 3055
rect -25163 3011 -25107 3055
rect -25063 3011 -25007 3055
rect -24963 3011 -24907 3055
rect -24863 3011 -24807 3055
rect -24763 3011 -24707 3055
rect -24663 3011 -24607 3055
rect -24563 3011 -24507 3055
rect -24463 3011 -24407 3055
rect -24363 3011 -24307 3055
rect -24263 3011 -24207 3055
rect -24163 3011 -24107 3055
rect -24063 3011 -24007 3055
rect -23963 3011 -23907 3055
rect -23863 3011 -23407 3055
rect -23363 3011 -23307 3055
rect -23263 3011 -23207 3055
rect -23163 3011 -23107 3055
rect -23063 3011 -23007 3055
rect -22963 3011 -22907 3055
rect -22863 3011 -22807 3055
rect -22763 3011 -22707 3055
rect -22663 3011 -22607 3055
rect -22563 3011 -22507 3055
rect -22463 3011 -22407 3055
rect -22363 3011 -22307 3055
rect -22263 3011 -22207 3055
rect -22163 3011 -22107 3055
rect -22063 3011 -22007 3055
rect -21963 3011 -21907 3055
rect -21863 3011 -21407 3055
rect -21363 3011 -21307 3055
rect -21263 3011 -21207 3055
rect -21163 3011 -21107 3055
rect -21063 3011 -21007 3055
rect -20963 3011 -20907 3055
rect -20863 3011 -20807 3055
rect -20763 3011 -20707 3055
rect -20663 3011 -20607 3055
rect -20563 3011 -20507 3055
rect -20463 3011 -20407 3055
rect -20363 3011 -20307 3055
rect -20263 3011 -20207 3055
rect -20163 3011 -20107 3055
rect -20063 3011 -20007 3055
rect -19963 3011 -19907 3055
rect -19863 3011 -18301 3055
rect -105430 2955 -18301 3011
rect -105430 2911 -27407 2955
rect -27363 2911 -27307 2955
rect -27263 2911 -27207 2955
rect -27163 2911 -27107 2955
rect -27063 2911 -27007 2955
rect -26963 2911 -26907 2955
rect -26863 2911 -26807 2955
rect -26763 2911 -26707 2955
rect -26663 2911 -26607 2955
rect -26563 2911 -26507 2955
rect -26463 2911 -26407 2955
rect -26363 2911 -26307 2955
rect -26263 2911 -26207 2955
rect -26163 2911 -26107 2955
rect -26063 2911 -26007 2955
rect -25963 2911 -25907 2955
rect -25863 2911 -25407 2955
rect -25363 2911 -25307 2955
rect -25263 2911 -25207 2955
rect -25163 2911 -25107 2955
rect -25063 2911 -25007 2955
rect -24963 2911 -24907 2955
rect -24863 2911 -24807 2955
rect -24763 2911 -24707 2955
rect -24663 2911 -24607 2955
rect -24563 2911 -24507 2955
rect -24463 2911 -24407 2955
rect -24363 2911 -24307 2955
rect -24263 2911 -24207 2955
rect -24163 2911 -24107 2955
rect -24063 2911 -24007 2955
rect -23963 2911 -23907 2955
rect -23863 2911 -23407 2955
rect -23363 2911 -23307 2955
rect -23263 2911 -23207 2955
rect -23163 2911 -23107 2955
rect -23063 2911 -23007 2955
rect -22963 2911 -22907 2955
rect -22863 2911 -22807 2955
rect -22763 2911 -22707 2955
rect -22663 2911 -22607 2955
rect -22563 2911 -22507 2955
rect -22463 2911 -22407 2955
rect -22363 2911 -22307 2955
rect -22263 2911 -22207 2955
rect -22163 2911 -22107 2955
rect -22063 2911 -22007 2955
rect -21963 2911 -21907 2955
rect -21863 2911 -21407 2955
rect -21363 2911 -21307 2955
rect -21263 2911 -21207 2955
rect -21163 2911 -21107 2955
rect -21063 2911 -21007 2955
rect -20963 2911 -20907 2955
rect -20863 2911 -20807 2955
rect -20763 2911 -20707 2955
rect -20663 2911 -20607 2955
rect -20563 2911 -20507 2955
rect -20463 2911 -20407 2955
rect -20363 2911 -20307 2955
rect -20263 2911 -20207 2955
rect -20163 2911 -20107 2955
rect -20063 2911 -20007 2955
rect -19963 2911 -19907 2955
rect -19863 2911 -18301 2955
rect -105430 2855 -18301 2911
rect -105430 2811 -27407 2855
rect -27363 2811 -27307 2855
rect -27263 2811 -27207 2855
rect -27163 2811 -27107 2855
rect -27063 2811 -27007 2855
rect -26963 2811 -26907 2855
rect -26863 2811 -26807 2855
rect -26763 2811 -26707 2855
rect -26663 2811 -26607 2855
rect -26563 2811 -26507 2855
rect -26463 2811 -26407 2855
rect -26363 2811 -26307 2855
rect -26263 2811 -26207 2855
rect -26163 2811 -26107 2855
rect -26063 2811 -26007 2855
rect -25963 2811 -25907 2855
rect -25863 2811 -25407 2855
rect -25363 2811 -25307 2855
rect -25263 2811 -25207 2855
rect -25163 2811 -25107 2855
rect -25063 2811 -25007 2855
rect -24963 2811 -24907 2855
rect -24863 2811 -24807 2855
rect -24763 2811 -24707 2855
rect -24663 2811 -24607 2855
rect -24563 2811 -24507 2855
rect -24463 2811 -24407 2855
rect -24363 2811 -24307 2855
rect -24263 2811 -24207 2855
rect -24163 2811 -24107 2855
rect -24063 2811 -24007 2855
rect -23963 2811 -23907 2855
rect -23863 2811 -23407 2855
rect -23363 2811 -23307 2855
rect -23263 2811 -23207 2855
rect -23163 2811 -23107 2855
rect -23063 2811 -23007 2855
rect -22963 2811 -22907 2855
rect -22863 2811 -22807 2855
rect -22763 2811 -22707 2855
rect -22663 2811 -22607 2855
rect -22563 2811 -22507 2855
rect -22463 2811 -22407 2855
rect -22363 2811 -22307 2855
rect -22263 2811 -22207 2855
rect -22163 2811 -22107 2855
rect -22063 2811 -22007 2855
rect -21963 2811 -21907 2855
rect -21863 2811 -21407 2855
rect -21363 2811 -21307 2855
rect -21263 2811 -21207 2855
rect -21163 2811 -21107 2855
rect -21063 2811 -21007 2855
rect -20963 2811 -20907 2855
rect -20863 2811 -20807 2855
rect -20763 2811 -20707 2855
rect -20663 2811 -20607 2855
rect -20563 2811 -20507 2855
rect -20463 2811 -20407 2855
rect -20363 2811 -20307 2855
rect -20263 2811 -20207 2855
rect -20163 2811 -20107 2855
rect -20063 2811 -20007 2855
rect -19963 2811 -19907 2855
rect -19863 2811 -18301 2855
rect -105430 2755 -18301 2811
rect -105430 2711 -27407 2755
rect -27363 2711 -27307 2755
rect -27263 2711 -27207 2755
rect -27163 2711 -27107 2755
rect -27063 2711 -27007 2755
rect -26963 2711 -26907 2755
rect -26863 2711 -26807 2755
rect -26763 2711 -26707 2755
rect -26663 2711 -26607 2755
rect -26563 2711 -26507 2755
rect -26463 2711 -26407 2755
rect -26363 2711 -26307 2755
rect -26263 2711 -26207 2755
rect -26163 2711 -26107 2755
rect -26063 2711 -26007 2755
rect -25963 2711 -25907 2755
rect -25863 2711 -25407 2755
rect -25363 2711 -25307 2755
rect -25263 2711 -25207 2755
rect -25163 2711 -25107 2755
rect -25063 2711 -25007 2755
rect -24963 2711 -24907 2755
rect -24863 2711 -24807 2755
rect -24763 2711 -24707 2755
rect -24663 2711 -24607 2755
rect -24563 2711 -24507 2755
rect -24463 2711 -24407 2755
rect -24363 2711 -24307 2755
rect -24263 2711 -24207 2755
rect -24163 2711 -24107 2755
rect -24063 2711 -24007 2755
rect -23963 2711 -23907 2755
rect -23863 2711 -23407 2755
rect -23363 2711 -23307 2755
rect -23263 2711 -23207 2755
rect -23163 2711 -23107 2755
rect -23063 2711 -23007 2755
rect -22963 2711 -22907 2755
rect -22863 2711 -22807 2755
rect -22763 2711 -22707 2755
rect -22663 2711 -22607 2755
rect -22563 2711 -22507 2755
rect -22463 2711 -22407 2755
rect -22363 2711 -22307 2755
rect -22263 2711 -22207 2755
rect -22163 2711 -22107 2755
rect -22063 2711 -22007 2755
rect -21963 2711 -21907 2755
rect -21863 2711 -21407 2755
rect -21363 2711 -21307 2755
rect -21263 2711 -21207 2755
rect -21163 2711 -21107 2755
rect -21063 2711 -21007 2755
rect -20963 2711 -20907 2755
rect -20863 2711 -20807 2755
rect -20763 2711 -20707 2755
rect -20663 2711 -20607 2755
rect -20563 2711 -20507 2755
rect -20463 2711 -20407 2755
rect -20363 2711 -20307 2755
rect -20263 2711 -20207 2755
rect -20163 2711 -20107 2755
rect -20063 2711 -20007 2755
rect -19963 2711 -19907 2755
rect -19863 2711 -18301 2755
rect -105430 2655 -18301 2711
rect -105430 2611 -27407 2655
rect -27363 2611 -27307 2655
rect -27263 2611 -27207 2655
rect -27163 2611 -27107 2655
rect -27063 2611 -27007 2655
rect -26963 2611 -26907 2655
rect -26863 2611 -26807 2655
rect -26763 2611 -26707 2655
rect -26663 2611 -26607 2655
rect -26563 2611 -26507 2655
rect -26463 2611 -26407 2655
rect -26363 2611 -26307 2655
rect -26263 2611 -26207 2655
rect -26163 2611 -26107 2655
rect -26063 2611 -26007 2655
rect -25963 2611 -25907 2655
rect -25863 2611 -25407 2655
rect -25363 2611 -25307 2655
rect -25263 2611 -25207 2655
rect -25163 2611 -25107 2655
rect -25063 2611 -25007 2655
rect -24963 2611 -24907 2655
rect -24863 2611 -24807 2655
rect -24763 2611 -24707 2655
rect -24663 2611 -24607 2655
rect -24563 2611 -24507 2655
rect -24463 2611 -24407 2655
rect -24363 2611 -24307 2655
rect -24263 2611 -24207 2655
rect -24163 2611 -24107 2655
rect -24063 2611 -24007 2655
rect -23963 2611 -23907 2655
rect -23863 2611 -23407 2655
rect -23363 2611 -23307 2655
rect -23263 2611 -23207 2655
rect -23163 2611 -23107 2655
rect -23063 2611 -23007 2655
rect -22963 2611 -22907 2655
rect -22863 2611 -22807 2655
rect -22763 2611 -22707 2655
rect -22663 2611 -22607 2655
rect -22563 2611 -22507 2655
rect -22463 2611 -22407 2655
rect -22363 2611 -22307 2655
rect -22263 2611 -22207 2655
rect -22163 2611 -22107 2655
rect -22063 2611 -22007 2655
rect -21963 2611 -21907 2655
rect -21863 2611 -21407 2655
rect -21363 2611 -21307 2655
rect -21263 2611 -21207 2655
rect -21163 2611 -21107 2655
rect -21063 2611 -21007 2655
rect -20963 2611 -20907 2655
rect -20863 2611 -20807 2655
rect -20763 2611 -20707 2655
rect -20663 2611 -20607 2655
rect -20563 2611 -20507 2655
rect -20463 2611 -20407 2655
rect -20363 2611 -20307 2655
rect -20263 2611 -20207 2655
rect -20163 2611 -20107 2655
rect -20063 2611 -20007 2655
rect -19963 2611 -19907 2655
rect -19863 2611 -18301 2655
rect -105430 2555 -18301 2611
rect -105430 2511 -27407 2555
rect -27363 2511 -27307 2555
rect -27263 2511 -27207 2555
rect -27163 2511 -27107 2555
rect -27063 2511 -27007 2555
rect -26963 2511 -26907 2555
rect -26863 2511 -26807 2555
rect -26763 2511 -26707 2555
rect -26663 2511 -26607 2555
rect -26563 2511 -26507 2555
rect -26463 2511 -26407 2555
rect -26363 2511 -26307 2555
rect -26263 2511 -26207 2555
rect -26163 2511 -26107 2555
rect -26063 2511 -26007 2555
rect -25963 2511 -25907 2555
rect -25863 2511 -25407 2555
rect -25363 2511 -25307 2555
rect -25263 2511 -25207 2555
rect -25163 2511 -25107 2555
rect -25063 2511 -25007 2555
rect -24963 2511 -24907 2555
rect -24863 2511 -24807 2555
rect -24763 2511 -24707 2555
rect -24663 2511 -24607 2555
rect -24563 2511 -24507 2555
rect -24463 2511 -24407 2555
rect -24363 2511 -24307 2555
rect -24263 2511 -24207 2555
rect -24163 2511 -24107 2555
rect -24063 2511 -24007 2555
rect -23963 2511 -23907 2555
rect -23863 2511 -23407 2555
rect -23363 2511 -23307 2555
rect -23263 2511 -23207 2555
rect -23163 2511 -23107 2555
rect -23063 2511 -23007 2555
rect -22963 2511 -22907 2555
rect -22863 2511 -22807 2555
rect -22763 2511 -22707 2555
rect -22663 2511 -22607 2555
rect -22563 2511 -22507 2555
rect -22463 2511 -22407 2555
rect -22363 2511 -22307 2555
rect -22263 2511 -22207 2555
rect -22163 2511 -22107 2555
rect -22063 2511 -22007 2555
rect -21963 2511 -21907 2555
rect -21863 2511 -21407 2555
rect -21363 2511 -21307 2555
rect -21263 2511 -21207 2555
rect -21163 2511 -21107 2555
rect -21063 2511 -21007 2555
rect -20963 2511 -20907 2555
rect -20863 2511 -20807 2555
rect -20763 2511 -20707 2555
rect -20663 2511 -20607 2555
rect -20563 2511 -20507 2555
rect -20463 2511 -20407 2555
rect -20363 2511 -20307 2555
rect -20263 2511 -20207 2555
rect -20163 2511 -20107 2555
rect -20063 2511 -20007 2555
rect -19963 2511 -19907 2555
rect -19863 2511 -18301 2555
rect -105430 2455 -18301 2511
rect -105430 2411 -27407 2455
rect -27363 2411 -27307 2455
rect -27263 2411 -27207 2455
rect -27163 2411 -27107 2455
rect -27063 2411 -27007 2455
rect -26963 2411 -26907 2455
rect -26863 2411 -26807 2455
rect -26763 2411 -26707 2455
rect -26663 2411 -26607 2455
rect -26563 2411 -26507 2455
rect -26463 2411 -26407 2455
rect -26363 2411 -26307 2455
rect -26263 2411 -26207 2455
rect -26163 2411 -26107 2455
rect -26063 2411 -26007 2455
rect -25963 2411 -25907 2455
rect -25863 2411 -25407 2455
rect -25363 2411 -25307 2455
rect -25263 2411 -25207 2455
rect -25163 2411 -25107 2455
rect -25063 2411 -25007 2455
rect -24963 2411 -24907 2455
rect -24863 2411 -24807 2455
rect -24763 2411 -24707 2455
rect -24663 2411 -24607 2455
rect -24563 2411 -24507 2455
rect -24463 2411 -24407 2455
rect -24363 2411 -24307 2455
rect -24263 2411 -24207 2455
rect -24163 2411 -24107 2455
rect -24063 2411 -24007 2455
rect -23963 2411 -23907 2455
rect -23863 2411 -23407 2455
rect -23363 2411 -23307 2455
rect -23263 2411 -23207 2455
rect -23163 2411 -23107 2455
rect -23063 2411 -23007 2455
rect -22963 2411 -22907 2455
rect -22863 2411 -22807 2455
rect -22763 2411 -22707 2455
rect -22663 2411 -22607 2455
rect -22563 2411 -22507 2455
rect -22463 2411 -22407 2455
rect -22363 2411 -22307 2455
rect -22263 2411 -22207 2455
rect -22163 2411 -22107 2455
rect -22063 2411 -22007 2455
rect -21963 2411 -21907 2455
rect -21863 2411 -21407 2455
rect -21363 2411 -21307 2455
rect -21263 2411 -21207 2455
rect -21163 2411 -21107 2455
rect -21063 2411 -21007 2455
rect -20963 2411 -20907 2455
rect -20863 2411 -20807 2455
rect -20763 2411 -20707 2455
rect -20663 2411 -20607 2455
rect -20563 2411 -20507 2455
rect -20463 2411 -20407 2455
rect -20363 2411 -20307 2455
rect -20263 2411 -20207 2455
rect -20163 2411 -20107 2455
rect -20063 2411 -20007 2455
rect -19963 2411 -19907 2455
rect -19863 2411 -18301 2455
rect -105430 2355 -18301 2411
rect -105430 2311 -27407 2355
rect -27363 2311 -27307 2355
rect -27263 2311 -27207 2355
rect -27163 2311 -27107 2355
rect -27063 2311 -27007 2355
rect -26963 2311 -26907 2355
rect -26863 2311 -26807 2355
rect -26763 2311 -26707 2355
rect -26663 2311 -26607 2355
rect -26563 2311 -26507 2355
rect -26463 2311 -26407 2355
rect -26363 2311 -26307 2355
rect -26263 2311 -26207 2355
rect -26163 2311 -26107 2355
rect -26063 2311 -26007 2355
rect -25963 2311 -25907 2355
rect -25863 2311 -25407 2355
rect -25363 2311 -25307 2355
rect -25263 2311 -25207 2355
rect -25163 2311 -25107 2355
rect -25063 2311 -25007 2355
rect -24963 2311 -24907 2355
rect -24863 2311 -24807 2355
rect -24763 2311 -24707 2355
rect -24663 2311 -24607 2355
rect -24563 2311 -24507 2355
rect -24463 2311 -24407 2355
rect -24363 2311 -24307 2355
rect -24263 2311 -24207 2355
rect -24163 2311 -24107 2355
rect -24063 2311 -24007 2355
rect -23963 2311 -23907 2355
rect -23863 2311 -23407 2355
rect -23363 2311 -23307 2355
rect -23263 2311 -23207 2355
rect -23163 2311 -23107 2355
rect -23063 2311 -23007 2355
rect -22963 2311 -22907 2355
rect -22863 2311 -22807 2355
rect -22763 2311 -22707 2355
rect -22663 2311 -22607 2355
rect -22563 2311 -22507 2355
rect -22463 2311 -22407 2355
rect -22363 2311 -22307 2355
rect -22263 2311 -22207 2355
rect -22163 2311 -22107 2355
rect -22063 2311 -22007 2355
rect -21963 2311 -21907 2355
rect -21863 2311 -21407 2355
rect -21363 2311 -21307 2355
rect -21263 2311 -21207 2355
rect -21163 2311 -21107 2355
rect -21063 2311 -21007 2355
rect -20963 2311 -20907 2355
rect -20863 2311 -20807 2355
rect -20763 2311 -20707 2355
rect -20663 2311 -20607 2355
rect -20563 2311 -20507 2355
rect -20463 2311 -20407 2355
rect -20363 2311 -20307 2355
rect -20263 2311 -20207 2355
rect -20163 2311 -20107 2355
rect -20063 2311 -20007 2355
rect -19963 2311 -19907 2355
rect -19863 2311 -18301 2355
rect -105430 2255 -18301 2311
rect -105430 2211 -27407 2255
rect -27363 2211 -27307 2255
rect -27263 2211 -27207 2255
rect -27163 2211 -27107 2255
rect -27063 2211 -27007 2255
rect -26963 2211 -26907 2255
rect -26863 2211 -26807 2255
rect -26763 2211 -26707 2255
rect -26663 2211 -26607 2255
rect -26563 2211 -26507 2255
rect -26463 2211 -26407 2255
rect -26363 2211 -26307 2255
rect -26263 2211 -26207 2255
rect -26163 2211 -26107 2255
rect -26063 2211 -26007 2255
rect -25963 2211 -25907 2255
rect -25863 2211 -25407 2255
rect -25363 2211 -25307 2255
rect -25263 2211 -25207 2255
rect -25163 2211 -25107 2255
rect -25063 2211 -25007 2255
rect -24963 2211 -24907 2255
rect -24863 2211 -24807 2255
rect -24763 2211 -24707 2255
rect -24663 2211 -24607 2255
rect -24563 2211 -24507 2255
rect -24463 2211 -24407 2255
rect -24363 2211 -24307 2255
rect -24263 2211 -24207 2255
rect -24163 2211 -24107 2255
rect -24063 2211 -24007 2255
rect -23963 2211 -23907 2255
rect -23863 2211 -23407 2255
rect -23363 2211 -23307 2255
rect -23263 2211 -23207 2255
rect -23163 2211 -23107 2255
rect -23063 2211 -23007 2255
rect -22963 2211 -22907 2255
rect -22863 2211 -22807 2255
rect -22763 2211 -22707 2255
rect -22663 2211 -22607 2255
rect -22563 2211 -22507 2255
rect -22463 2211 -22407 2255
rect -22363 2211 -22307 2255
rect -22263 2211 -22207 2255
rect -22163 2211 -22107 2255
rect -22063 2211 -22007 2255
rect -21963 2211 -21907 2255
rect -21863 2211 -21407 2255
rect -21363 2211 -21307 2255
rect -21263 2211 -21207 2255
rect -21163 2211 -21107 2255
rect -21063 2211 -21007 2255
rect -20963 2211 -20907 2255
rect -20863 2211 -20807 2255
rect -20763 2211 -20707 2255
rect -20663 2211 -20607 2255
rect -20563 2211 -20507 2255
rect -20463 2211 -20407 2255
rect -20363 2211 -20307 2255
rect -20263 2211 -20207 2255
rect -20163 2211 -20107 2255
rect -20063 2211 -20007 2255
rect -19963 2211 -19907 2255
rect -19863 2211 -18301 2255
rect -105430 2155 -18301 2211
rect -105430 2111 -27407 2155
rect -27363 2111 -27307 2155
rect -27263 2111 -27207 2155
rect -27163 2111 -27107 2155
rect -27063 2111 -27007 2155
rect -26963 2111 -26907 2155
rect -26863 2111 -26807 2155
rect -26763 2111 -26707 2155
rect -26663 2111 -26607 2155
rect -26563 2111 -26507 2155
rect -26463 2111 -26407 2155
rect -26363 2111 -26307 2155
rect -26263 2111 -26207 2155
rect -26163 2111 -26107 2155
rect -26063 2111 -26007 2155
rect -25963 2111 -25907 2155
rect -25863 2111 -25407 2155
rect -25363 2111 -25307 2155
rect -25263 2111 -25207 2155
rect -25163 2111 -25107 2155
rect -25063 2111 -25007 2155
rect -24963 2111 -24907 2155
rect -24863 2111 -24807 2155
rect -24763 2111 -24707 2155
rect -24663 2111 -24607 2155
rect -24563 2111 -24507 2155
rect -24463 2111 -24407 2155
rect -24363 2111 -24307 2155
rect -24263 2111 -24207 2155
rect -24163 2111 -24107 2155
rect -24063 2111 -24007 2155
rect -23963 2111 -23907 2155
rect -23863 2111 -23407 2155
rect -23363 2111 -23307 2155
rect -23263 2111 -23207 2155
rect -23163 2111 -23107 2155
rect -23063 2111 -23007 2155
rect -22963 2111 -22907 2155
rect -22863 2111 -22807 2155
rect -22763 2111 -22707 2155
rect -22663 2111 -22607 2155
rect -22563 2111 -22507 2155
rect -22463 2111 -22407 2155
rect -22363 2111 -22307 2155
rect -22263 2111 -22207 2155
rect -22163 2111 -22107 2155
rect -22063 2111 -22007 2155
rect -21963 2111 -21907 2155
rect -21863 2111 -21407 2155
rect -21363 2111 -21307 2155
rect -21263 2111 -21207 2155
rect -21163 2111 -21107 2155
rect -21063 2111 -21007 2155
rect -20963 2111 -20907 2155
rect -20863 2111 -20807 2155
rect -20763 2111 -20707 2155
rect -20663 2111 -20607 2155
rect -20563 2111 -20507 2155
rect -20463 2111 -20407 2155
rect -20363 2111 -20307 2155
rect -20263 2111 -20207 2155
rect -20163 2111 -20107 2155
rect -20063 2111 -20007 2155
rect -19963 2111 -19907 2155
rect -19863 2111 -18301 2155
rect -105430 2055 -18301 2111
rect -105430 2011 -27407 2055
rect -27363 2011 -27307 2055
rect -27263 2011 -27207 2055
rect -27163 2011 -27107 2055
rect -27063 2011 -27007 2055
rect -26963 2011 -26907 2055
rect -26863 2011 -26807 2055
rect -26763 2011 -26707 2055
rect -26663 2011 -26607 2055
rect -26563 2011 -26507 2055
rect -26463 2011 -26407 2055
rect -26363 2011 -26307 2055
rect -26263 2011 -26207 2055
rect -26163 2011 -26107 2055
rect -26063 2011 -26007 2055
rect -25963 2011 -25907 2055
rect -25863 2011 -25407 2055
rect -25363 2011 -25307 2055
rect -25263 2011 -25207 2055
rect -25163 2011 -25107 2055
rect -25063 2011 -25007 2055
rect -24963 2011 -24907 2055
rect -24863 2011 -24807 2055
rect -24763 2011 -24707 2055
rect -24663 2011 -24607 2055
rect -24563 2011 -24507 2055
rect -24463 2011 -24407 2055
rect -24363 2011 -24307 2055
rect -24263 2011 -24207 2055
rect -24163 2011 -24107 2055
rect -24063 2011 -24007 2055
rect -23963 2011 -23907 2055
rect -23863 2011 -23407 2055
rect -23363 2011 -23307 2055
rect -23263 2011 -23207 2055
rect -23163 2011 -23107 2055
rect -23063 2011 -23007 2055
rect -22963 2011 -22907 2055
rect -22863 2011 -22807 2055
rect -22763 2011 -22707 2055
rect -22663 2011 -22607 2055
rect -22563 2011 -22507 2055
rect -22463 2011 -22407 2055
rect -22363 2011 -22307 2055
rect -22263 2011 -22207 2055
rect -22163 2011 -22107 2055
rect -22063 2011 -22007 2055
rect -21963 2011 -21907 2055
rect -21863 2011 -21407 2055
rect -21363 2011 -21307 2055
rect -21263 2011 -21207 2055
rect -21163 2011 -21107 2055
rect -21063 2011 -21007 2055
rect -20963 2011 -20907 2055
rect -20863 2011 -20807 2055
rect -20763 2011 -20707 2055
rect -20663 2011 -20607 2055
rect -20563 2011 -20507 2055
rect -20463 2011 -20407 2055
rect -20363 2011 -20307 2055
rect -20263 2011 -20207 2055
rect -20163 2011 -20107 2055
rect -20063 2011 -20007 2055
rect -19963 2011 -19907 2055
rect -19863 2011 -18301 2055
rect -105430 379 -18301 2011
rect 120915 3016 124714 3140
rect 120915 2353 122315 3016
rect 123454 2353 124714 3016
rect -105430 -135314 -96269 379
rect -16721 -2958 118225 -2106
rect 120915 -2958 124714 2353
rect -16721 -4472 125401 -2958
rect -16721 -4804 118225 -4472
rect 120915 -4668 124714 -4472
rect -16721 -7154 -3437 -4804
rect -16721 -7374 -12772 -7154
rect -12552 -7374 -12302 -7154
rect -12082 -7374 -11832 -7154
rect -11612 -7374 -11362 -7154
rect -11142 -7374 -10892 -7154
rect -10672 -7374 -10422 -7154
rect -10202 -7374 -9952 -7154
rect -9732 -7374 -9482 -7154
rect -9262 -7374 -9012 -7154
rect -8792 -7374 -8542 -7154
rect -8322 -7374 -8072 -7154
rect -7852 -7374 -7602 -7154
rect -7382 -7374 -7132 -7154
rect -6912 -7374 -6662 -7154
rect -6442 -7374 -3437 -7154
rect -16721 -8175 -3437 -7374
rect 7194 -9756 18364 -7194
rect 7194 -9800 9195 -9756
rect 9239 -9800 9295 -9756
rect 9339 -9800 9395 -9756
rect 9439 -9800 9495 -9756
rect 9539 -9800 9595 -9756
rect 9639 -9800 9695 -9756
rect 9739 -9800 9795 -9756
rect 9839 -9800 9895 -9756
rect 9939 -9800 9995 -9756
rect 10039 -9800 10095 -9756
rect 10139 -9800 10195 -9756
rect 10239 -9800 10295 -9756
rect 10339 -9800 10395 -9756
rect 10439 -9800 10495 -9756
rect 10539 -9800 10595 -9756
rect 10639 -9800 10695 -9756
rect 10739 -9800 11195 -9756
rect 11239 -9800 11295 -9756
rect 11339 -9800 11395 -9756
rect 11439 -9800 11495 -9756
rect 11539 -9800 11595 -9756
rect 11639 -9800 11695 -9756
rect 11739 -9800 11795 -9756
rect 11839 -9800 11895 -9756
rect 11939 -9800 11995 -9756
rect 12039 -9800 12095 -9756
rect 12139 -9800 12195 -9756
rect 12239 -9800 12295 -9756
rect 12339 -9800 12395 -9756
rect 12439 -9800 12495 -9756
rect 12539 -9800 12595 -9756
rect 12639 -9800 12695 -9756
rect 12739 -9800 13195 -9756
rect 13239 -9800 13295 -9756
rect 13339 -9800 13395 -9756
rect 13439 -9800 13495 -9756
rect 13539 -9800 13595 -9756
rect 13639 -9800 13695 -9756
rect 13739 -9800 13795 -9756
rect 13839 -9800 13895 -9756
rect 13939 -9800 13995 -9756
rect 14039 -9800 14095 -9756
rect 14139 -9800 14195 -9756
rect 14239 -9800 14295 -9756
rect 14339 -9800 14395 -9756
rect 14439 -9800 14495 -9756
rect 14539 -9800 14595 -9756
rect 14639 -9800 14695 -9756
rect 14739 -9800 15195 -9756
rect 15239 -9800 15295 -9756
rect 15339 -9800 15395 -9756
rect 15439 -9800 15495 -9756
rect 15539 -9800 15595 -9756
rect 15639 -9800 15695 -9756
rect 15739 -9800 15795 -9756
rect 15839 -9800 15895 -9756
rect 15939 -9800 15995 -9756
rect 16039 -9800 16095 -9756
rect 16139 -9800 16195 -9756
rect 16239 -9800 16295 -9756
rect 16339 -9800 16395 -9756
rect 16439 -9800 16495 -9756
rect 16539 -9800 16595 -9756
rect 16639 -9800 16695 -9756
rect 16739 -9800 18364 -9756
rect 7194 -9856 18364 -9800
rect 7194 -9900 9195 -9856
rect 9239 -9900 9295 -9856
rect 9339 -9900 9395 -9856
rect 9439 -9900 9495 -9856
rect 9539 -9900 9595 -9856
rect 9639 -9900 9695 -9856
rect 9739 -9900 9795 -9856
rect 9839 -9900 9895 -9856
rect 9939 -9900 9995 -9856
rect 10039 -9900 10095 -9856
rect 10139 -9900 10195 -9856
rect 10239 -9900 10295 -9856
rect 10339 -9900 10395 -9856
rect 10439 -9900 10495 -9856
rect 10539 -9900 10595 -9856
rect 10639 -9900 10695 -9856
rect 10739 -9900 11195 -9856
rect 11239 -9900 11295 -9856
rect 11339 -9900 11395 -9856
rect 11439 -9900 11495 -9856
rect 11539 -9900 11595 -9856
rect 11639 -9900 11695 -9856
rect 11739 -9900 11795 -9856
rect 11839 -9900 11895 -9856
rect 11939 -9900 11995 -9856
rect 12039 -9900 12095 -9856
rect 12139 -9900 12195 -9856
rect 12239 -9900 12295 -9856
rect 12339 -9900 12395 -9856
rect 12439 -9900 12495 -9856
rect 12539 -9900 12595 -9856
rect 12639 -9900 12695 -9856
rect 12739 -9900 13195 -9856
rect 13239 -9900 13295 -9856
rect 13339 -9900 13395 -9856
rect 13439 -9900 13495 -9856
rect 13539 -9900 13595 -9856
rect 13639 -9900 13695 -9856
rect 13739 -9900 13795 -9856
rect 13839 -9900 13895 -9856
rect 13939 -9900 13995 -9856
rect 14039 -9900 14095 -9856
rect 14139 -9900 14195 -9856
rect 14239 -9900 14295 -9856
rect 14339 -9900 14395 -9856
rect 14439 -9900 14495 -9856
rect 14539 -9900 14595 -9856
rect 14639 -9900 14695 -9856
rect 14739 -9900 15195 -9856
rect 15239 -9900 15295 -9856
rect 15339 -9900 15395 -9856
rect 15439 -9900 15495 -9856
rect 15539 -9900 15595 -9856
rect 15639 -9900 15695 -9856
rect 15739 -9900 15795 -9856
rect 15839 -9900 15895 -9856
rect 15939 -9900 15995 -9856
rect 16039 -9900 16095 -9856
rect 16139 -9900 16195 -9856
rect 16239 -9900 16295 -9856
rect 16339 -9900 16395 -9856
rect 16439 -9900 16495 -9856
rect 16539 -9900 16595 -9856
rect 16639 -9900 16695 -9856
rect 16739 -9900 18364 -9856
rect 7194 -9956 18364 -9900
rect 7194 -10000 9195 -9956
rect 9239 -10000 9295 -9956
rect 9339 -10000 9395 -9956
rect 9439 -10000 9495 -9956
rect 9539 -10000 9595 -9956
rect 9639 -10000 9695 -9956
rect 9739 -10000 9795 -9956
rect 9839 -10000 9895 -9956
rect 9939 -10000 9995 -9956
rect 10039 -10000 10095 -9956
rect 10139 -10000 10195 -9956
rect 10239 -10000 10295 -9956
rect 10339 -10000 10395 -9956
rect 10439 -10000 10495 -9956
rect 10539 -10000 10595 -9956
rect 10639 -10000 10695 -9956
rect 10739 -10000 11195 -9956
rect 11239 -10000 11295 -9956
rect 11339 -10000 11395 -9956
rect 11439 -10000 11495 -9956
rect 11539 -10000 11595 -9956
rect 11639 -10000 11695 -9956
rect 11739 -10000 11795 -9956
rect 11839 -10000 11895 -9956
rect 11939 -10000 11995 -9956
rect 12039 -10000 12095 -9956
rect 12139 -10000 12195 -9956
rect 12239 -10000 12295 -9956
rect 12339 -10000 12395 -9956
rect 12439 -10000 12495 -9956
rect 12539 -10000 12595 -9956
rect 12639 -10000 12695 -9956
rect 12739 -10000 13195 -9956
rect 13239 -10000 13295 -9956
rect 13339 -10000 13395 -9956
rect 13439 -10000 13495 -9956
rect 13539 -10000 13595 -9956
rect 13639 -10000 13695 -9956
rect 13739 -10000 13795 -9956
rect 13839 -10000 13895 -9956
rect 13939 -10000 13995 -9956
rect 14039 -10000 14095 -9956
rect 14139 -10000 14195 -9956
rect 14239 -10000 14295 -9956
rect 14339 -10000 14395 -9956
rect 14439 -10000 14495 -9956
rect 14539 -10000 14595 -9956
rect 14639 -10000 14695 -9956
rect 14739 -10000 15195 -9956
rect 15239 -10000 15295 -9956
rect 15339 -10000 15395 -9956
rect 15439 -10000 15495 -9956
rect 15539 -10000 15595 -9956
rect 15639 -10000 15695 -9956
rect 15739 -10000 15795 -9956
rect 15839 -10000 15895 -9956
rect 15939 -10000 15995 -9956
rect 16039 -10000 16095 -9956
rect 16139 -10000 16195 -9956
rect 16239 -10000 16295 -9956
rect 16339 -10000 16395 -9956
rect 16439 -10000 16495 -9956
rect 16539 -10000 16595 -9956
rect 16639 -10000 16695 -9956
rect 16739 -10000 18364 -9956
rect 7194 -10056 18364 -10000
rect 7194 -10100 9195 -10056
rect 9239 -10100 9295 -10056
rect 9339 -10100 9395 -10056
rect 9439 -10100 9495 -10056
rect 9539 -10100 9595 -10056
rect 9639 -10100 9695 -10056
rect 9739 -10100 9795 -10056
rect 9839 -10100 9895 -10056
rect 9939 -10100 9995 -10056
rect 10039 -10100 10095 -10056
rect 10139 -10100 10195 -10056
rect 10239 -10100 10295 -10056
rect 10339 -10100 10395 -10056
rect 10439 -10100 10495 -10056
rect 10539 -10100 10595 -10056
rect 10639 -10100 10695 -10056
rect 10739 -10100 11195 -10056
rect 11239 -10100 11295 -10056
rect 11339 -10100 11395 -10056
rect 11439 -10100 11495 -10056
rect 11539 -10100 11595 -10056
rect 11639 -10100 11695 -10056
rect 11739 -10100 11795 -10056
rect 11839 -10100 11895 -10056
rect 11939 -10100 11995 -10056
rect 12039 -10100 12095 -10056
rect 12139 -10100 12195 -10056
rect 12239 -10100 12295 -10056
rect 12339 -10100 12395 -10056
rect 12439 -10100 12495 -10056
rect 12539 -10100 12595 -10056
rect 12639 -10100 12695 -10056
rect 12739 -10100 13195 -10056
rect 13239 -10100 13295 -10056
rect 13339 -10100 13395 -10056
rect 13439 -10100 13495 -10056
rect 13539 -10100 13595 -10056
rect 13639 -10100 13695 -10056
rect 13739 -10100 13795 -10056
rect 13839 -10100 13895 -10056
rect 13939 -10100 13995 -10056
rect 14039 -10100 14095 -10056
rect 14139 -10100 14195 -10056
rect 14239 -10100 14295 -10056
rect 14339 -10100 14395 -10056
rect 14439 -10100 14495 -10056
rect 14539 -10100 14595 -10056
rect 14639 -10100 14695 -10056
rect 14739 -10100 15195 -10056
rect 15239 -10100 15295 -10056
rect 15339 -10100 15395 -10056
rect 15439 -10100 15495 -10056
rect 15539 -10100 15595 -10056
rect 15639 -10100 15695 -10056
rect 15739 -10100 15795 -10056
rect 15839 -10100 15895 -10056
rect 15939 -10100 15995 -10056
rect 16039 -10100 16095 -10056
rect 16139 -10100 16195 -10056
rect 16239 -10100 16295 -10056
rect 16339 -10100 16395 -10056
rect 16439 -10100 16495 -10056
rect 16539 -10100 16595 -10056
rect 16639 -10100 16695 -10056
rect 16739 -10100 18364 -10056
rect 7194 -10156 18364 -10100
rect 7194 -10200 9195 -10156
rect 9239 -10200 9295 -10156
rect 9339 -10200 9395 -10156
rect 9439 -10200 9495 -10156
rect 9539 -10200 9595 -10156
rect 9639 -10200 9695 -10156
rect 9739 -10200 9795 -10156
rect 9839 -10200 9895 -10156
rect 9939 -10200 9995 -10156
rect 10039 -10200 10095 -10156
rect 10139 -10200 10195 -10156
rect 10239 -10200 10295 -10156
rect 10339 -10200 10395 -10156
rect 10439 -10200 10495 -10156
rect 10539 -10200 10595 -10156
rect 10639 -10200 10695 -10156
rect 10739 -10200 11195 -10156
rect 11239 -10200 11295 -10156
rect 11339 -10200 11395 -10156
rect 11439 -10200 11495 -10156
rect 11539 -10200 11595 -10156
rect 11639 -10200 11695 -10156
rect 11739 -10200 11795 -10156
rect 11839 -10200 11895 -10156
rect 11939 -10200 11995 -10156
rect 12039 -10200 12095 -10156
rect 12139 -10200 12195 -10156
rect 12239 -10200 12295 -10156
rect 12339 -10200 12395 -10156
rect 12439 -10200 12495 -10156
rect 12539 -10200 12595 -10156
rect 12639 -10200 12695 -10156
rect 12739 -10200 13195 -10156
rect 13239 -10200 13295 -10156
rect 13339 -10200 13395 -10156
rect 13439 -10200 13495 -10156
rect 13539 -10200 13595 -10156
rect 13639 -10200 13695 -10156
rect 13739 -10200 13795 -10156
rect 13839 -10200 13895 -10156
rect 13939 -10200 13995 -10156
rect 14039 -10200 14095 -10156
rect 14139 -10200 14195 -10156
rect 14239 -10200 14295 -10156
rect 14339 -10200 14395 -10156
rect 14439 -10200 14495 -10156
rect 14539 -10200 14595 -10156
rect 14639 -10200 14695 -10156
rect 14739 -10200 15195 -10156
rect 15239 -10200 15295 -10156
rect 15339 -10200 15395 -10156
rect 15439 -10200 15495 -10156
rect 15539 -10200 15595 -10156
rect 15639 -10200 15695 -10156
rect 15739 -10200 15795 -10156
rect 15839 -10200 15895 -10156
rect 15939 -10200 15995 -10156
rect 16039 -10200 16095 -10156
rect 16139 -10200 16195 -10156
rect 16239 -10200 16295 -10156
rect 16339 -10200 16395 -10156
rect 16439 -10200 16495 -10156
rect 16539 -10200 16595 -10156
rect 16639 -10200 16695 -10156
rect 16739 -10200 18364 -10156
rect 7194 -10256 18364 -10200
rect 7194 -10300 9195 -10256
rect 9239 -10300 9295 -10256
rect 9339 -10300 9395 -10256
rect 9439 -10300 9495 -10256
rect 9539 -10300 9595 -10256
rect 9639 -10300 9695 -10256
rect 9739 -10300 9795 -10256
rect 9839 -10300 9895 -10256
rect 9939 -10300 9995 -10256
rect 10039 -10300 10095 -10256
rect 10139 -10300 10195 -10256
rect 10239 -10300 10295 -10256
rect 10339 -10300 10395 -10256
rect 10439 -10300 10495 -10256
rect 10539 -10300 10595 -10256
rect 10639 -10300 10695 -10256
rect 10739 -10300 11195 -10256
rect 11239 -10300 11295 -10256
rect 11339 -10300 11395 -10256
rect 11439 -10300 11495 -10256
rect 11539 -10300 11595 -10256
rect 11639 -10300 11695 -10256
rect 11739 -10300 11795 -10256
rect 11839 -10300 11895 -10256
rect 11939 -10300 11995 -10256
rect 12039 -10300 12095 -10256
rect 12139 -10300 12195 -10256
rect 12239 -10300 12295 -10256
rect 12339 -10300 12395 -10256
rect 12439 -10300 12495 -10256
rect 12539 -10300 12595 -10256
rect 12639 -10300 12695 -10256
rect 12739 -10300 13195 -10256
rect 13239 -10300 13295 -10256
rect 13339 -10300 13395 -10256
rect 13439 -10300 13495 -10256
rect 13539 -10300 13595 -10256
rect 13639 -10300 13695 -10256
rect 13739 -10300 13795 -10256
rect 13839 -10300 13895 -10256
rect 13939 -10300 13995 -10256
rect 14039 -10300 14095 -10256
rect 14139 -10300 14195 -10256
rect 14239 -10300 14295 -10256
rect 14339 -10300 14395 -10256
rect 14439 -10300 14495 -10256
rect 14539 -10300 14595 -10256
rect 14639 -10300 14695 -10256
rect 14739 -10300 15195 -10256
rect 15239 -10300 15295 -10256
rect 15339 -10300 15395 -10256
rect 15439 -10300 15495 -10256
rect 15539 -10300 15595 -10256
rect 15639 -10300 15695 -10256
rect 15739 -10300 15795 -10256
rect 15839 -10300 15895 -10256
rect 15939 -10300 15995 -10256
rect 16039 -10300 16095 -10256
rect 16139 -10300 16195 -10256
rect 16239 -10300 16295 -10256
rect 16339 -10300 16395 -10256
rect 16439 -10300 16495 -10256
rect 16539 -10300 16595 -10256
rect 16639 -10300 16695 -10256
rect 16739 -10300 18364 -10256
rect 7194 -10356 18364 -10300
rect 7194 -10400 9195 -10356
rect 9239 -10400 9295 -10356
rect 9339 -10400 9395 -10356
rect 9439 -10400 9495 -10356
rect 9539 -10400 9595 -10356
rect 9639 -10400 9695 -10356
rect 9739 -10400 9795 -10356
rect 9839 -10400 9895 -10356
rect 9939 -10400 9995 -10356
rect 10039 -10400 10095 -10356
rect 10139 -10400 10195 -10356
rect 10239 -10400 10295 -10356
rect 10339 -10400 10395 -10356
rect 10439 -10400 10495 -10356
rect 10539 -10400 10595 -10356
rect 10639 -10400 10695 -10356
rect 10739 -10400 11195 -10356
rect 11239 -10400 11295 -10356
rect 11339 -10400 11395 -10356
rect 11439 -10400 11495 -10356
rect 11539 -10400 11595 -10356
rect 11639 -10400 11695 -10356
rect 11739 -10400 11795 -10356
rect 11839 -10400 11895 -10356
rect 11939 -10400 11995 -10356
rect 12039 -10400 12095 -10356
rect 12139 -10400 12195 -10356
rect 12239 -10400 12295 -10356
rect 12339 -10400 12395 -10356
rect 12439 -10400 12495 -10356
rect 12539 -10400 12595 -10356
rect 12639 -10400 12695 -10356
rect 12739 -10400 13195 -10356
rect 13239 -10400 13295 -10356
rect 13339 -10400 13395 -10356
rect 13439 -10400 13495 -10356
rect 13539 -10400 13595 -10356
rect 13639 -10400 13695 -10356
rect 13739 -10400 13795 -10356
rect 13839 -10400 13895 -10356
rect 13939 -10400 13995 -10356
rect 14039 -10400 14095 -10356
rect 14139 -10400 14195 -10356
rect 14239 -10400 14295 -10356
rect 14339 -10400 14395 -10356
rect 14439 -10400 14495 -10356
rect 14539 -10400 14595 -10356
rect 14639 -10400 14695 -10356
rect 14739 -10400 15195 -10356
rect 15239 -10400 15295 -10356
rect 15339 -10400 15395 -10356
rect 15439 -10400 15495 -10356
rect 15539 -10400 15595 -10356
rect 15639 -10400 15695 -10356
rect 15739 -10400 15795 -10356
rect 15839 -10400 15895 -10356
rect 15939 -10400 15995 -10356
rect 16039 -10400 16095 -10356
rect 16139 -10400 16195 -10356
rect 16239 -10400 16295 -10356
rect 16339 -10400 16395 -10356
rect 16439 -10400 16495 -10356
rect 16539 -10400 16595 -10356
rect 16639 -10400 16695 -10356
rect 16739 -10400 18364 -10356
rect 7194 -10456 18364 -10400
rect 7194 -10500 9195 -10456
rect 9239 -10500 9295 -10456
rect 9339 -10500 9395 -10456
rect 9439 -10500 9495 -10456
rect 9539 -10500 9595 -10456
rect 9639 -10500 9695 -10456
rect 9739 -10500 9795 -10456
rect 9839 -10500 9895 -10456
rect 9939 -10500 9995 -10456
rect 10039 -10500 10095 -10456
rect 10139 -10500 10195 -10456
rect 10239 -10500 10295 -10456
rect 10339 -10500 10395 -10456
rect 10439 -10500 10495 -10456
rect 10539 -10500 10595 -10456
rect 10639 -10500 10695 -10456
rect 10739 -10500 11195 -10456
rect 11239 -10500 11295 -10456
rect 11339 -10500 11395 -10456
rect 11439 -10500 11495 -10456
rect 11539 -10500 11595 -10456
rect 11639 -10500 11695 -10456
rect 11739 -10500 11795 -10456
rect 11839 -10500 11895 -10456
rect 11939 -10500 11995 -10456
rect 12039 -10500 12095 -10456
rect 12139 -10500 12195 -10456
rect 12239 -10500 12295 -10456
rect 12339 -10500 12395 -10456
rect 12439 -10500 12495 -10456
rect 12539 -10500 12595 -10456
rect 12639 -10500 12695 -10456
rect 12739 -10500 13195 -10456
rect 13239 -10500 13295 -10456
rect 13339 -10500 13395 -10456
rect 13439 -10500 13495 -10456
rect 13539 -10500 13595 -10456
rect 13639 -10500 13695 -10456
rect 13739 -10500 13795 -10456
rect 13839 -10500 13895 -10456
rect 13939 -10500 13995 -10456
rect 14039 -10500 14095 -10456
rect 14139 -10500 14195 -10456
rect 14239 -10500 14295 -10456
rect 14339 -10500 14395 -10456
rect 14439 -10500 14495 -10456
rect 14539 -10500 14595 -10456
rect 14639 -10500 14695 -10456
rect 14739 -10500 15195 -10456
rect 15239 -10500 15295 -10456
rect 15339 -10500 15395 -10456
rect 15439 -10500 15495 -10456
rect 15539 -10500 15595 -10456
rect 15639 -10500 15695 -10456
rect 15739 -10500 15795 -10456
rect 15839 -10500 15895 -10456
rect 15939 -10500 15995 -10456
rect 16039 -10500 16095 -10456
rect 16139 -10500 16195 -10456
rect 16239 -10500 16295 -10456
rect 16339 -10500 16395 -10456
rect 16439 -10500 16495 -10456
rect 16539 -10500 16595 -10456
rect 16639 -10500 16695 -10456
rect 16739 -10500 18364 -10456
rect 7194 -10556 18364 -10500
rect 7194 -10600 9195 -10556
rect 9239 -10600 9295 -10556
rect 9339 -10600 9395 -10556
rect 9439 -10600 9495 -10556
rect 9539 -10600 9595 -10556
rect 9639 -10600 9695 -10556
rect 9739 -10600 9795 -10556
rect 9839 -10600 9895 -10556
rect 9939 -10600 9995 -10556
rect 10039 -10600 10095 -10556
rect 10139 -10600 10195 -10556
rect 10239 -10600 10295 -10556
rect 10339 -10600 10395 -10556
rect 10439 -10600 10495 -10556
rect 10539 -10600 10595 -10556
rect 10639 -10600 10695 -10556
rect 10739 -10600 11195 -10556
rect 11239 -10600 11295 -10556
rect 11339 -10600 11395 -10556
rect 11439 -10600 11495 -10556
rect 11539 -10600 11595 -10556
rect 11639 -10600 11695 -10556
rect 11739 -10600 11795 -10556
rect 11839 -10600 11895 -10556
rect 11939 -10600 11995 -10556
rect 12039 -10600 12095 -10556
rect 12139 -10600 12195 -10556
rect 12239 -10600 12295 -10556
rect 12339 -10600 12395 -10556
rect 12439 -10600 12495 -10556
rect 12539 -10600 12595 -10556
rect 12639 -10600 12695 -10556
rect 12739 -10600 13195 -10556
rect 13239 -10600 13295 -10556
rect 13339 -10600 13395 -10556
rect 13439 -10600 13495 -10556
rect 13539 -10600 13595 -10556
rect 13639 -10600 13695 -10556
rect 13739 -10600 13795 -10556
rect 13839 -10600 13895 -10556
rect 13939 -10600 13995 -10556
rect 14039 -10600 14095 -10556
rect 14139 -10600 14195 -10556
rect 14239 -10600 14295 -10556
rect 14339 -10600 14395 -10556
rect 14439 -10600 14495 -10556
rect 14539 -10600 14595 -10556
rect 14639 -10600 14695 -10556
rect 14739 -10600 15195 -10556
rect 15239 -10600 15295 -10556
rect 15339 -10600 15395 -10556
rect 15439 -10600 15495 -10556
rect 15539 -10600 15595 -10556
rect 15639 -10600 15695 -10556
rect 15739 -10600 15795 -10556
rect 15839 -10600 15895 -10556
rect 15939 -10600 15995 -10556
rect 16039 -10600 16095 -10556
rect 16139 -10600 16195 -10556
rect 16239 -10600 16295 -10556
rect 16339 -10600 16395 -10556
rect 16439 -10600 16495 -10556
rect 16539 -10600 16595 -10556
rect 16639 -10600 16695 -10556
rect 16739 -10600 18364 -10556
rect 7194 -10656 18364 -10600
rect 7194 -10700 9195 -10656
rect 9239 -10700 9295 -10656
rect 9339 -10700 9395 -10656
rect 9439 -10700 9495 -10656
rect 9539 -10700 9595 -10656
rect 9639 -10700 9695 -10656
rect 9739 -10700 9795 -10656
rect 9839 -10700 9895 -10656
rect 9939 -10700 9995 -10656
rect 10039 -10700 10095 -10656
rect 10139 -10700 10195 -10656
rect 10239 -10700 10295 -10656
rect 10339 -10700 10395 -10656
rect 10439 -10700 10495 -10656
rect 10539 -10700 10595 -10656
rect 10639 -10700 10695 -10656
rect 10739 -10700 11195 -10656
rect 11239 -10700 11295 -10656
rect 11339 -10700 11395 -10656
rect 11439 -10700 11495 -10656
rect 11539 -10700 11595 -10656
rect 11639 -10700 11695 -10656
rect 11739 -10700 11795 -10656
rect 11839 -10700 11895 -10656
rect 11939 -10700 11995 -10656
rect 12039 -10700 12095 -10656
rect 12139 -10700 12195 -10656
rect 12239 -10700 12295 -10656
rect 12339 -10700 12395 -10656
rect 12439 -10700 12495 -10656
rect 12539 -10700 12595 -10656
rect 12639 -10700 12695 -10656
rect 12739 -10700 13195 -10656
rect 13239 -10700 13295 -10656
rect 13339 -10700 13395 -10656
rect 13439 -10700 13495 -10656
rect 13539 -10700 13595 -10656
rect 13639 -10700 13695 -10656
rect 13739 -10700 13795 -10656
rect 13839 -10700 13895 -10656
rect 13939 -10700 13995 -10656
rect 14039 -10700 14095 -10656
rect 14139 -10700 14195 -10656
rect 14239 -10700 14295 -10656
rect 14339 -10700 14395 -10656
rect 14439 -10700 14495 -10656
rect 14539 -10700 14595 -10656
rect 14639 -10700 14695 -10656
rect 14739 -10700 15195 -10656
rect 15239 -10700 15295 -10656
rect 15339 -10700 15395 -10656
rect 15439 -10700 15495 -10656
rect 15539 -10700 15595 -10656
rect 15639 -10700 15695 -10656
rect 15739 -10700 15795 -10656
rect 15839 -10700 15895 -10656
rect 15939 -10700 15995 -10656
rect 16039 -10700 16095 -10656
rect 16139 -10700 16195 -10656
rect 16239 -10700 16295 -10656
rect 16339 -10700 16395 -10656
rect 16439 -10700 16495 -10656
rect 16539 -10700 16595 -10656
rect 16639 -10700 16695 -10656
rect 16739 -10700 18364 -10656
rect 7194 -10756 18364 -10700
rect 7194 -10800 9195 -10756
rect 9239 -10800 9295 -10756
rect 9339 -10800 9395 -10756
rect 9439 -10800 9495 -10756
rect 9539 -10800 9595 -10756
rect 9639 -10800 9695 -10756
rect 9739 -10800 9795 -10756
rect 9839 -10800 9895 -10756
rect 9939 -10800 9995 -10756
rect 10039 -10800 10095 -10756
rect 10139 -10800 10195 -10756
rect 10239 -10800 10295 -10756
rect 10339 -10800 10395 -10756
rect 10439 -10800 10495 -10756
rect 10539 -10800 10595 -10756
rect 10639 -10800 10695 -10756
rect 10739 -10800 11195 -10756
rect 11239 -10800 11295 -10756
rect 11339 -10800 11395 -10756
rect 11439 -10800 11495 -10756
rect 11539 -10800 11595 -10756
rect 11639 -10800 11695 -10756
rect 11739 -10800 11795 -10756
rect 11839 -10800 11895 -10756
rect 11939 -10800 11995 -10756
rect 12039 -10800 12095 -10756
rect 12139 -10800 12195 -10756
rect 12239 -10800 12295 -10756
rect 12339 -10800 12395 -10756
rect 12439 -10800 12495 -10756
rect 12539 -10800 12595 -10756
rect 12639 -10800 12695 -10756
rect 12739 -10800 13195 -10756
rect 13239 -10800 13295 -10756
rect 13339 -10800 13395 -10756
rect 13439 -10800 13495 -10756
rect 13539 -10800 13595 -10756
rect 13639 -10800 13695 -10756
rect 13739 -10800 13795 -10756
rect 13839 -10800 13895 -10756
rect 13939 -10800 13995 -10756
rect 14039 -10800 14095 -10756
rect 14139 -10800 14195 -10756
rect 14239 -10800 14295 -10756
rect 14339 -10800 14395 -10756
rect 14439 -10800 14495 -10756
rect 14539 -10800 14595 -10756
rect 14639 -10800 14695 -10756
rect 14739 -10800 15195 -10756
rect 15239 -10800 15295 -10756
rect 15339 -10800 15395 -10756
rect 15439 -10800 15495 -10756
rect 15539 -10800 15595 -10756
rect 15639 -10800 15695 -10756
rect 15739 -10800 15795 -10756
rect 15839 -10800 15895 -10756
rect 15939 -10800 15995 -10756
rect 16039 -10800 16095 -10756
rect 16139 -10800 16195 -10756
rect 16239 -10800 16295 -10756
rect 16339 -10800 16395 -10756
rect 16439 -10800 16495 -10756
rect 16539 -10800 16595 -10756
rect 16639 -10800 16695 -10756
rect 16739 -10800 18364 -10756
rect 7194 -10856 18364 -10800
rect 7194 -10900 9195 -10856
rect 9239 -10900 9295 -10856
rect 9339 -10900 9395 -10856
rect 9439 -10900 9495 -10856
rect 9539 -10900 9595 -10856
rect 9639 -10900 9695 -10856
rect 9739 -10900 9795 -10856
rect 9839 -10900 9895 -10856
rect 9939 -10900 9995 -10856
rect 10039 -10900 10095 -10856
rect 10139 -10900 10195 -10856
rect 10239 -10900 10295 -10856
rect 10339 -10900 10395 -10856
rect 10439 -10900 10495 -10856
rect 10539 -10900 10595 -10856
rect 10639 -10900 10695 -10856
rect 10739 -10900 11195 -10856
rect 11239 -10900 11295 -10856
rect 11339 -10900 11395 -10856
rect 11439 -10900 11495 -10856
rect 11539 -10900 11595 -10856
rect 11639 -10900 11695 -10856
rect 11739 -10900 11795 -10856
rect 11839 -10900 11895 -10856
rect 11939 -10900 11995 -10856
rect 12039 -10900 12095 -10856
rect 12139 -10900 12195 -10856
rect 12239 -10900 12295 -10856
rect 12339 -10900 12395 -10856
rect 12439 -10900 12495 -10856
rect 12539 -10900 12595 -10856
rect 12639 -10900 12695 -10856
rect 12739 -10900 13195 -10856
rect 13239 -10900 13295 -10856
rect 13339 -10900 13395 -10856
rect 13439 -10900 13495 -10856
rect 13539 -10900 13595 -10856
rect 13639 -10900 13695 -10856
rect 13739 -10900 13795 -10856
rect 13839 -10900 13895 -10856
rect 13939 -10900 13995 -10856
rect 14039 -10900 14095 -10856
rect 14139 -10900 14195 -10856
rect 14239 -10900 14295 -10856
rect 14339 -10900 14395 -10856
rect 14439 -10900 14495 -10856
rect 14539 -10900 14595 -10856
rect 14639 -10900 14695 -10856
rect 14739 -10900 15195 -10856
rect 15239 -10900 15295 -10856
rect 15339 -10900 15395 -10856
rect 15439 -10900 15495 -10856
rect 15539 -10900 15595 -10856
rect 15639 -10900 15695 -10856
rect 15739 -10900 15795 -10856
rect 15839 -10900 15895 -10856
rect 15939 -10900 15995 -10856
rect 16039 -10900 16095 -10856
rect 16139 -10900 16195 -10856
rect 16239 -10900 16295 -10856
rect 16339 -10900 16395 -10856
rect 16439 -10900 16495 -10856
rect 16539 -10900 16595 -10856
rect 16639 -10900 16695 -10856
rect 16739 -10900 18364 -10856
rect 7194 -10956 18364 -10900
rect 7194 -11000 9195 -10956
rect 9239 -11000 9295 -10956
rect 9339 -11000 9395 -10956
rect 9439 -11000 9495 -10956
rect 9539 -11000 9595 -10956
rect 9639 -11000 9695 -10956
rect 9739 -11000 9795 -10956
rect 9839 -11000 9895 -10956
rect 9939 -11000 9995 -10956
rect 10039 -11000 10095 -10956
rect 10139 -11000 10195 -10956
rect 10239 -11000 10295 -10956
rect 10339 -11000 10395 -10956
rect 10439 -11000 10495 -10956
rect 10539 -11000 10595 -10956
rect 10639 -11000 10695 -10956
rect 10739 -11000 11195 -10956
rect 11239 -11000 11295 -10956
rect 11339 -11000 11395 -10956
rect 11439 -11000 11495 -10956
rect 11539 -11000 11595 -10956
rect 11639 -11000 11695 -10956
rect 11739 -11000 11795 -10956
rect 11839 -11000 11895 -10956
rect 11939 -11000 11995 -10956
rect 12039 -11000 12095 -10956
rect 12139 -11000 12195 -10956
rect 12239 -11000 12295 -10956
rect 12339 -11000 12395 -10956
rect 12439 -11000 12495 -10956
rect 12539 -11000 12595 -10956
rect 12639 -11000 12695 -10956
rect 12739 -11000 13195 -10956
rect 13239 -11000 13295 -10956
rect 13339 -11000 13395 -10956
rect 13439 -11000 13495 -10956
rect 13539 -11000 13595 -10956
rect 13639 -11000 13695 -10956
rect 13739 -11000 13795 -10956
rect 13839 -11000 13895 -10956
rect 13939 -11000 13995 -10956
rect 14039 -11000 14095 -10956
rect 14139 -11000 14195 -10956
rect 14239 -11000 14295 -10956
rect 14339 -11000 14395 -10956
rect 14439 -11000 14495 -10956
rect 14539 -11000 14595 -10956
rect 14639 -11000 14695 -10956
rect 14739 -11000 15195 -10956
rect 15239 -11000 15295 -10956
rect 15339 -11000 15395 -10956
rect 15439 -11000 15495 -10956
rect 15539 -11000 15595 -10956
rect 15639 -11000 15695 -10956
rect 15739 -11000 15795 -10956
rect 15839 -11000 15895 -10956
rect 15939 -11000 15995 -10956
rect 16039 -11000 16095 -10956
rect 16139 -11000 16195 -10956
rect 16239 -11000 16295 -10956
rect 16339 -11000 16395 -10956
rect 16439 -11000 16495 -10956
rect 16539 -11000 16595 -10956
rect 16639 -11000 16695 -10956
rect 16739 -11000 18364 -10956
rect -16409 -13436 -2893 -11009
rect -16409 -13656 -12784 -13436
rect -12564 -13656 -12314 -13436
rect -12094 -13656 -11844 -13436
rect -11624 -13656 -11374 -13436
rect -11154 -13656 -10904 -13436
rect -10684 -13656 -10434 -13436
rect -10214 -13656 -9964 -13436
rect -9744 -13656 -9494 -13436
rect -9274 -13656 -9024 -13436
rect -8804 -13656 -8554 -13436
rect -8334 -13656 -8084 -13436
rect -7864 -13656 -7614 -13436
rect -7394 -13656 -7144 -13436
rect -6924 -13656 -6674 -13436
rect -6454 -13656 -2893 -13436
rect -105430 -135358 -104783 -135314
rect -104739 -135358 -104683 -135314
rect -104639 -135358 -104583 -135314
rect -104539 -135358 -104483 -135314
rect -104439 -135358 -104383 -135314
rect -104339 -135358 -104283 -135314
rect -104239 -135358 -104183 -135314
rect -104139 -135358 -104083 -135314
rect -104039 -135358 -103983 -135314
rect -103939 -135358 -103883 -135314
rect -103839 -135358 -103783 -135314
rect -103739 -135358 -103683 -135314
rect -103639 -135358 -103583 -135314
rect -103539 -135358 -103483 -135314
rect -103439 -135358 -103383 -135314
rect -103339 -135358 -103283 -135314
rect -103239 -135358 -102783 -135314
rect -102739 -135358 -102683 -135314
rect -102639 -135358 -102583 -135314
rect -102539 -135358 -102483 -135314
rect -102439 -135358 -102383 -135314
rect -102339 -135358 -102283 -135314
rect -102239 -135358 -102183 -135314
rect -102139 -135358 -102083 -135314
rect -102039 -135358 -101983 -135314
rect -101939 -135358 -101883 -135314
rect -101839 -135358 -101783 -135314
rect -101739 -135358 -101683 -135314
rect -101639 -135358 -101583 -135314
rect -101539 -135358 -101483 -135314
rect -101439 -135358 -101383 -135314
rect -101339 -135358 -101283 -135314
rect -101239 -135358 -100783 -135314
rect -100739 -135358 -100683 -135314
rect -100639 -135358 -100583 -135314
rect -100539 -135358 -100483 -135314
rect -100439 -135358 -100383 -135314
rect -100339 -135358 -100283 -135314
rect -100239 -135358 -100183 -135314
rect -100139 -135358 -100083 -135314
rect -100039 -135358 -99983 -135314
rect -99939 -135358 -99883 -135314
rect -99839 -135358 -99783 -135314
rect -99739 -135358 -99683 -135314
rect -99639 -135358 -99583 -135314
rect -99539 -135358 -99483 -135314
rect -99439 -135358 -99383 -135314
rect -99339 -135358 -99283 -135314
rect -99239 -135358 -98783 -135314
rect -98739 -135358 -98683 -135314
rect -98639 -135358 -98583 -135314
rect -98539 -135358 -98483 -135314
rect -98439 -135358 -98383 -135314
rect -98339 -135358 -98283 -135314
rect -98239 -135358 -98183 -135314
rect -98139 -135358 -98083 -135314
rect -98039 -135358 -97983 -135314
rect -97939 -135358 -97883 -135314
rect -97839 -135358 -97783 -135314
rect -97739 -135358 -97683 -135314
rect -97639 -135358 -97583 -135314
rect -97539 -135358 -97483 -135314
rect -97439 -135358 -97383 -135314
rect -97339 -135358 -97283 -135314
rect -97239 -135358 -96269 -135314
rect -105430 -135414 -96269 -135358
rect -105430 -135458 -104783 -135414
rect -104739 -135458 -104683 -135414
rect -104639 -135458 -104583 -135414
rect -104539 -135458 -104483 -135414
rect -104439 -135458 -104383 -135414
rect -104339 -135458 -104283 -135414
rect -104239 -135458 -104183 -135414
rect -104139 -135458 -104083 -135414
rect -104039 -135458 -103983 -135414
rect -103939 -135458 -103883 -135414
rect -103839 -135458 -103783 -135414
rect -103739 -135458 -103683 -135414
rect -103639 -135458 -103583 -135414
rect -103539 -135458 -103483 -135414
rect -103439 -135458 -103383 -135414
rect -103339 -135458 -103283 -135414
rect -103239 -135458 -102783 -135414
rect -102739 -135458 -102683 -135414
rect -102639 -135458 -102583 -135414
rect -102539 -135458 -102483 -135414
rect -102439 -135458 -102383 -135414
rect -102339 -135458 -102283 -135414
rect -102239 -135458 -102183 -135414
rect -102139 -135458 -102083 -135414
rect -102039 -135458 -101983 -135414
rect -101939 -135458 -101883 -135414
rect -101839 -135458 -101783 -135414
rect -101739 -135458 -101683 -135414
rect -101639 -135458 -101583 -135414
rect -101539 -135458 -101483 -135414
rect -101439 -135458 -101383 -135414
rect -101339 -135458 -101283 -135414
rect -101239 -135458 -100783 -135414
rect -100739 -135458 -100683 -135414
rect -100639 -135458 -100583 -135414
rect -100539 -135458 -100483 -135414
rect -100439 -135458 -100383 -135414
rect -100339 -135458 -100283 -135414
rect -100239 -135458 -100183 -135414
rect -100139 -135458 -100083 -135414
rect -100039 -135458 -99983 -135414
rect -99939 -135458 -99883 -135414
rect -99839 -135458 -99783 -135414
rect -99739 -135458 -99683 -135414
rect -99639 -135458 -99583 -135414
rect -99539 -135458 -99483 -135414
rect -99439 -135458 -99383 -135414
rect -99339 -135458 -99283 -135414
rect -99239 -135458 -98783 -135414
rect -98739 -135458 -98683 -135414
rect -98639 -135458 -98583 -135414
rect -98539 -135458 -98483 -135414
rect -98439 -135458 -98383 -135414
rect -98339 -135458 -98283 -135414
rect -98239 -135458 -98183 -135414
rect -98139 -135458 -98083 -135414
rect -98039 -135458 -97983 -135414
rect -97939 -135458 -97883 -135414
rect -97839 -135458 -97783 -135414
rect -97739 -135458 -97683 -135414
rect -97639 -135458 -97583 -135414
rect -97539 -135458 -97483 -135414
rect -97439 -135458 -97383 -135414
rect -97339 -135458 -97283 -135414
rect -97239 -135458 -96269 -135414
rect -105430 -135514 -96269 -135458
rect -105430 -135558 -104783 -135514
rect -104739 -135558 -104683 -135514
rect -104639 -135558 -104583 -135514
rect -104539 -135558 -104483 -135514
rect -104439 -135558 -104383 -135514
rect -104339 -135558 -104283 -135514
rect -104239 -135558 -104183 -135514
rect -104139 -135558 -104083 -135514
rect -104039 -135558 -103983 -135514
rect -103939 -135558 -103883 -135514
rect -103839 -135558 -103783 -135514
rect -103739 -135558 -103683 -135514
rect -103639 -135558 -103583 -135514
rect -103539 -135558 -103483 -135514
rect -103439 -135558 -103383 -135514
rect -103339 -135558 -103283 -135514
rect -103239 -135558 -102783 -135514
rect -102739 -135558 -102683 -135514
rect -102639 -135558 -102583 -135514
rect -102539 -135558 -102483 -135514
rect -102439 -135558 -102383 -135514
rect -102339 -135558 -102283 -135514
rect -102239 -135558 -102183 -135514
rect -102139 -135558 -102083 -135514
rect -102039 -135558 -101983 -135514
rect -101939 -135558 -101883 -135514
rect -101839 -135558 -101783 -135514
rect -101739 -135558 -101683 -135514
rect -101639 -135558 -101583 -135514
rect -101539 -135558 -101483 -135514
rect -101439 -135558 -101383 -135514
rect -101339 -135558 -101283 -135514
rect -101239 -135558 -100783 -135514
rect -100739 -135558 -100683 -135514
rect -100639 -135558 -100583 -135514
rect -100539 -135558 -100483 -135514
rect -100439 -135558 -100383 -135514
rect -100339 -135558 -100283 -135514
rect -100239 -135558 -100183 -135514
rect -100139 -135558 -100083 -135514
rect -100039 -135558 -99983 -135514
rect -99939 -135558 -99883 -135514
rect -99839 -135558 -99783 -135514
rect -99739 -135558 -99683 -135514
rect -99639 -135558 -99583 -135514
rect -99539 -135558 -99483 -135514
rect -99439 -135558 -99383 -135514
rect -99339 -135558 -99283 -135514
rect -99239 -135558 -98783 -135514
rect -98739 -135558 -98683 -135514
rect -98639 -135558 -98583 -135514
rect -98539 -135558 -98483 -135514
rect -98439 -135558 -98383 -135514
rect -98339 -135558 -98283 -135514
rect -98239 -135558 -98183 -135514
rect -98139 -135558 -98083 -135514
rect -98039 -135558 -97983 -135514
rect -97939 -135558 -97883 -135514
rect -97839 -135558 -97783 -135514
rect -97739 -135558 -97683 -135514
rect -97639 -135558 -97583 -135514
rect -97539 -135558 -97483 -135514
rect -97439 -135558 -97383 -135514
rect -97339 -135558 -97283 -135514
rect -97239 -135558 -96269 -135514
rect -105430 -135614 -96269 -135558
rect -105430 -135658 -104783 -135614
rect -104739 -135658 -104683 -135614
rect -104639 -135658 -104583 -135614
rect -104539 -135658 -104483 -135614
rect -104439 -135658 -104383 -135614
rect -104339 -135658 -104283 -135614
rect -104239 -135658 -104183 -135614
rect -104139 -135658 -104083 -135614
rect -104039 -135658 -103983 -135614
rect -103939 -135658 -103883 -135614
rect -103839 -135658 -103783 -135614
rect -103739 -135658 -103683 -135614
rect -103639 -135658 -103583 -135614
rect -103539 -135658 -103483 -135614
rect -103439 -135658 -103383 -135614
rect -103339 -135658 -103283 -135614
rect -103239 -135658 -102783 -135614
rect -102739 -135658 -102683 -135614
rect -102639 -135658 -102583 -135614
rect -102539 -135658 -102483 -135614
rect -102439 -135658 -102383 -135614
rect -102339 -135658 -102283 -135614
rect -102239 -135658 -102183 -135614
rect -102139 -135658 -102083 -135614
rect -102039 -135658 -101983 -135614
rect -101939 -135658 -101883 -135614
rect -101839 -135658 -101783 -135614
rect -101739 -135658 -101683 -135614
rect -101639 -135658 -101583 -135614
rect -101539 -135658 -101483 -135614
rect -101439 -135658 -101383 -135614
rect -101339 -135658 -101283 -135614
rect -101239 -135658 -100783 -135614
rect -100739 -135658 -100683 -135614
rect -100639 -135658 -100583 -135614
rect -100539 -135658 -100483 -135614
rect -100439 -135658 -100383 -135614
rect -100339 -135658 -100283 -135614
rect -100239 -135658 -100183 -135614
rect -100139 -135658 -100083 -135614
rect -100039 -135658 -99983 -135614
rect -99939 -135658 -99883 -135614
rect -99839 -135658 -99783 -135614
rect -99739 -135658 -99683 -135614
rect -99639 -135658 -99583 -135614
rect -99539 -135658 -99483 -135614
rect -99439 -135658 -99383 -135614
rect -99339 -135658 -99283 -135614
rect -99239 -135658 -98783 -135614
rect -98739 -135658 -98683 -135614
rect -98639 -135658 -98583 -135614
rect -98539 -135658 -98483 -135614
rect -98439 -135658 -98383 -135614
rect -98339 -135658 -98283 -135614
rect -98239 -135658 -98183 -135614
rect -98139 -135658 -98083 -135614
rect -98039 -135658 -97983 -135614
rect -97939 -135658 -97883 -135614
rect -97839 -135658 -97783 -135614
rect -97739 -135658 -97683 -135614
rect -97639 -135658 -97583 -135614
rect -97539 -135658 -97483 -135614
rect -97439 -135658 -97383 -135614
rect -97339 -135658 -97283 -135614
rect -97239 -135658 -96269 -135614
rect -105430 -135714 -96269 -135658
rect -105430 -135758 -104783 -135714
rect -104739 -135758 -104683 -135714
rect -104639 -135758 -104583 -135714
rect -104539 -135758 -104483 -135714
rect -104439 -135758 -104383 -135714
rect -104339 -135758 -104283 -135714
rect -104239 -135758 -104183 -135714
rect -104139 -135758 -104083 -135714
rect -104039 -135758 -103983 -135714
rect -103939 -135758 -103883 -135714
rect -103839 -135758 -103783 -135714
rect -103739 -135758 -103683 -135714
rect -103639 -135758 -103583 -135714
rect -103539 -135758 -103483 -135714
rect -103439 -135758 -103383 -135714
rect -103339 -135758 -103283 -135714
rect -103239 -135758 -102783 -135714
rect -102739 -135758 -102683 -135714
rect -102639 -135758 -102583 -135714
rect -102539 -135758 -102483 -135714
rect -102439 -135758 -102383 -135714
rect -102339 -135758 -102283 -135714
rect -102239 -135758 -102183 -135714
rect -102139 -135758 -102083 -135714
rect -102039 -135758 -101983 -135714
rect -101939 -135758 -101883 -135714
rect -101839 -135758 -101783 -135714
rect -101739 -135758 -101683 -135714
rect -101639 -135758 -101583 -135714
rect -101539 -135758 -101483 -135714
rect -101439 -135758 -101383 -135714
rect -101339 -135758 -101283 -135714
rect -101239 -135758 -100783 -135714
rect -100739 -135758 -100683 -135714
rect -100639 -135758 -100583 -135714
rect -100539 -135758 -100483 -135714
rect -100439 -135758 -100383 -135714
rect -100339 -135758 -100283 -135714
rect -100239 -135758 -100183 -135714
rect -100139 -135758 -100083 -135714
rect -100039 -135758 -99983 -135714
rect -99939 -135758 -99883 -135714
rect -99839 -135758 -99783 -135714
rect -99739 -135758 -99683 -135714
rect -99639 -135758 -99583 -135714
rect -99539 -135758 -99483 -135714
rect -99439 -135758 -99383 -135714
rect -99339 -135758 -99283 -135714
rect -99239 -135758 -98783 -135714
rect -98739 -135758 -98683 -135714
rect -98639 -135758 -98583 -135714
rect -98539 -135758 -98483 -135714
rect -98439 -135758 -98383 -135714
rect -98339 -135758 -98283 -135714
rect -98239 -135758 -98183 -135714
rect -98139 -135758 -98083 -135714
rect -98039 -135758 -97983 -135714
rect -97939 -135758 -97883 -135714
rect -97839 -135758 -97783 -135714
rect -97739 -135758 -97683 -135714
rect -97639 -135758 -97583 -135714
rect -97539 -135758 -97483 -135714
rect -97439 -135758 -97383 -135714
rect -97339 -135758 -97283 -135714
rect -97239 -135758 -96269 -135714
rect -105430 -135814 -96269 -135758
rect -105430 -135858 -104783 -135814
rect -104739 -135858 -104683 -135814
rect -104639 -135858 -104583 -135814
rect -104539 -135858 -104483 -135814
rect -104439 -135858 -104383 -135814
rect -104339 -135858 -104283 -135814
rect -104239 -135858 -104183 -135814
rect -104139 -135858 -104083 -135814
rect -104039 -135858 -103983 -135814
rect -103939 -135858 -103883 -135814
rect -103839 -135858 -103783 -135814
rect -103739 -135858 -103683 -135814
rect -103639 -135858 -103583 -135814
rect -103539 -135858 -103483 -135814
rect -103439 -135858 -103383 -135814
rect -103339 -135858 -103283 -135814
rect -103239 -135858 -102783 -135814
rect -102739 -135858 -102683 -135814
rect -102639 -135858 -102583 -135814
rect -102539 -135858 -102483 -135814
rect -102439 -135858 -102383 -135814
rect -102339 -135858 -102283 -135814
rect -102239 -135858 -102183 -135814
rect -102139 -135858 -102083 -135814
rect -102039 -135858 -101983 -135814
rect -101939 -135858 -101883 -135814
rect -101839 -135858 -101783 -135814
rect -101739 -135858 -101683 -135814
rect -101639 -135858 -101583 -135814
rect -101539 -135858 -101483 -135814
rect -101439 -135858 -101383 -135814
rect -101339 -135858 -101283 -135814
rect -101239 -135858 -100783 -135814
rect -100739 -135858 -100683 -135814
rect -100639 -135858 -100583 -135814
rect -100539 -135858 -100483 -135814
rect -100439 -135858 -100383 -135814
rect -100339 -135858 -100283 -135814
rect -100239 -135858 -100183 -135814
rect -100139 -135858 -100083 -135814
rect -100039 -135858 -99983 -135814
rect -99939 -135858 -99883 -135814
rect -99839 -135858 -99783 -135814
rect -99739 -135858 -99683 -135814
rect -99639 -135858 -99583 -135814
rect -99539 -135858 -99483 -135814
rect -99439 -135858 -99383 -135814
rect -99339 -135858 -99283 -135814
rect -99239 -135858 -98783 -135814
rect -98739 -135858 -98683 -135814
rect -98639 -135858 -98583 -135814
rect -98539 -135858 -98483 -135814
rect -98439 -135858 -98383 -135814
rect -98339 -135858 -98283 -135814
rect -98239 -135858 -98183 -135814
rect -98139 -135858 -98083 -135814
rect -98039 -135858 -97983 -135814
rect -97939 -135858 -97883 -135814
rect -97839 -135858 -97783 -135814
rect -97739 -135858 -97683 -135814
rect -97639 -135858 -97583 -135814
rect -97539 -135858 -97483 -135814
rect -97439 -135858 -97383 -135814
rect -97339 -135858 -97283 -135814
rect -97239 -135858 -96269 -135814
rect -105430 -135914 -96269 -135858
rect -105430 -135958 -104783 -135914
rect -104739 -135958 -104683 -135914
rect -104639 -135958 -104583 -135914
rect -104539 -135958 -104483 -135914
rect -104439 -135958 -104383 -135914
rect -104339 -135958 -104283 -135914
rect -104239 -135958 -104183 -135914
rect -104139 -135958 -104083 -135914
rect -104039 -135958 -103983 -135914
rect -103939 -135958 -103883 -135914
rect -103839 -135958 -103783 -135914
rect -103739 -135958 -103683 -135914
rect -103639 -135958 -103583 -135914
rect -103539 -135958 -103483 -135914
rect -103439 -135958 -103383 -135914
rect -103339 -135958 -103283 -135914
rect -103239 -135958 -102783 -135914
rect -102739 -135958 -102683 -135914
rect -102639 -135958 -102583 -135914
rect -102539 -135958 -102483 -135914
rect -102439 -135958 -102383 -135914
rect -102339 -135958 -102283 -135914
rect -102239 -135958 -102183 -135914
rect -102139 -135958 -102083 -135914
rect -102039 -135958 -101983 -135914
rect -101939 -135958 -101883 -135914
rect -101839 -135958 -101783 -135914
rect -101739 -135958 -101683 -135914
rect -101639 -135958 -101583 -135914
rect -101539 -135958 -101483 -135914
rect -101439 -135958 -101383 -135914
rect -101339 -135958 -101283 -135914
rect -101239 -135958 -100783 -135914
rect -100739 -135958 -100683 -135914
rect -100639 -135958 -100583 -135914
rect -100539 -135958 -100483 -135914
rect -100439 -135958 -100383 -135914
rect -100339 -135958 -100283 -135914
rect -100239 -135958 -100183 -135914
rect -100139 -135958 -100083 -135914
rect -100039 -135958 -99983 -135914
rect -99939 -135958 -99883 -135914
rect -99839 -135958 -99783 -135914
rect -99739 -135958 -99683 -135914
rect -99639 -135958 -99583 -135914
rect -99539 -135958 -99483 -135914
rect -99439 -135958 -99383 -135914
rect -99339 -135958 -99283 -135914
rect -99239 -135958 -98783 -135914
rect -98739 -135958 -98683 -135914
rect -98639 -135958 -98583 -135914
rect -98539 -135958 -98483 -135914
rect -98439 -135958 -98383 -135914
rect -98339 -135958 -98283 -135914
rect -98239 -135958 -98183 -135914
rect -98139 -135958 -98083 -135914
rect -98039 -135958 -97983 -135914
rect -97939 -135958 -97883 -135914
rect -97839 -135958 -97783 -135914
rect -97739 -135958 -97683 -135914
rect -97639 -135958 -97583 -135914
rect -97539 -135958 -97483 -135914
rect -97439 -135958 -97383 -135914
rect -97339 -135958 -97283 -135914
rect -97239 -135958 -96269 -135914
rect -105430 -136014 -96269 -135958
rect -105430 -136058 -104783 -136014
rect -104739 -136058 -104683 -136014
rect -104639 -136058 -104583 -136014
rect -104539 -136058 -104483 -136014
rect -104439 -136058 -104383 -136014
rect -104339 -136058 -104283 -136014
rect -104239 -136058 -104183 -136014
rect -104139 -136058 -104083 -136014
rect -104039 -136058 -103983 -136014
rect -103939 -136058 -103883 -136014
rect -103839 -136058 -103783 -136014
rect -103739 -136058 -103683 -136014
rect -103639 -136058 -103583 -136014
rect -103539 -136058 -103483 -136014
rect -103439 -136058 -103383 -136014
rect -103339 -136058 -103283 -136014
rect -103239 -136058 -102783 -136014
rect -102739 -136058 -102683 -136014
rect -102639 -136058 -102583 -136014
rect -102539 -136058 -102483 -136014
rect -102439 -136058 -102383 -136014
rect -102339 -136058 -102283 -136014
rect -102239 -136058 -102183 -136014
rect -102139 -136058 -102083 -136014
rect -102039 -136058 -101983 -136014
rect -101939 -136058 -101883 -136014
rect -101839 -136058 -101783 -136014
rect -101739 -136058 -101683 -136014
rect -101639 -136058 -101583 -136014
rect -101539 -136058 -101483 -136014
rect -101439 -136058 -101383 -136014
rect -101339 -136058 -101283 -136014
rect -101239 -136058 -100783 -136014
rect -100739 -136058 -100683 -136014
rect -100639 -136058 -100583 -136014
rect -100539 -136058 -100483 -136014
rect -100439 -136058 -100383 -136014
rect -100339 -136058 -100283 -136014
rect -100239 -136058 -100183 -136014
rect -100139 -136058 -100083 -136014
rect -100039 -136058 -99983 -136014
rect -99939 -136058 -99883 -136014
rect -99839 -136058 -99783 -136014
rect -99739 -136058 -99683 -136014
rect -99639 -136058 -99583 -136014
rect -99539 -136058 -99483 -136014
rect -99439 -136058 -99383 -136014
rect -99339 -136058 -99283 -136014
rect -99239 -136058 -98783 -136014
rect -98739 -136058 -98683 -136014
rect -98639 -136058 -98583 -136014
rect -98539 -136058 -98483 -136014
rect -98439 -136058 -98383 -136014
rect -98339 -136058 -98283 -136014
rect -98239 -136058 -98183 -136014
rect -98139 -136058 -98083 -136014
rect -98039 -136058 -97983 -136014
rect -97939 -136058 -97883 -136014
rect -97839 -136058 -97783 -136014
rect -97739 -136058 -97683 -136014
rect -97639 -136058 -97583 -136014
rect -97539 -136058 -97483 -136014
rect -97439 -136058 -97383 -136014
rect -97339 -136058 -97283 -136014
rect -97239 -136058 -96269 -136014
rect -105430 -136114 -96269 -136058
rect -105430 -136158 -104783 -136114
rect -104739 -136158 -104683 -136114
rect -104639 -136158 -104583 -136114
rect -104539 -136158 -104483 -136114
rect -104439 -136158 -104383 -136114
rect -104339 -136158 -104283 -136114
rect -104239 -136158 -104183 -136114
rect -104139 -136158 -104083 -136114
rect -104039 -136158 -103983 -136114
rect -103939 -136158 -103883 -136114
rect -103839 -136158 -103783 -136114
rect -103739 -136158 -103683 -136114
rect -103639 -136158 -103583 -136114
rect -103539 -136158 -103483 -136114
rect -103439 -136158 -103383 -136114
rect -103339 -136158 -103283 -136114
rect -103239 -136158 -102783 -136114
rect -102739 -136158 -102683 -136114
rect -102639 -136158 -102583 -136114
rect -102539 -136158 -102483 -136114
rect -102439 -136158 -102383 -136114
rect -102339 -136158 -102283 -136114
rect -102239 -136158 -102183 -136114
rect -102139 -136158 -102083 -136114
rect -102039 -136158 -101983 -136114
rect -101939 -136158 -101883 -136114
rect -101839 -136158 -101783 -136114
rect -101739 -136158 -101683 -136114
rect -101639 -136158 -101583 -136114
rect -101539 -136158 -101483 -136114
rect -101439 -136158 -101383 -136114
rect -101339 -136158 -101283 -136114
rect -101239 -136158 -100783 -136114
rect -100739 -136158 -100683 -136114
rect -100639 -136158 -100583 -136114
rect -100539 -136158 -100483 -136114
rect -100439 -136158 -100383 -136114
rect -100339 -136158 -100283 -136114
rect -100239 -136158 -100183 -136114
rect -100139 -136158 -100083 -136114
rect -100039 -136158 -99983 -136114
rect -99939 -136158 -99883 -136114
rect -99839 -136158 -99783 -136114
rect -99739 -136158 -99683 -136114
rect -99639 -136158 -99583 -136114
rect -99539 -136158 -99483 -136114
rect -99439 -136158 -99383 -136114
rect -99339 -136158 -99283 -136114
rect -99239 -136158 -98783 -136114
rect -98739 -136158 -98683 -136114
rect -98639 -136158 -98583 -136114
rect -98539 -136158 -98483 -136114
rect -98439 -136158 -98383 -136114
rect -98339 -136158 -98283 -136114
rect -98239 -136158 -98183 -136114
rect -98139 -136158 -98083 -136114
rect -98039 -136158 -97983 -136114
rect -97939 -136158 -97883 -136114
rect -97839 -136158 -97783 -136114
rect -97739 -136158 -97683 -136114
rect -97639 -136158 -97583 -136114
rect -97539 -136158 -97483 -136114
rect -97439 -136158 -97383 -136114
rect -97339 -136158 -97283 -136114
rect -97239 -136158 -96269 -136114
rect -105430 -136214 -96269 -136158
rect -105430 -136258 -104783 -136214
rect -104739 -136258 -104683 -136214
rect -104639 -136258 -104583 -136214
rect -104539 -136258 -104483 -136214
rect -104439 -136258 -104383 -136214
rect -104339 -136258 -104283 -136214
rect -104239 -136258 -104183 -136214
rect -104139 -136258 -104083 -136214
rect -104039 -136258 -103983 -136214
rect -103939 -136258 -103883 -136214
rect -103839 -136258 -103783 -136214
rect -103739 -136258 -103683 -136214
rect -103639 -136258 -103583 -136214
rect -103539 -136258 -103483 -136214
rect -103439 -136258 -103383 -136214
rect -103339 -136258 -103283 -136214
rect -103239 -136258 -102783 -136214
rect -102739 -136258 -102683 -136214
rect -102639 -136258 -102583 -136214
rect -102539 -136258 -102483 -136214
rect -102439 -136258 -102383 -136214
rect -102339 -136258 -102283 -136214
rect -102239 -136258 -102183 -136214
rect -102139 -136258 -102083 -136214
rect -102039 -136258 -101983 -136214
rect -101939 -136258 -101883 -136214
rect -101839 -136258 -101783 -136214
rect -101739 -136258 -101683 -136214
rect -101639 -136258 -101583 -136214
rect -101539 -136258 -101483 -136214
rect -101439 -136258 -101383 -136214
rect -101339 -136258 -101283 -136214
rect -101239 -136258 -100783 -136214
rect -100739 -136258 -100683 -136214
rect -100639 -136258 -100583 -136214
rect -100539 -136258 -100483 -136214
rect -100439 -136258 -100383 -136214
rect -100339 -136258 -100283 -136214
rect -100239 -136258 -100183 -136214
rect -100139 -136258 -100083 -136214
rect -100039 -136258 -99983 -136214
rect -99939 -136258 -99883 -136214
rect -99839 -136258 -99783 -136214
rect -99739 -136258 -99683 -136214
rect -99639 -136258 -99583 -136214
rect -99539 -136258 -99483 -136214
rect -99439 -136258 -99383 -136214
rect -99339 -136258 -99283 -136214
rect -99239 -136258 -98783 -136214
rect -98739 -136258 -98683 -136214
rect -98639 -136258 -98583 -136214
rect -98539 -136258 -98483 -136214
rect -98439 -136258 -98383 -136214
rect -98339 -136258 -98283 -136214
rect -98239 -136258 -98183 -136214
rect -98139 -136258 -98083 -136214
rect -98039 -136258 -97983 -136214
rect -97939 -136258 -97883 -136214
rect -97839 -136258 -97783 -136214
rect -97739 -136258 -97683 -136214
rect -97639 -136258 -97583 -136214
rect -97539 -136258 -97483 -136214
rect -97439 -136258 -97383 -136214
rect -97339 -136258 -97283 -136214
rect -97239 -136258 -96269 -136214
rect -105430 -136314 -96269 -136258
rect -105430 -136358 -104783 -136314
rect -104739 -136358 -104683 -136314
rect -104639 -136358 -104583 -136314
rect -104539 -136358 -104483 -136314
rect -104439 -136358 -104383 -136314
rect -104339 -136358 -104283 -136314
rect -104239 -136358 -104183 -136314
rect -104139 -136358 -104083 -136314
rect -104039 -136358 -103983 -136314
rect -103939 -136358 -103883 -136314
rect -103839 -136358 -103783 -136314
rect -103739 -136358 -103683 -136314
rect -103639 -136358 -103583 -136314
rect -103539 -136358 -103483 -136314
rect -103439 -136358 -103383 -136314
rect -103339 -136358 -103283 -136314
rect -103239 -136358 -102783 -136314
rect -102739 -136358 -102683 -136314
rect -102639 -136358 -102583 -136314
rect -102539 -136358 -102483 -136314
rect -102439 -136358 -102383 -136314
rect -102339 -136358 -102283 -136314
rect -102239 -136358 -102183 -136314
rect -102139 -136358 -102083 -136314
rect -102039 -136358 -101983 -136314
rect -101939 -136358 -101883 -136314
rect -101839 -136358 -101783 -136314
rect -101739 -136358 -101683 -136314
rect -101639 -136358 -101583 -136314
rect -101539 -136358 -101483 -136314
rect -101439 -136358 -101383 -136314
rect -101339 -136358 -101283 -136314
rect -101239 -136358 -100783 -136314
rect -100739 -136358 -100683 -136314
rect -100639 -136358 -100583 -136314
rect -100539 -136358 -100483 -136314
rect -100439 -136358 -100383 -136314
rect -100339 -136358 -100283 -136314
rect -100239 -136358 -100183 -136314
rect -100139 -136358 -100083 -136314
rect -100039 -136358 -99983 -136314
rect -99939 -136358 -99883 -136314
rect -99839 -136358 -99783 -136314
rect -99739 -136358 -99683 -136314
rect -99639 -136358 -99583 -136314
rect -99539 -136358 -99483 -136314
rect -99439 -136358 -99383 -136314
rect -99339 -136358 -99283 -136314
rect -99239 -136358 -98783 -136314
rect -98739 -136358 -98683 -136314
rect -98639 -136358 -98583 -136314
rect -98539 -136358 -98483 -136314
rect -98439 -136358 -98383 -136314
rect -98339 -136358 -98283 -136314
rect -98239 -136358 -98183 -136314
rect -98139 -136358 -98083 -136314
rect -98039 -136358 -97983 -136314
rect -97939 -136358 -97883 -136314
rect -97839 -136358 -97783 -136314
rect -97739 -136358 -97683 -136314
rect -97639 -136358 -97583 -136314
rect -97539 -136358 -97483 -136314
rect -97439 -136358 -97383 -136314
rect -97339 -136358 -97283 -136314
rect -97239 -136358 -96269 -136314
rect -105430 -136414 -96269 -136358
rect -105430 -136458 -104783 -136414
rect -104739 -136458 -104683 -136414
rect -104639 -136458 -104583 -136414
rect -104539 -136458 -104483 -136414
rect -104439 -136458 -104383 -136414
rect -104339 -136458 -104283 -136414
rect -104239 -136458 -104183 -136414
rect -104139 -136458 -104083 -136414
rect -104039 -136458 -103983 -136414
rect -103939 -136458 -103883 -136414
rect -103839 -136458 -103783 -136414
rect -103739 -136458 -103683 -136414
rect -103639 -136458 -103583 -136414
rect -103539 -136458 -103483 -136414
rect -103439 -136458 -103383 -136414
rect -103339 -136458 -103283 -136414
rect -103239 -136458 -102783 -136414
rect -102739 -136458 -102683 -136414
rect -102639 -136458 -102583 -136414
rect -102539 -136458 -102483 -136414
rect -102439 -136458 -102383 -136414
rect -102339 -136458 -102283 -136414
rect -102239 -136458 -102183 -136414
rect -102139 -136458 -102083 -136414
rect -102039 -136458 -101983 -136414
rect -101939 -136458 -101883 -136414
rect -101839 -136458 -101783 -136414
rect -101739 -136458 -101683 -136414
rect -101639 -136458 -101583 -136414
rect -101539 -136458 -101483 -136414
rect -101439 -136458 -101383 -136414
rect -101339 -136458 -101283 -136414
rect -101239 -136458 -100783 -136414
rect -100739 -136458 -100683 -136414
rect -100639 -136458 -100583 -136414
rect -100539 -136458 -100483 -136414
rect -100439 -136458 -100383 -136414
rect -100339 -136458 -100283 -136414
rect -100239 -136458 -100183 -136414
rect -100139 -136458 -100083 -136414
rect -100039 -136458 -99983 -136414
rect -99939 -136458 -99883 -136414
rect -99839 -136458 -99783 -136414
rect -99739 -136458 -99683 -136414
rect -99639 -136458 -99583 -136414
rect -99539 -136458 -99483 -136414
rect -99439 -136458 -99383 -136414
rect -99339 -136458 -99283 -136414
rect -99239 -136458 -98783 -136414
rect -98739 -136458 -98683 -136414
rect -98639 -136458 -98583 -136414
rect -98539 -136458 -98483 -136414
rect -98439 -136458 -98383 -136414
rect -98339 -136458 -98283 -136414
rect -98239 -136458 -98183 -136414
rect -98139 -136458 -98083 -136414
rect -98039 -136458 -97983 -136414
rect -97939 -136458 -97883 -136414
rect -97839 -136458 -97783 -136414
rect -97739 -136458 -97683 -136414
rect -97639 -136458 -97583 -136414
rect -97539 -136458 -97483 -136414
rect -97439 -136458 -97383 -136414
rect -97339 -136458 -97283 -136414
rect -97239 -136458 -96269 -136414
rect -105430 -136514 -96269 -136458
rect -105430 -136558 -104783 -136514
rect -104739 -136558 -104683 -136514
rect -104639 -136558 -104583 -136514
rect -104539 -136558 -104483 -136514
rect -104439 -136558 -104383 -136514
rect -104339 -136558 -104283 -136514
rect -104239 -136558 -104183 -136514
rect -104139 -136558 -104083 -136514
rect -104039 -136558 -103983 -136514
rect -103939 -136558 -103883 -136514
rect -103839 -136558 -103783 -136514
rect -103739 -136558 -103683 -136514
rect -103639 -136558 -103583 -136514
rect -103539 -136558 -103483 -136514
rect -103439 -136558 -103383 -136514
rect -103339 -136558 -103283 -136514
rect -103239 -136558 -102783 -136514
rect -102739 -136558 -102683 -136514
rect -102639 -136558 -102583 -136514
rect -102539 -136558 -102483 -136514
rect -102439 -136558 -102383 -136514
rect -102339 -136558 -102283 -136514
rect -102239 -136558 -102183 -136514
rect -102139 -136558 -102083 -136514
rect -102039 -136558 -101983 -136514
rect -101939 -136558 -101883 -136514
rect -101839 -136558 -101783 -136514
rect -101739 -136558 -101683 -136514
rect -101639 -136558 -101583 -136514
rect -101539 -136558 -101483 -136514
rect -101439 -136558 -101383 -136514
rect -101339 -136558 -101283 -136514
rect -101239 -136558 -100783 -136514
rect -100739 -136558 -100683 -136514
rect -100639 -136558 -100583 -136514
rect -100539 -136558 -100483 -136514
rect -100439 -136558 -100383 -136514
rect -100339 -136558 -100283 -136514
rect -100239 -136558 -100183 -136514
rect -100139 -136558 -100083 -136514
rect -100039 -136558 -99983 -136514
rect -99939 -136558 -99883 -136514
rect -99839 -136558 -99783 -136514
rect -99739 -136558 -99683 -136514
rect -99639 -136558 -99583 -136514
rect -99539 -136558 -99483 -136514
rect -99439 -136558 -99383 -136514
rect -99339 -136558 -99283 -136514
rect -99239 -136558 -98783 -136514
rect -98739 -136558 -98683 -136514
rect -98639 -136558 -98583 -136514
rect -98539 -136558 -98483 -136514
rect -98439 -136558 -98383 -136514
rect -98339 -136558 -98283 -136514
rect -98239 -136558 -98183 -136514
rect -98139 -136558 -98083 -136514
rect -98039 -136558 -97983 -136514
rect -97939 -136558 -97883 -136514
rect -97839 -136558 -97783 -136514
rect -97739 -136558 -97683 -136514
rect -97639 -136558 -97583 -136514
rect -97539 -136558 -97483 -136514
rect -97439 -136558 -97383 -136514
rect -97339 -136558 -97283 -136514
rect -97239 -136558 -96269 -136514
rect -105430 -136614 -96269 -136558
rect -105430 -136658 -104783 -136614
rect -104739 -136658 -104683 -136614
rect -104639 -136658 -104583 -136614
rect -104539 -136658 -104483 -136614
rect -104439 -136658 -104383 -136614
rect -104339 -136658 -104283 -136614
rect -104239 -136658 -104183 -136614
rect -104139 -136658 -104083 -136614
rect -104039 -136658 -103983 -136614
rect -103939 -136658 -103883 -136614
rect -103839 -136658 -103783 -136614
rect -103739 -136658 -103683 -136614
rect -103639 -136658 -103583 -136614
rect -103539 -136658 -103483 -136614
rect -103439 -136658 -103383 -136614
rect -103339 -136658 -103283 -136614
rect -103239 -136658 -102783 -136614
rect -102739 -136658 -102683 -136614
rect -102639 -136658 -102583 -136614
rect -102539 -136658 -102483 -136614
rect -102439 -136658 -102383 -136614
rect -102339 -136658 -102283 -136614
rect -102239 -136658 -102183 -136614
rect -102139 -136658 -102083 -136614
rect -102039 -136658 -101983 -136614
rect -101939 -136658 -101883 -136614
rect -101839 -136658 -101783 -136614
rect -101739 -136658 -101683 -136614
rect -101639 -136658 -101583 -136614
rect -101539 -136658 -101483 -136614
rect -101439 -136658 -101383 -136614
rect -101339 -136658 -101283 -136614
rect -101239 -136658 -100783 -136614
rect -100739 -136658 -100683 -136614
rect -100639 -136658 -100583 -136614
rect -100539 -136658 -100483 -136614
rect -100439 -136658 -100383 -136614
rect -100339 -136658 -100283 -136614
rect -100239 -136658 -100183 -136614
rect -100139 -136658 -100083 -136614
rect -100039 -136658 -99983 -136614
rect -99939 -136658 -99883 -136614
rect -99839 -136658 -99783 -136614
rect -99739 -136658 -99683 -136614
rect -99639 -136658 -99583 -136614
rect -99539 -136658 -99483 -136614
rect -99439 -136658 -99383 -136614
rect -99339 -136658 -99283 -136614
rect -99239 -136658 -98783 -136614
rect -98739 -136658 -98683 -136614
rect -98639 -136658 -98583 -136614
rect -98539 -136658 -98483 -136614
rect -98439 -136658 -98383 -136614
rect -98339 -136658 -98283 -136614
rect -98239 -136658 -98183 -136614
rect -98139 -136658 -98083 -136614
rect -98039 -136658 -97983 -136614
rect -97939 -136658 -97883 -136614
rect -97839 -136658 -97783 -136614
rect -97739 -136658 -97683 -136614
rect -97639 -136658 -97583 -136614
rect -97539 -136658 -97483 -136614
rect -97439 -136658 -97383 -136614
rect -97339 -136658 -97283 -136614
rect -97239 -136658 -96269 -136614
rect -105430 -136714 -96269 -136658
rect -105430 -136758 -104783 -136714
rect -104739 -136758 -104683 -136714
rect -104639 -136758 -104583 -136714
rect -104539 -136758 -104483 -136714
rect -104439 -136758 -104383 -136714
rect -104339 -136758 -104283 -136714
rect -104239 -136758 -104183 -136714
rect -104139 -136758 -104083 -136714
rect -104039 -136758 -103983 -136714
rect -103939 -136758 -103883 -136714
rect -103839 -136758 -103783 -136714
rect -103739 -136758 -103683 -136714
rect -103639 -136758 -103583 -136714
rect -103539 -136758 -103483 -136714
rect -103439 -136758 -103383 -136714
rect -103339 -136758 -103283 -136714
rect -103239 -136758 -102783 -136714
rect -102739 -136758 -102683 -136714
rect -102639 -136758 -102583 -136714
rect -102539 -136758 -102483 -136714
rect -102439 -136758 -102383 -136714
rect -102339 -136758 -102283 -136714
rect -102239 -136758 -102183 -136714
rect -102139 -136758 -102083 -136714
rect -102039 -136758 -101983 -136714
rect -101939 -136758 -101883 -136714
rect -101839 -136758 -101783 -136714
rect -101739 -136758 -101683 -136714
rect -101639 -136758 -101583 -136714
rect -101539 -136758 -101483 -136714
rect -101439 -136758 -101383 -136714
rect -101339 -136758 -101283 -136714
rect -101239 -136758 -100783 -136714
rect -100739 -136758 -100683 -136714
rect -100639 -136758 -100583 -136714
rect -100539 -136758 -100483 -136714
rect -100439 -136758 -100383 -136714
rect -100339 -136758 -100283 -136714
rect -100239 -136758 -100183 -136714
rect -100139 -136758 -100083 -136714
rect -100039 -136758 -99983 -136714
rect -99939 -136758 -99883 -136714
rect -99839 -136758 -99783 -136714
rect -99739 -136758 -99683 -136714
rect -99639 -136758 -99583 -136714
rect -99539 -136758 -99483 -136714
rect -99439 -136758 -99383 -136714
rect -99339 -136758 -99283 -136714
rect -99239 -136758 -98783 -136714
rect -98739 -136758 -98683 -136714
rect -98639 -136758 -98583 -136714
rect -98539 -136758 -98483 -136714
rect -98439 -136758 -98383 -136714
rect -98339 -136758 -98283 -136714
rect -98239 -136758 -98183 -136714
rect -98139 -136758 -98083 -136714
rect -98039 -136758 -97983 -136714
rect -97939 -136758 -97883 -136714
rect -97839 -136758 -97783 -136714
rect -97739 -136758 -97683 -136714
rect -97639 -136758 -97583 -136714
rect -97539 -136758 -97483 -136714
rect -97439 -136758 -97383 -136714
rect -97339 -136758 -97283 -136714
rect -97239 -136758 -96269 -136714
rect -105430 -136814 -96269 -136758
rect -105430 -136858 -104783 -136814
rect -104739 -136858 -104683 -136814
rect -104639 -136858 -104583 -136814
rect -104539 -136858 -104483 -136814
rect -104439 -136858 -104383 -136814
rect -104339 -136858 -104283 -136814
rect -104239 -136858 -104183 -136814
rect -104139 -136858 -104083 -136814
rect -104039 -136858 -103983 -136814
rect -103939 -136858 -103883 -136814
rect -103839 -136858 -103783 -136814
rect -103739 -136858 -103683 -136814
rect -103639 -136858 -103583 -136814
rect -103539 -136858 -103483 -136814
rect -103439 -136858 -103383 -136814
rect -103339 -136858 -103283 -136814
rect -103239 -136858 -102783 -136814
rect -102739 -136858 -102683 -136814
rect -102639 -136858 -102583 -136814
rect -102539 -136858 -102483 -136814
rect -102439 -136858 -102383 -136814
rect -102339 -136858 -102283 -136814
rect -102239 -136858 -102183 -136814
rect -102139 -136858 -102083 -136814
rect -102039 -136858 -101983 -136814
rect -101939 -136858 -101883 -136814
rect -101839 -136858 -101783 -136814
rect -101739 -136858 -101683 -136814
rect -101639 -136858 -101583 -136814
rect -101539 -136858 -101483 -136814
rect -101439 -136858 -101383 -136814
rect -101339 -136858 -101283 -136814
rect -101239 -136858 -100783 -136814
rect -100739 -136858 -100683 -136814
rect -100639 -136858 -100583 -136814
rect -100539 -136858 -100483 -136814
rect -100439 -136858 -100383 -136814
rect -100339 -136858 -100283 -136814
rect -100239 -136858 -100183 -136814
rect -100139 -136858 -100083 -136814
rect -100039 -136858 -99983 -136814
rect -99939 -136858 -99883 -136814
rect -99839 -136858 -99783 -136814
rect -99739 -136858 -99683 -136814
rect -99639 -136858 -99583 -136814
rect -99539 -136858 -99483 -136814
rect -99439 -136858 -99383 -136814
rect -99339 -136858 -99283 -136814
rect -99239 -136858 -98783 -136814
rect -98739 -136858 -98683 -136814
rect -98639 -136858 -98583 -136814
rect -98539 -136858 -98483 -136814
rect -98439 -136858 -98383 -136814
rect -98339 -136858 -98283 -136814
rect -98239 -136858 -98183 -136814
rect -98139 -136858 -98083 -136814
rect -98039 -136858 -97983 -136814
rect -97939 -136858 -97883 -136814
rect -97839 -136858 -97783 -136814
rect -97739 -136858 -97683 -136814
rect -97639 -136858 -97583 -136814
rect -97539 -136858 -97483 -136814
rect -97439 -136858 -97383 -136814
rect -97339 -136858 -97283 -136814
rect -97239 -136858 -96269 -136814
rect -105430 -137375 -96269 -136858
rect -87194 -24366 -71799 -23015
rect -87194 -24410 -82799 -24366
rect -82755 -24410 -82699 -24366
rect -82655 -24410 -82599 -24366
rect -82555 -24410 -82499 -24366
rect -82455 -24410 -82399 -24366
rect -82355 -24410 -82299 -24366
rect -82255 -24410 -82199 -24366
rect -82155 -24410 -82099 -24366
rect -82055 -24410 -81999 -24366
rect -81955 -24410 -81899 -24366
rect -81855 -24410 -81799 -24366
rect -81755 -24410 -81699 -24366
rect -81655 -24410 -81599 -24366
rect -81555 -24410 -81499 -24366
rect -81455 -24410 -81399 -24366
rect -81355 -24410 -81299 -24366
rect -81255 -24410 -80799 -24366
rect -80755 -24410 -80699 -24366
rect -80655 -24410 -80599 -24366
rect -80555 -24410 -80499 -24366
rect -80455 -24410 -80399 -24366
rect -80355 -24410 -80299 -24366
rect -80255 -24410 -80199 -24366
rect -80155 -24410 -80099 -24366
rect -80055 -24410 -79999 -24366
rect -79955 -24410 -79899 -24366
rect -79855 -24410 -79799 -24366
rect -79755 -24410 -79699 -24366
rect -79655 -24410 -79599 -24366
rect -79555 -24410 -79499 -24366
rect -79455 -24410 -79399 -24366
rect -79355 -24410 -79299 -24366
rect -79255 -24410 -78799 -24366
rect -78755 -24410 -78699 -24366
rect -78655 -24410 -78599 -24366
rect -78555 -24410 -78499 -24366
rect -78455 -24410 -78399 -24366
rect -78355 -24410 -78299 -24366
rect -78255 -24410 -78199 -24366
rect -78155 -24410 -78099 -24366
rect -78055 -24410 -77999 -24366
rect -77955 -24410 -77899 -24366
rect -77855 -24410 -77799 -24366
rect -77755 -24410 -77699 -24366
rect -77655 -24410 -77599 -24366
rect -77555 -24410 -77499 -24366
rect -77455 -24410 -77399 -24366
rect -77355 -24410 -77299 -24366
rect -77255 -24410 -76799 -24366
rect -76755 -24410 -76699 -24366
rect -76655 -24410 -76599 -24366
rect -76555 -24410 -76499 -24366
rect -76455 -24410 -76399 -24366
rect -76355 -24410 -76299 -24366
rect -76255 -24410 -76199 -24366
rect -76155 -24410 -76099 -24366
rect -76055 -24410 -75999 -24366
rect -75955 -24410 -75899 -24366
rect -75855 -24410 -75799 -24366
rect -75755 -24410 -75699 -24366
rect -75655 -24410 -75599 -24366
rect -75555 -24410 -75499 -24366
rect -75455 -24410 -75399 -24366
rect -75355 -24410 -75299 -24366
rect -75255 -24410 -71799 -24366
rect -87194 -24466 -71799 -24410
rect -87194 -24510 -82799 -24466
rect -82755 -24510 -82699 -24466
rect -82655 -24510 -82599 -24466
rect -82555 -24510 -82499 -24466
rect -82455 -24510 -82399 -24466
rect -82355 -24510 -82299 -24466
rect -82255 -24510 -82199 -24466
rect -82155 -24510 -82099 -24466
rect -82055 -24510 -81999 -24466
rect -81955 -24510 -81899 -24466
rect -81855 -24510 -81799 -24466
rect -81755 -24510 -81699 -24466
rect -81655 -24510 -81599 -24466
rect -81555 -24510 -81499 -24466
rect -81455 -24510 -81399 -24466
rect -81355 -24510 -81299 -24466
rect -81255 -24510 -80799 -24466
rect -80755 -24510 -80699 -24466
rect -80655 -24510 -80599 -24466
rect -80555 -24510 -80499 -24466
rect -80455 -24510 -80399 -24466
rect -80355 -24510 -80299 -24466
rect -80255 -24510 -80199 -24466
rect -80155 -24510 -80099 -24466
rect -80055 -24510 -79999 -24466
rect -79955 -24510 -79899 -24466
rect -79855 -24510 -79799 -24466
rect -79755 -24510 -79699 -24466
rect -79655 -24510 -79599 -24466
rect -79555 -24510 -79499 -24466
rect -79455 -24510 -79399 -24466
rect -79355 -24510 -79299 -24466
rect -79255 -24510 -78799 -24466
rect -78755 -24510 -78699 -24466
rect -78655 -24510 -78599 -24466
rect -78555 -24510 -78499 -24466
rect -78455 -24510 -78399 -24466
rect -78355 -24510 -78299 -24466
rect -78255 -24510 -78199 -24466
rect -78155 -24510 -78099 -24466
rect -78055 -24510 -77999 -24466
rect -77955 -24510 -77899 -24466
rect -77855 -24510 -77799 -24466
rect -77755 -24510 -77699 -24466
rect -77655 -24510 -77599 -24466
rect -77555 -24510 -77499 -24466
rect -77455 -24510 -77399 -24466
rect -77355 -24510 -77299 -24466
rect -77255 -24510 -76799 -24466
rect -76755 -24510 -76699 -24466
rect -76655 -24510 -76599 -24466
rect -76555 -24510 -76499 -24466
rect -76455 -24510 -76399 -24466
rect -76355 -24510 -76299 -24466
rect -76255 -24510 -76199 -24466
rect -76155 -24510 -76099 -24466
rect -76055 -24510 -75999 -24466
rect -75955 -24510 -75899 -24466
rect -75855 -24510 -75799 -24466
rect -75755 -24510 -75699 -24466
rect -75655 -24510 -75599 -24466
rect -75555 -24510 -75499 -24466
rect -75455 -24510 -75399 -24466
rect -75355 -24510 -75299 -24466
rect -75255 -24510 -71799 -24466
rect -87194 -24566 -71799 -24510
rect -87194 -24610 -82799 -24566
rect -82755 -24610 -82699 -24566
rect -82655 -24610 -82599 -24566
rect -82555 -24610 -82499 -24566
rect -82455 -24610 -82399 -24566
rect -82355 -24610 -82299 -24566
rect -82255 -24610 -82199 -24566
rect -82155 -24610 -82099 -24566
rect -82055 -24610 -81999 -24566
rect -81955 -24610 -81899 -24566
rect -81855 -24610 -81799 -24566
rect -81755 -24610 -81699 -24566
rect -81655 -24610 -81599 -24566
rect -81555 -24610 -81499 -24566
rect -81455 -24610 -81399 -24566
rect -81355 -24610 -81299 -24566
rect -81255 -24610 -80799 -24566
rect -80755 -24610 -80699 -24566
rect -80655 -24610 -80599 -24566
rect -80555 -24610 -80499 -24566
rect -80455 -24610 -80399 -24566
rect -80355 -24610 -80299 -24566
rect -80255 -24610 -80199 -24566
rect -80155 -24610 -80099 -24566
rect -80055 -24610 -79999 -24566
rect -79955 -24610 -79899 -24566
rect -79855 -24610 -79799 -24566
rect -79755 -24610 -79699 -24566
rect -79655 -24610 -79599 -24566
rect -79555 -24610 -79499 -24566
rect -79455 -24610 -79399 -24566
rect -79355 -24610 -79299 -24566
rect -79255 -24610 -78799 -24566
rect -78755 -24610 -78699 -24566
rect -78655 -24610 -78599 -24566
rect -78555 -24610 -78499 -24566
rect -78455 -24610 -78399 -24566
rect -78355 -24610 -78299 -24566
rect -78255 -24610 -78199 -24566
rect -78155 -24610 -78099 -24566
rect -78055 -24610 -77999 -24566
rect -77955 -24610 -77899 -24566
rect -77855 -24610 -77799 -24566
rect -77755 -24610 -77699 -24566
rect -77655 -24610 -77599 -24566
rect -77555 -24610 -77499 -24566
rect -77455 -24610 -77399 -24566
rect -77355 -24610 -77299 -24566
rect -77255 -24610 -76799 -24566
rect -76755 -24610 -76699 -24566
rect -76655 -24610 -76599 -24566
rect -76555 -24610 -76499 -24566
rect -76455 -24610 -76399 -24566
rect -76355 -24610 -76299 -24566
rect -76255 -24610 -76199 -24566
rect -76155 -24610 -76099 -24566
rect -76055 -24610 -75999 -24566
rect -75955 -24610 -75899 -24566
rect -75855 -24610 -75799 -24566
rect -75755 -24610 -75699 -24566
rect -75655 -24610 -75599 -24566
rect -75555 -24610 -75499 -24566
rect -75455 -24610 -75399 -24566
rect -75355 -24610 -75299 -24566
rect -75255 -24610 -71799 -24566
rect -87194 -24666 -71799 -24610
rect -87194 -24710 -82799 -24666
rect -82755 -24710 -82699 -24666
rect -82655 -24710 -82599 -24666
rect -82555 -24710 -82499 -24666
rect -82455 -24710 -82399 -24666
rect -82355 -24710 -82299 -24666
rect -82255 -24710 -82199 -24666
rect -82155 -24710 -82099 -24666
rect -82055 -24710 -81999 -24666
rect -81955 -24710 -81899 -24666
rect -81855 -24710 -81799 -24666
rect -81755 -24710 -81699 -24666
rect -81655 -24710 -81599 -24666
rect -81555 -24710 -81499 -24666
rect -81455 -24710 -81399 -24666
rect -81355 -24710 -81299 -24666
rect -81255 -24710 -80799 -24666
rect -80755 -24710 -80699 -24666
rect -80655 -24710 -80599 -24666
rect -80555 -24710 -80499 -24666
rect -80455 -24710 -80399 -24666
rect -80355 -24710 -80299 -24666
rect -80255 -24710 -80199 -24666
rect -80155 -24710 -80099 -24666
rect -80055 -24710 -79999 -24666
rect -79955 -24710 -79899 -24666
rect -79855 -24710 -79799 -24666
rect -79755 -24710 -79699 -24666
rect -79655 -24710 -79599 -24666
rect -79555 -24710 -79499 -24666
rect -79455 -24710 -79399 -24666
rect -79355 -24710 -79299 -24666
rect -79255 -24710 -78799 -24666
rect -78755 -24710 -78699 -24666
rect -78655 -24710 -78599 -24666
rect -78555 -24710 -78499 -24666
rect -78455 -24710 -78399 -24666
rect -78355 -24710 -78299 -24666
rect -78255 -24710 -78199 -24666
rect -78155 -24710 -78099 -24666
rect -78055 -24710 -77999 -24666
rect -77955 -24710 -77899 -24666
rect -77855 -24710 -77799 -24666
rect -77755 -24710 -77699 -24666
rect -77655 -24710 -77599 -24666
rect -77555 -24710 -77499 -24666
rect -77455 -24710 -77399 -24666
rect -77355 -24710 -77299 -24666
rect -77255 -24710 -76799 -24666
rect -76755 -24710 -76699 -24666
rect -76655 -24710 -76599 -24666
rect -76555 -24710 -76499 -24666
rect -76455 -24710 -76399 -24666
rect -76355 -24710 -76299 -24666
rect -76255 -24710 -76199 -24666
rect -76155 -24710 -76099 -24666
rect -76055 -24710 -75999 -24666
rect -75955 -24710 -75899 -24666
rect -75855 -24710 -75799 -24666
rect -75755 -24710 -75699 -24666
rect -75655 -24710 -75599 -24666
rect -75555 -24710 -75499 -24666
rect -75455 -24710 -75399 -24666
rect -75355 -24710 -75299 -24666
rect -75255 -24710 -71799 -24666
rect -87194 -24766 -71799 -24710
rect -87194 -24810 -82799 -24766
rect -82755 -24810 -82699 -24766
rect -82655 -24810 -82599 -24766
rect -82555 -24810 -82499 -24766
rect -82455 -24810 -82399 -24766
rect -82355 -24810 -82299 -24766
rect -82255 -24810 -82199 -24766
rect -82155 -24810 -82099 -24766
rect -82055 -24810 -81999 -24766
rect -81955 -24810 -81899 -24766
rect -81855 -24810 -81799 -24766
rect -81755 -24810 -81699 -24766
rect -81655 -24810 -81599 -24766
rect -81555 -24810 -81499 -24766
rect -81455 -24810 -81399 -24766
rect -81355 -24810 -81299 -24766
rect -81255 -24810 -80799 -24766
rect -80755 -24810 -80699 -24766
rect -80655 -24810 -80599 -24766
rect -80555 -24810 -80499 -24766
rect -80455 -24810 -80399 -24766
rect -80355 -24810 -80299 -24766
rect -80255 -24810 -80199 -24766
rect -80155 -24810 -80099 -24766
rect -80055 -24810 -79999 -24766
rect -79955 -24810 -79899 -24766
rect -79855 -24810 -79799 -24766
rect -79755 -24810 -79699 -24766
rect -79655 -24810 -79599 -24766
rect -79555 -24810 -79499 -24766
rect -79455 -24810 -79399 -24766
rect -79355 -24810 -79299 -24766
rect -79255 -24810 -78799 -24766
rect -78755 -24810 -78699 -24766
rect -78655 -24810 -78599 -24766
rect -78555 -24810 -78499 -24766
rect -78455 -24810 -78399 -24766
rect -78355 -24810 -78299 -24766
rect -78255 -24810 -78199 -24766
rect -78155 -24810 -78099 -24766
rect -78055 -24810 -77999 -24766
rect -77955 -24810 -77899 -24766
rect -77855 -24810 -77799 -24766
rect -77755 -24810 -77699 -24766
rect -77655 -24810 -77599 -24766
rect -77555 -24810 -77499 -24766
rect -77455 -24810 -77399 -24766
rect -77355 -24810 -77299 -24766
rect -77255 -24810 -76799 -24766
rect -76755 -24810 -76699 -24766
rect -76655 -24810 -76599 -24766
rect -76555 -24810 -76499 -24766
rect -76455 -24810 -76399 -24766
rect -76355 -24810 -76299 -24766
rect -76255 -24810 -76199 -24766
rect -76155 -24810 -76099 -24766
rect -76055 -24810 -75999 -24766
rect -75955 -24810 -75899 -24766
rect -75855 -24810 -75799 -24766
rect -75755 -24810 -75699 -24766
rect -75655 -24810 -75599 -24766
rect -75555 -24810 -75499 -24766
rect -75455 -24810 -75399 -24766
rect -75355 -24810 -75299 -24766
rect -75255 -24810 -71799 -24766
rect -87194 -24866 -71799 -24810
rect -87194 -24910 -82799 -24866
rect -82755 -24910 -82699 -24866
rect -82655 -24910 -82599 -24866
rect -82555 -24910 -82499 -24866
rect -82455 -24910 -82399 -24866
rect -82355 -24910 -82299 -24866
rect -82255 -24910 -82199 -24866
rect -82155 -24910 -82099 -24866
rect -82055 -24910 -81999 -24866
rect -81955 -24910 -81899 -24866
rect -81855 -24910 -81799 -24866
rect -81755 -24910 -81699 -24866
rect -81655 -24910 -81599 -24866
rect -81555 -24910 -81499 -24866
rect -81455 -24910 -81399 -24866
rect -81355 -24910 -81299 -24866
rect -81255 -24910 -80799 -24866
rect -80755 -24910 -80699 -24866
rect -80655 -24910 -80599 -24866
rect -80555 -24910 -80499 -24866
rect -80455 -24910 -80399 -24866
rect -80355 -24910 -80299 -24866
rect -80255 -24910 -80199 -24866
rect -80155 -24910 -80099 -24866
rect -80055 -24910 -79999 -24866
rect -79955 -24910 -79899 -24866
rect -79855 -24910 -79799 -24866
rect -79755 -24910 -79699 -24866
rect -79655 -24910 -79599 -24866
rect -79555 -24910 -79499 -24866
rect -79455 -24910 -79399 -24866
rect -79355 -24910 -79299 -24866
rect -79255 -24910 -78799 -24866
rect -78755 -24910 -78699 -24866
rect -78655 -24910 -78599 -24866
rect -78555 -24910 -78499 -24866
rect -78455 -24910 -78399 -24866
rect -78355 -24910 -78299 -24866
rect -78255 -24910 -78199 -24866
rect -78155 -24910 -78099 -24866
rect -78055 -24910 -77999 -24866
rect -77955 -24910 -77899 -24866
rect -77855 -24910 -77799 -24866
rect -77755 -24910 -77699 -24866
rect -77655 -24910 -77599 -24866
rect -77555 -24910 -77499 -24866
rect -77455 -24910 -77399 -24866
rect -77355 -24910 -77299 -24866
rect -77255 -24910 -76799 -24866
rect -76755 -24910 -76699 -24866
rect -76655 -24910 -76599 -24866
rect -76555 -24910 -76499 -24866
rect -76455 -24910 -76399 -24866
rect -76355 -24910 -76299 -24866
rect -76255 -24910 -76199 -24866
rect -76155 -24910 -76099 -24866
rect -76055 -24910 -75999 -24866
rect -75955 -24910 -75899 -24866
rect -75855 -24910 -75799 -24866
rect -75755 -24910 -75699 -24866
rect -75655 -24910 -75599 -24866
rect -75555 -24910 -75499 -24866
rect -75455 -24910 -75399 -24866
rect -75355 -24910 -75299 -24866
rect -75255 -24910 -71799 -24866
rect -87194 -24966 -71799 -24910
rect -87194 -25010 -82799 -24966
rect -82755 -25010 -82699 -24966
rect -82655 -25010 -82599 -24966
rect -82555 -25010 -82499 -24966
rect -82455 -25010 -82399 -24966
rect -82355 -25010 -82299 -24966
rect -82255 -25010 -82199 -24966
rect -82155 -25010 -82099 -24966
rect -82055 -25010 -81999 -24966
rect -81955 -25010 -81899 -24966
rect -81855 -25010 -81799 -24966
rect -81755 -25010 -81699 -24966
rect -81655 -25010 -81599 -24966
rect -81555 -25010 -81499 -24966
rect -81455 -25010 -81399 -24966
rect -81355 -25010 -81299 -24966
rect -81255 -25010 -80799 -24966
rect -80755 -25010 -80699 -24966
rect -80655 -25010 -80599 -24966
rect -80555 -25010 -80499 -24966
rect -80455 -25010 -80399 -24966
rect -80355 -25010 -80299 -24966
rect -80255 -25010 -80199 -24966
rect -80155 -25010 -80099 -24966
rect -80055 -25010 -79999 -24966
rect -79955 -25010 -79899 -24966
rect -79855 -25010 -79799 -24966
rect -79755 -25010 -79699 -24966
rect -79655 -25010 -79599 -24966
rect -79555 -25010 -79499 -24966
rect -79455 -25010 -79399 -24966
rect -79355 -25010 -79299 -24966
rect -79255 -25010 -78799 -24966
rect -78755 -25010 -78699 -24966
rect -78655 -25010 -78599 -24966
rect -78555 -25010 -78499 -24966
rect -78455 -25010 -78399 -24966
rect -78355 -25010 -78299 -24966
rect -78255 -25010 -78199 -24966
rect -78155 -25010 -78099 -24966
rect -78055 -25010 -77999 -24966
rect -77955 -25010 -77899 -24966
rect -77855 -25010 -77799 -24966
rect -77755 -25010 -77699 -24966
rect -77655 -25010 -77599 -24966
rect -77555 -25010 -77499 -24966
rect -77455 -25010 -77399 -24966
rect -77355 -25010 -77299 -24966
rect -77255 -25010 -76799 -24966
rect -76755 -25010 -76699 -24966
rect -76655 -25010 -76599 -24966
rect -76555 -25010 -76499 -24966
rect -76455 -25010 -76399 -24966
rect -76355 -25010 -76299 -24966
rect -76255 -25010 -76199 -24966
rect -76155 -25010 -76099 -24966
rect -76055 -25010 -75999 -24966
rect -75955 -25010 -75899 -24966
rect -75855 -25010 -75799 -24966
rect -75755 -25010 -75699 -24966
rect -75655 -25010 -75599 -24966
rect -75555 -25010 -75499 -24966
rect -75455 -25010 -75399 -24966
rect -75355 -25010 -75299 -24966
rect -75255 -25010 -71799 -24966
rect -87194 -25066 -71799 -25010
rect -87194 -25110 -82799 -25066
rect -82755 -25110 -82699 -25066
rect -82655 -25110 -82599 -25066
rect -82555 -25110 -82499 -25066
rect -82455 -25110 -82399 -25066
rect -82355 -25110 -82299 -25066
rect -82255 -25110 -82199 -25066
rect -82155 -25110 -82099 -25066
rect -82055 -25110 -81999 -25066
rect -81955 -25110 -81899 -25066
rect -81855 -25110 -81799 -25066
rect -81755 -25110 -81699 -25066
rect -81655 -25110 -81599 -25066
rect -81555 -25110 -81499 -25066
rect -81455 -25110 -81399 -25066
rect -81355 -25110 -81299 -25066
rect -81255 -25110 -80799 -25066
rect -80755 -25110 -80699 -25066
rect -80655 -25110 -80599 -25066
rect -80555 -25110 -80499 -25066
rect -80455 -25110 -80399 -25066
rect -80355 -25110 -80299 -25066
rect -80255 -25110 -80199 -25066
rect -80155 -25110 -80099 -25066
rect -80055 -25110 -79999 -25066
rect -79955 -25110 -79899 -25066
rect -79855 -25110 -79799 -25066
rect -79755 -25110 -79699 -25066
rect -79655 -25110 -79599 -25066
rect -79555 -25110 -79499 -25066
rect -79455 -25110 -79399 -25066
rect -79355 -25110 -79299 -25066
rect -79255 -25110 -78799 -25066
rect -78755 -25110 -78699 -25066
rect -78655 -25110 -78599 -25066
rect -78555 -25110 -78499 -25066
rect -78455 -25110 -78399 -25066
rect -78355 -25110 -78299 -25066
rect -78255 -25110 -78199 -25066
rect -78155 -25110 -78099 -25066
rect -78055 -25110 -77999 -25066
rect -77955 -25110 -77899 -25066
rect -77855 -25110 -77799 -25066
rect -77755 -25110 -77699 -25066
rect -77655 -25110 -77599 -25066
rect -77555 -25110 -77499 -25066
rect -77455 -25110 -77399 -25066
rect -77355 -25110 -77299 -25066
rect -77255 -25110 -76799 -25066
rect -76755 -25110 -76699 -25066
rect -76655 -25110 -76599 -25066
rect -76555 -25110 -76499 -25066
rect -76455 -25110 -76399 -25066
rect -76355 -25110 -76299 -25066
rect -76255 -25110 -76199 -25066
rect -76155 -25110 -76099 -25066
rect -76055 -25110 -75999 -25066
rect -75955 -25110 -75899 -25066
rect -75855 -25110 -75799 -25066
rect -75755 -25110 -75699 -25066
rect -75655 -25110 -75599 -25066
rect -75555 -25110 -75499 -25066
rect -75455 -25110 -75399 -25066
rect -75355 -25110 -75299 -25066
rect -75255 -25110 -71799 -25066
rect -87194 -25166 -71799 -25110
rect -87194 -25210 -82799 -25166
rect -82755 -25210 -82699 -25166
rect -82655 -25210 -82599 -25166
rect -82555 -25210 -82499 -25166
rect -82455 -25210 -82399 -25166
rect -82355 -25210 -82299 -25166
rect -82255 -25210 -82199 -25166
rect -82155 -25210 -82099 -25166
rect -82055 -25210 -81999 -25166
rect -81955 -25210 -81899 -25166
rect -81855 -25210 -81799 -25166
rect -81755 -25210 -81699 -25166
rect -81655 -25210 -81599 -25166
rect -81555 -25210 -81499 -25166
rect -81455 -25210 -81399 -25166
rect -81355 -25210 -81299 -25166
rect -81255 -25210 -80799 -25166
rect -80755 -25210 -80699 -25166
rect -80655 -25210 -80599 -25166
rect -80555 -25210 -80499 -25166
rect -80455 -25210 -80399 -25166
rect -80355 -25210 -80299 -25166
rect -80255 -25210 -80199 -25166
rect -80155 -25210 -80099 -25166
rect -80055 -25210 -79999 -25166
rect -79955 -25210 -79899 -25166
rect -79855 -25210 -79799 -25166
rect -79755 -25210 -79699 -25166
rect -79655 -25210 -79599 -25166
rect -79555 -25210 -79499 -25166
rect -79455 -25210 -79399 -25166
rect -79355 -25210 -79299 -25166
rect -79255 -25210 -78799 -25166
rect -78755 -25210 -78699 -25166
rect -78655 -25210 -78599 -25166
rect -78555 -25210 -78499 -25166
rect -78455 -25210 -78399 -25166
rect -78355 -25210 -78299 -25166
rect -78255 -25210 -78199 -25166
rect -78155 -25210 -78099 -25166
rect -78055 -25210 -77999 -25166
rect -77955 -25210 -77899 -25166
rect -77855 -25210 -77799 -25166
rect -77755 -25210 -77699 -25166
rect -77655 -25210 -77599 -25166
rect -77555 -25210 -77499 -25166
rect -77455 -25210 -77399 -25166
rect -77355 -25210 -77299 -25166
rect -77255 -25210 -76799 -25166
rect -76755 -25210 -76699 -25166
rect -76655 -25210 -76599 -25166
rect -76555 -25210 -76499 -25166
rect -76455 -25210 -76399 -25166
rect -76355 -25210 -76299 -25166
rect -76255 -25210 -76199 -25166
rect -76155 -25210 -76099 -25166
rect -76055 -25210 -75999 -25166
rect -75955 -25210 -75899 -25166
rect -75855 -25210 -75799 -25166
rect -75755 -25210 -75699 -25166
rect -75655 -25210 -75599 -25166
rect -75555 -25210 -75499 -25166
rect -75455 -25210 -75399 -25166
rect -75355 -25210 -75299 -25166
rect -75255 -25210 -71799 -25166
rect -87194 -25266 -71799 -25210
rect -87194 -25310 -82799 -25266
rect -82755 -25310 -82699 -25266
rect -82655 -25310 -82599 -25266
rect -82555 -25310 -82499 -25266
rect -82455 -25310 -82399 -25266
rect -82355 -25310 -82299 -25266
rect -82255 -25310 -82199 -25266
rect -82155 -25310 -82099 -25266
rect -82055 -25310 -81999 -25266
rect -81955 -25310 -81899 -25266
rect -81855 -25310 -81799 -25266
rect -81755 -25310 -81699 -25266
rect -81655 -25310 -81599 -25266
rect -81555 -25310 -81499 -25266
rect -81455 -25310 -81399 -25266
rect -81355 -25310 -81299 -25266
rect -81255 -25310 -80799 -25266
rect -80755 -25310 -80699 -25266
rect -80655 -25310 -80599 -25266
rect -80555 -25310 -80499 -25266
rect -80455 -25310 -80399 -25266
rect -80355 -25310 -80299 -25266
rect -80255 -25310 -80199 -25266
rect -80155 -25310 -80099 -25266
rect -80055 -25310 -79999 -25266
rect -79955 -25310 -79899 -25266
rect -79855 -25310 -79799 -25266
rect -79755 -25310 -79699 -25266
rect -79655 -25310 -79599 -25266
rect -79555 -25310 -79499 -25266
rect -79455 -25310 -79399 -25266
rect -79355 -25310 -79299 -25266
rect -79255 -25310 -78799 -25266
rect -78755 -25310 -78699 -25266
rect -78655 -25310 -78599 -25266
rect -78555 -25310 -78499 -25266
rect -78455 -25310 -78399 -25266
rect -78355 -25310 -78299 -25266
rect -78255 -25310 -78199 -25266
rect -78155 -25310 -78099 -25266
rect -78055 -25310 -77999 -25266
rect -77955 -25310 -77899 -25266
rect -77855 -25310 -77799 -25266
rect -77755 -25310 -77699 -25266
rect -77655 -25310 -77599 -25266
rect -77555 -25310 -77499 -25266
rect -77455 -25310 -77399 -25266
rect -77355 -25310 -77299 -25266
rect -77255 -25310 -76799 -25266
rect -76755 -25310 -76699 -25266
rect -76655 -25310 -76599 -25266
rect -76555 -25310 -76499 -25266
rect -76455 -25310 -76399 -25266
rect -76355 -25310 -76299 -25266
rect -76255 -25310 -76199 -25266
rect -76155 -25310 -76099 -25266
rect -76055 -25310 -75999 -25266
rect -75955 -25310 -75899 -25266
rect -75855 -25310 -75799 -25266
rect -75755 -25310 -75699 -25266
rect -75655 -25310 -75599 -25266
rect -75555 -25310 -75499 -25266
rect -75455 -25310 -75399 -25266
rect -75355 -25310 -75299 -25266
rect -75255 -25310 -71799 -25266
rect -87194 -25366 -71799 -25310
rect -87194 -25410 -82799 -25366
rect -82755 -25410 -82699 -25366
rect -82655 -25410 -82599 -25366
rect -82555 -25410 -82499 -25366
rect -82455 -25410 -82399 -25366
rect -82355 -25410 -82299 -25366
rect -82255 -25410 -82199 -25366
rect -82155 -25410 -82099 -25366
rect -82055 -25410 -81999 -25366
rect -81955 -25410 -81899 -25366
rect -81855 -25410 -81799 -25366
rect -81755 -25410 -81699 -25366
rect -81655 -25410 -81599 -25366
rect -81555 -25410 -81499 -25366
rect -81455 -25410 -81399 -25366
rect -81355 -25410 -81299 -25366
rect -81255 -25410 -80799 -25366
rect -80755 -25410 -80699 -25366
rect -80655 -25410 -80599 -25366
rect -80555 -25410 -80499 -25366
rect -80455 -25410 -80399 -25366
rect -80355 -25410 -80299 -25366
rect -80255 -25410 -80199 -25366
rect -80155 -25410 -80099 -25366
rect -80055 -25410 -79999 -25366
rect -79955 -25410 -79899 -25366
rect -79855 -25410 -79799 -25366
rect -79755 -25410 -79699 -25366
rect -79655 -25410 -79599 -25366
rect -79555 -25410 -79499 -25366
rect -79455 -25410 -79399 -25366
rect -79355 -25410 -79299 -25366
rect -79255 -25410 -78799 -25366
rect -78755 -25410 -78699 -25366
rect -78655 -25410 -78599 -25366
rect -78555 -25410 -78499 -25366
rect -78455 -25410 -78399 -25366
rect -78355 -25410 -78299 -25366
rect -78255 -25410 -78199 -25366
rect -78155 -25410 -78099 -25366
rect -78055 -25410 -77999 -25366
rect -77955 -25410 -77899 -25366
rect -77855 -25410 -77799 -25366
rect -77755 -25410 -77699 -25366
rect -77655 -25410 -77599 -25366
rect -77555 -25410 -77499 -25366
rect -77455 -25410 -77399 -25366
rect -77355 -25410 -77299 -25366
rect -77255 -25410 -76799 -25366
rect -76755 -25410 -76699 -25366
rect -76655 -25410 -76599 -25366
rect -76555 -25410 -76499 -25366
rect -76455 -25410 -76399 -25366
rect -76355 -25410 -76299 -25366
rect -76255 -25410 -76199 -25366
rect -76155 -25410 -76099 -25366
rect -76055 -25410 -75999 -25366
rect -75955 -25410 -75899 -25366
rect -75855 -25410 -75799 -25366
rect -75755 -25410 -75699 -25366
rect -75655 -25410 -75599 -25366
rect -75555 -25410 -75499 -25366
rect -75455 -25410 -75399 -25366
rect -75355 -25410 -75299 -25366
rect -75255 -25410 -71799 -25366
rect -87194 -25466 -71799 -25410
rect -87194 -25510 -82799 -25466
rect -82755 -25510 -82699 -25466
rect -82655 -25510 -82599 -25466
rect -82555 -25510 -82499 -25466
rect -82455 -25510 -82399 -25466
rect -82355 -25510 -82299 -25466
rect -82255 -25510 -82199 -25466
rect -82155 -25510 -82099 -25466
rect -82055 -25510 -81999 -25466
rect -81955 -25510 -81899 -25466
rect -81855 -25510 -81799 -25466
rect -81755 -25510 -81699 -25466
rect -81655 -25510 -81599 -25466
rect -81555 -25510 -81499 -25466
rect -81455 -25510 -81399 -25466
rect -81355 -25510 -81299 -25466
rect -81255 -25510 -80799 -25466
rect -80755 -25510 -80699 -25466
rect -80655 -25510 -80599 -25466
rect -80555 -25510 -80499 -25466
rect -80455 -25510 -80399 -25466
rect -80355 -25510 -80299 -25466
rect -80255 -25510 -80199 -25466
rect -80155 -25510 -80099 -25466
rect -80055 -25510 -79999 -25466
rect -79955 -25510 -79899 -25466
rect -79855 -25510 -79799 -25466
rect -79755 -25510 -79699 -25466
rect -79655 -25510 -79599 -25466
rect -79555 -25510 -79499 -25466
rect -79455 -25510 -79399 -25466
rect -79355 -25510 -79299 -25466
rect -79255 -25510 -78799 -25466
rect -78755 -25510 -78699 -25466
rect -78655 -25510 -78599 -25466
rect -78555 -25510 -78499 -25466
rect -78455 -25510 -78399 -25466
rect -78355 -25510 -78299 -25466
rect -78255 -25510 -78199 -25466
rect -78155 -25510 -78099 -25466
rect -78055 -25510 -77999 -25466
rect -77955 -25510 -77899 -25466
rect -77855 -25510 -77799 -25466
rect -77755 -25510 -77699 -25466
rect -77655 -25510 -77599 -25466
rect -77555 -25510 -77499 -25466
rect -77455 -25510 -77399 -25466
rect -77355 -25510 -77299 -25466
rect -77255 -25510 -76799 -25466
rect -76755 -25510 -76699 -25466
rect -76655 -25510 -76599 -25466
rect -76555 -25510 -76499 -25466
rect -76455 -25510 -76399 -25466
rect -76355 -25510 -76299 -25466
rect -76255 -25510 -76199 -25466
rect -76155 -25510 -76099 -25466
rect -76055 -25510 -75999 -25466
rect -75955 -25510 -75899 -25466
rect -75855 -25510 -75799 -25466
rect -75755 -25510 -75699 -25466
rect -75655 -25510 -75599 -25466
rect -75555 -25510 -75499 -25466
rect -75455 -25510 -75399 -25466
rect -75355 -25510 -75299 -25466
rect -75255 -25510 -71799 -25466
rect -87194 -25566 -71799 -25510
rect -87194 -25610 -82799 -25566
rect -82755 -25610 -82699 -25566
rect -82655 -25610 -82599 -25566
rect -82555 -25610 -82499 -25566
rect -82455 -25610 -82399 -25566
rect -82355 -25610 -82299 -25566
rect -82255 -25610 -82199 -25566
rect -82155 -25610 -82099 -25566
rect -82055 -25610 -81999 -25566
rect -81955 -25610 -81899 -25566
rect -81855 -25610 -81799 -25566
rect -81755 -25610 -81699 -25566
rect -81655 -25610 -81599 -25566
rect -81555 -25610 -81499 -25566
rect -81455 -25610 -81399 -25566
rect -81355 -25610 -81299 -25566
rect -81255 -25610 -80799 -25566
rect -80755 -25610 -80699 -25566
rect -80655 -25610 -80599 -25566
rect -80555 -25610 -80499 -25566
rect -80455 -25610 -80399 -25566
rect -80355 -25610 -80299 -25566
rect -80255 -25610 -80199 -25566
rect -80155 -25610 -80099 -25566
rect -80055 -25610 -79999 -25566
rect -79955 -25610 -79899 -25566
rect -79855 -25610 -79799 -25566
rect -79755 -25610 -79699 -25566
rect -79655 -25610 -79599 -25566
rect -79555 -25610 -79499 -25566
rect -79455 -25610 -79399 -25566
rect -79355 -25610 -79299 -25566
rect -79255 -25610 -78799 -25566
rect -78755 -25610 -78699 -25566
rect -78655 -25610 -78599 -25566
rect -78555 -25610 -78499 -25566
rect -78455 -25610 -78399 -25566
rect -78355 -25610 -78299 -25566
rect -78255 -25610 -78199 -25566
rect -78155 -25610 -78099 -25566
rect -78055 -25610 -77999 -25566
rect -77955 -25610 -77899 -25566
rect -77855 -25610 -77799 -25566
rect -77755 -25610 -77699 -25566
rect -77655 -25610 -77599 -25566
rect -77555 -25610 -77499 -25566
rect -77455 -25610 -77399 -25566
rect -77355 -25610 -77299 -25566
rect -77255 -25610 -76799 -25566
rect -76755 -25610 -76699 -25566
rect -76655 -25610 -76599 -25566
rect -76555 -25610 -76499 -25566
rect -76455 -25610 -76399 -25566
rect -76355 -25610 -76299 -25566
rect -76255 -25610 -76199 -25566
rect -76155 -25610 -76099 -25566
rect -76055 -25610 -75999 -25566
rect -75955 -25610 -75899 -25566
rect -75855 -25610 -75799 -25566
rect -75755 -25610 -75699 -25566
rect -75655 -25610 -75599 -25566
rect -75555 -25610 -75499 -25566
rect -75455 -25610 -75399 -25566
rect -75355 -25610 -75299 -25566
rect -75255 -25610 -71799 -25566
rect -87194 -25666 -71799 -25610
rect -87194 -25710 -82799 -25666
rect -82755 -25710 -82699 -25666
rect -82655 -25710 -82599 -25666
rect -82555 -25710 -82499 -25666
rect -82455 -25710 -82399 -25666
rect -82355 -25710 -82299 -25666
rect -82255 -25710 -82199 -25666
rect -82155 -25710 -82099 -25666
rect -82055 -25710 -81999 -25666
rect -81955 -25710 -81899 -25666
rect -81855 -25710 -81799 -25666
rect -81755 -25710 -81699 -25666
rect -81655 -25710 -81599 -25666
rect -81555 -25710 -81499 -25666
rect -81455 -25710 -81399 -25666
rect -81355 -25710 -81299 -25666
rect -81255 -25710 -80799 -25666
rect -80755 -25710 -80699 -25666
rect -80655 -25710 -80599 -25666
rect -80555 -25710 -80499 -25666
rect -80455 -25710 -80399 -25666
rect -80355 -25710 -80299 -25666
rect -80255 -25710 -80199 -25666
rect -80155 -25710 -80099 -25666
rect -80055 -25710 -79999 -25666
rect -79955 -25710 -79899 -25666
rect -79855 -25710 -79799 -25666
rect -79755 -25710 -79699 -25666
rect -79655 -25710 -79599 -25666
rect -79555 -25710 -79499 -25666
rect -79455 -25710 -79399 -25666
rect -79355 -25710 -79299 -25666
rect -79255 -25710 -78799 -25666
rect -78755 -25710 -78699 -25666
rect -78655 -25710 -78599 -25666
rect -78555 -25710 -78499 -25666
rect -78455 -25710 -78399 -25666
rect -78355 -25710 -78299 -25666
rect -78255 -25710 -78199 -25666
rect -78155 -25710 -78099 -25666
rect -78055 -25710 -77999 -25666
rect -77955 -25710 -77899 -25666
rect -77855 -25710 -77799 -25666
rect -77755 -25710 -77699 -25666
rect -77655 -25710 -77599 -25666
rect -77555 -25710 -77499 -25666
rect -77455 -25710 -77399 -25666
rect -77355 -25710 -77299 -25666
rect -77255 -25710 -76799 -25666
rect -76755 -25710 -76699 -25666
rect -76655 -25710 -76599 -25666
rect -76555 -25710 -76499 -25666
rect -76455 -25710 -76399 -25666
rect -76355 -25710 -76299 -25666
rect -76255 -25710 -76199 -25666
rect -76155 -25710 -76099 -25666
rect -76055 -25710 -75999 -25666
rect -75955 -25710 -75899 -25666
rect -75855 -25710 -75799 -25666
rect -75755 -25710 -75699 -25666
rect -75655 -25710 -75599 -25666
rect -75555 -25710 -75499 -25666
rect -75455 -25710 -75399 -25666
rect -75355 -25710 -75299 -25666
rect -75255 -25710 -71799 -25666
rect -87194 -25766 -71799 -25710
rect -87194 -25810 -82799 -25766
rect -82755 -25810 -82699 -25766
rect -82655 -25810 -82599 -25766
rect -82555 -25810 -82499 -25766
rect -82455 -25810 -82399 -25766
rect -82355 -25810 -82299 -25766
rect -82255 -25810 -82199 -25766
rect -82155 -25810 -82099 -25766
rect -82055 -25810 -81999 -25766
rect -81955 -25810 -81899 -25766
rect -81855 -25810 -81799 -25766
rect -81755 -25810 -81699 -25766
rect -81655 -25810 -81599 -25766
rect -81555 -25810 -81499 -25766
rect -81455 -25810 -81399 -25766
rect -81355 -25810 -81299 -25766
rect -81255 -25810 -80799 -25766
rect -80755 -25810 -80699 -25766
rect -80655 -25810 -80599 -25766
rect -80555 -25810 -80499 -25766
rect -80455 -25810 -80399 -25766
rect -80355 -25810 -80299 -25766
rect -80255 -25810 -80199 -25766
rect -80155 -25810 -80099 -25766
rect -80055 -25810 -79999 -25766
rect -79955 -25810 -79899 -25766
rect -79855 -25810 -79799 -25766
rect -79755 -25810 -79699 -25766
rect -79655 -25810 -79599 -25766
rect -79555 -25810 -79499 -25766
rect -79455 -25810 -79399 -25766
rect -79355 -25810 -79299 -25766
rect -79255 -25810 -78799 -25766
rect -78755 -25810 -78699 -25766
rect -78655 -25810 -78599 -25766
rect -78555 -25810 -78499 -25766
rect -78455 -25810 -78399 -25766
rect -78355 -25810 -78299 -25766
rect -78255 -25810 -78199 -25766
rect -78155 -25810 -78099 -25766
rect -78055 -25810 -77999 -25766
rect -77955 -25810 -77899 -25766
rect -77855 -25810 -77799 -25766
rect -77755 -25810 -77699 -25766
rect -77655 -25810 -77599 -25766
rect -77555 -25810 -77499 -25766
rect -77455 -25810 -77399 -25766
rect -77355 -25810 -77299 -25766
rect -77255 -25810 -76799 -25766
rect -76755 -25810 -76699 -25766
rect -76655 -25810 -76599 -25766
rect -76555 -25810 -76499 -25766
rect -76455 -25810 -76399 -25766
rect -76355 -25810 -76299 -25766
rect -76255 -25810 -76199 -25766
rect -76155 -25810 -76099 -25766
rect -76055 -25810 -75999 -25766
rect -75955 -25810 -75899 -25766
rect -75855 -25810 -75799 -25766
rect -75755 -25810 -75699 -25766
rect -75655 -25810 -75599 -25766
rect -75555 -25810 -75499 -25766
rect -75455 -25810 -75399 -25766
rect -75355 -25810 -75299 -25766
rect -75255 -25810 -71799 -25766
rect -87194 -25866 -71799 -25810
rect -87194 -25910 -82799 -25866
rect -82755 -25910 -82699 -25866
rect -82655 -25910 -82599 -25866
rect -82555 -25910 -82499 -25866
rect -82455 -25910 -82399 -25866
rect -82355 -25910 -82299 -25866
rect -82255 -25910 -82199 -25866
rect -82155 -25910 -82099 -25866
rect -82055 -25910 -81999 -25866
rect -81955 -25910 -81899 -25866
rect -81855 -25910 -81799 -25866
rect -81755 -25910 -81699 -25866
rect -81655 -25910 -81599 -25866
rect -81555 -25910 -81499 -25866
rect -81455 -25910 -81399 -25866
rect -81355 -25910 -81299 -25866
rect -81255 -25910 -80799 -25866
rect -80755 -25910 -80699 -25866
rect -80655 -25910 -80599 -25866
rect -80555 -25910 -80499 -25866
rect -80455 -25910 -80399 -25866
rect -80355 -25910 -80299 -25866
rect -80255 -25910 -80199 -25866
rect -80155 -25910 -80099 -25866
rect -80055 -25910 -79999 -25866
rect -79955 -25910 -79899 -25866
rect -79855 -25910 -79799 -25866
rect -79755 -25910 -79699 -25866
rect -79655 -25910 -79599 -25866
rect -79555 -25910 -79499 -25866
rect -79455 -25910 -79399 -25866
rect -79355 -25910 -79299 -25866
rect -79255 -25910 -78799 -25866
rect -78755 -25910 -78699 -25866
rect -78655 -25910 -78599 -25866
rect -78555 -25910 -78499 -25866
rect -78455 -25910 -78399 -25866
rect -78355 -25910 -78299 -25866
rect -78255 -25910 -78199 -25866
rect -78155 -25910 -78099 -25866
rect -78055 -25910 -77999 -25866
rect -77955 -25910 -77899 -25866
rect -77855 -25910 -77799 -25866
rect -77755 -25910 -77699 -25866
rect -77655 -25910 -77599 -25866
rect -77555 -25910 -77499 -25866
rect -77455 -25910 -77399 -25866
rect -77355 -25910 -77299 -25866
rect -77255 -25910 -76799 -25866
rect -76755 -25910 -76699 -25866
rect -76655 -25910 -76599 -25866
rect -76555 -25910 -76499 -25866
rect -76455 -25910 -76399 -25866
rect -76355 -25910 -76299 -25866
rect -76255 -25910 -76199 -25866
rect -76155 -25910 -76099 -25866
rect -76055 -25910 -75999 -25866
rect -75955 -25910 -75899 -25866
rect -75855 -25910 -75799 -25866
rect -75755 -25910 -75699 -25866
rect -75655 -25910 -75599 -25866
rect -75555 -25910 -75499 -25866
rect -75455 -25910 -75399 -25866
rect -75355 -25910 -75299 -25866
rect -75255 -25910 -71799 -25866
rect -87194 -80459 -71799 -25910
rect -87194 -80503 -82968 -80459
rect -82924 -80503 -82868 -80459
rect -82824 -80503 -82768 -80459
rect -82724 -80503 -82668 -80459
rect -82624 -80503 -82568 -80459
rect -82524 -80503 -82468 -80459
rect -82424 -80503 -82368 -80459
rect -82324 -80503 -82268 -80459
rect -82224 -80503 -82168 -80459
rect -82124 -80503 -82068 -80459
rect -82024 -80503 -81968 -80459
rect -81924 -80503 -81868 -80459
rect -81824 -80503 -81768 -80459
rect -81724 -80503 -81668 -80459
rect -81624 -80503 -81568 -80459
rect -81524 -80503 -81468 -80459
rect -81424 -80503 -80968 -80459
rect -80924 -80503 -80868 -80459
rect -80824 -80503 -80768 -80459
rect -80724 -80503 -80668 -80459
rect -80624 -80503 -80568 -80459
rect -80524 -80503 -80468 -80459
rect -80424 -80503 -80368 -80459
rect -80324 -80503 -80268 -80459
rect -80224 -80503 -80168 -80459
rect -80124 -80503 -80068 -80459
rect -80024 -80503 -79968 -80459
rect -79924 -80503 -79868 -80459
rect -79824 -80503 -79768 -80459
rect -79724 -80503 -79668 -80459
rect -79624 -80503 -79568 -80459
rect -79524 -80503 -79468 -80459
rect -79424 -80503 -78968 -80459
rect -78924 -80503 -78868 -80459
rect -78824 -80503 -78768 -80459
rect -78724 -80503 -78668 -80459
rect -78624 -80503 -78568 -80459
rect -78524 -80503 -78468 -80459
rect -78424 -80503 -78368 -80459
rect -78324 -80503 -78268 -80459
rect -78224 -80503 -78168 -80459
rect -78124 -80503 -78068 -80459
rect -78024 -80503 -77968 -80459
rect -77924 -80503 -77868 -80459
rect -77824 -80503 -77768 -80459
rect -77724 -80503 -77668 -80459
rect -77624 -80503 -77568 -80459
rect -77524 -80503 -77468 -80459
rect -77424 -80503 -76968 -80459
rect -76924 -80503 -76868 -80459
rect -76824 -80503 -76768 -80459
rect -76724 -80503 -76668 -80459
rect -76624 -80503 -76568 -80459
rect -76524 -80503 -76468 -80459
rect -76424 -80503 -76368 -80459
rect -76324 -80503 -76268 -80459
rect -76224 -80503 -76168 -80459
rect -76124 -80503 -76068 -80459
rect -76024 -80503 -75968 -80459
rect -75924 -80503 -75868 -80459
rect -75824 -80503 -75768 -80459
rect -75724 -80503 -75668 -80459
rect -75624 -80503 -75568 -80459
rect -75524 -80503 -75468 -80459
rect -75424 -80503 -71799 -80459
rect -87194 -80559 -71799 -80503
rect -87194 -80603 -82968 -80559
rect -82924 -80603 -82868 -80559
rect -82824 -80603 -82768 -80559
rect -82724 -80603 -82668 -80559
rect -82624 -80603 -82568 -80559
rect -82524 -80603 -82468 -80559
rect -82424 -80603 -82368 -80559
rect -82324 -80603 -82268 -80559
rect -82224 -80603 -82168 -80559
rect -82124 -80603 -82068 -80559
rect -82024 -80603 -81968 -80559
rect -81924 -80603 -81868 -80559
rect -81824 -80603 -81768 -80559
rect -81724 -80603 -81668 -80559
rect -81624 -80603 -81568 -80559
rect -81524 -80603 -81468 -80559
rect -81424 -80603 -80968 -80559
rect -80924 -80603 -80868 -80559
rect -80824 -80603 -80768 -80559
rect -80724 -80603 -80668 -80559
rect -80624 -80603 -80568 -80559
rect -80524 -80603 -80468 -80559
rect -80424 -80603 -80368 -80559
rect -80324 -80603 -80268 -80559
rect -80224 -80603 -80168 -80559
rect -80124 -80603 -80068 -80559
rect -80024 -80603 -79968 -80559
rect -79924 -80603 -79868 -80559
rect -79824 -80603 -79768 -80559
rect -79724 -80603 -79668 -80559
rect -79624 -80603 -79568 -80559
rect -79524 -80603 -79468 -80559
rect -79424 -80603 -78968 -80559
rect -78924 -80603 -78868 -80559
rect -78824 -80603 -78768 -80559
rect -78724 -80603 -78668 -80559
rect -78624 -80603 -78568 -80559
rect -78524 -80603 -78468 -80559
rect -78424 -80603 -78368 -80559
rect -78324 -80603 -78268 -80559
rect -78224 -80603 -78168 -80559
rect -78124 -80603 -78068 -80559
rect -78024 -80603 -77968 -80559
rect -77924 -80603 -77868 -80559
rect -77824 -80603 -77768 -80559
rect -77724 -80603 -77668 -80559
rect -77624 -80603 -77568 -80559
rect -77524 -80603 -77468 -80559
rect -77424 -80603 -76968 -80559
rect -76924 -80603 -76868 -80559
rect -76824 -80603 -76768 -80559
rect -76724 -80603 -76668 -80559
rect -76624 -80603 -76568 -80559
rect -76524 -80603 -76468 -80559
rect -76424 -80603 -76368 -80559
rect -76324 -80603 -76268 -80559
rect -76224 -80603 -76168 -80559
rect -76124 -80603 -76068 -80559
rect -76024 -80603 -75968 -80559
rect -75924 -80603 -75868 -80559
rect -75824 -80603 -75768 -80559
rect -75724 -80603 -75668 -80559
rect -75624 -80603 -75568 -80559
rect -75524 -80603 -75468 -80559
rect -75424 -80603 -71799 -80559
rect -87194 -80659 -71799 -80603
rect -87194 -80703 -82968 -80659
rect -82924 -80703 -82868 -80659
rect -82824 -80703 -82768 -80659
rect -82724 -80703 -82668 -80659
rect -82624 -80703 -82568 -80659
rect -82524 -80703 -82468 -80659
rect -82424 -80703 -82368 -80659
rect -82324 -80703 -82268 -80659
rect -82224 -80703 -82168 -80659
rect -82124 -80703 -82068 -80659
rect -82024 -80703 -81968 -80659
rect -81924 -80703 -81868 -80659
rect -81824 -80703 -81768 -80659
rect -81724 -80703 -81668 -80659
rect -81624 -80703 -81568 -80659
rect -81524 -80703 -81468 -80659
rect -81424 -80703 -80968 -80659
rect -80924 -80703 -80868 -80659
rect -80824 -80703 -80768 -80659
rect -80724 -80703 -80668 -80659
rect -80624 -80703 -80568 -80659
rect -80524 -80703 -80468 -80659
rect -80424 -80703 -80368 -80659
rect -80324 -80703 -80268 -80659
rect -80224 -80703 -80168 -80659
rect -80124 -80703 -80068 -80659
rect -80024 -80703 -79968 -80659
rect -79924 -80703 -79868 -80659
rect -79824 -80703 -79768 -80659
rect -79724 -80703 -79668 -80659
rect -79624 -80703 -79568 -80659
rect -79524 -80703 -79468 -80659
rect -79424 -80703 -78968 -80659
rect -78924 -80703 -78868 -80659
rect -78824 -80703 -78768 -80659
rect -78724 -80703 -78668 -80659
rect -78624 -80703 -78568 -80659
rect -78524 -80703 -78468 -80659
rect -78424 -80703 -78368 -80659
rect -78324 -80703 -78268 -80659
rect -78224 -80703 -78168 -80659
rect -78124 -80703 -78068 -80659
rect -78024 -80703 -77968 -80659
rect -77924 -80703 -77868 -80659
rect -77824 -80703 -77768 -80659
rect -77724 -80703 -77668 -80659
rect -77624 -80703 -77568 -80659
rect -77524 -80703 -77468 -80659
rect -77424 -80703 -76968 -80659
rect -76924 -80703 -76868 -80659
rect -76824 -80703 -76768 -80659
rect -76724 -80703 -76668 -80659
rect -76624 -80703 -76568 -80659
rect -76524 -80703 -76468 -80659
rect -76424 -80703 -76368 -80659
rect -76324 -80703 -76268 -80659
rect -76224 -80703 -76168 -80659
rect -76124 -80703 -76068 -80659
rect -76024 -80703 -75968 -80659
rect -75924 -80703 -75868 -80659
rect -75824 -80703 -75768 -80659
rect -75724 -80703 -75668 -80659
rect -75624 -80703 -75568 -80659
rect -75524 -80703 -75468 -80659
rect -75424 -80703 -71799 -80659
rect -87194 -80759 -71799 -80703
rect -87194 -80803 -82968 -80759
rect -82924 -80803 -82868 -80759
rect -82824 -80803 -82768 -80759
rect -82724 -80803 -82668 -80759
rect -82624 -80803 -82568 -80759
rect -82524 -80803 -82468 -80759
rect -82424 -80803 -82368 -80759
rect -82324 -80803 -82268 -80759
rect -82224 -80803 -82168 -80759
rect -82124 -80803 -82068 -80759
rect -82024 -80803 -81968 -80759
rect -81924 -80803 -81868 -80759
rect -81824 -80803 -81768 -80759
rect -81724 -80803 -81668 -80759
rect -81624 -80803 -81568 -80759
rect -81524 -80803 -81468 -80759
rect -81424 -80803 -80968 -80759
rect -80924 -80803 -80868 -80759
rect -80824 -80803 -80768 -80759
rect -80724 -80803 -80668 -80759
rect -80624 -80803 -80568 -80759
rect -80524 -80803 -80468 -80759
rect -80424 -80803 -80368 -80759
rect -80324 -80803 -80268 -80759
rect -80224 -80803 -80168 -80759
rect -80124 -80803 -80068 -80759
rect -80024 -80803 -79968 -80759
rect -79924 -80803 -79868 -80759
rect -79824 -80803 -79768 -80759
rect -79724 -80803 -79668 -80759
rect -79624 -80803 -79568 -80759
rect -79524 -80803 -79468 -80759
rect -79424 -80803 -78968 -80759
rect -78924 -80803 -78868 -80759
rect -78824 -80803 -78768 -80759
rect -78724 -80803 -78668 -80759
rect -78624 -80803 -78568 -80759
rect -78524 -80803 -78468 -80759
rect -78424 -80803 -78368 -80759
rect -78324 -80803 -78268 -80759
rect -78224 -80803 -78168 -80759
rect -78124 -80803 -78068 -80759
rect -78024 -80803 -77968 -80759
rect -77924 -80803 -77868 -80759
rect -77824 -80803 -77768 -80759
rect -77724 -80803 -77668 -80759
rect -77624 -80803 -77568 -80759
rect -77524 -80803 -77468 -80759
rect -77424 -80803 -76968 -80759
rect -76924 -80803 -76868 -80759
rect -76824 -80803 -76768 -80759
rect -76724 -80803 -76668 -80759
rect -76624 -80803 -76568 -80759
rect -76524 -80803 -76468 -80759
rect -76424 -80803 -76368 -80759
rect -76324 -80803 -76268 -80759
rect -76224 -80803 -76168 -80759
rect -76124 -80803 -76068 -80759
rect -76024 -80803 -75968 -80759
rect -75924 -80803 -75868 -80759
rect -75824 -80803 -75768 -80759
rect -75724 -80803 -75668 -80759
rect -75624 -80803 -75568 -80759
rect -75524 -80803 -75468 -80759
rect -75424 -80803 -71799 -80759
rect -87194 -80859 -71799 -80803
rect -87194 -80903 -82968 -80859
rect -82924 -80903 -82868 -80859
rect -82824 -80903 -82768 -80859
rect -82724 -80903 -82668 -80859
rect -82624 -80903 -82568 -80859
rect -82524 -80903 -82468 -80859
rect -82424 -80903 -82368 -80859
rect -82324 -80903 -82268 -80859
rect -82224 -80903 -82168 -80859
rect -82124 -80903 -82068 -80859
rect -82024 -80903 -81968 -80859
rect -81924 -80903 -81868 -80859
rect -81824 -80903 -81768 -80859
rect -81724 -80903 -81668 -80859
rect -81624 -80903 -81568 -80859
rect -81524 -80903 -81468 -80859
rect -81424 -80903 -80968 -80859
rect -80924 -80903 -80868 -80859
rect -80824 -80903 -80768 -80859
rect -80724 -80903 -80668 -80859
rect -80624 -80903 -80568 -80859
rect -80524 -80903 -80468 -80859
rect -80424 -80903 -80368 -80859
rect -80324 -80903 -80268 -80859
rect -80224 -80903 -80168 -80859
rect -80124 -80903 -80068 -80859
rect -80024 -80903 -79968 -80859
rect -79924 -80903 -79868 -80859
rect -79824 -80903 -79768 -80859
rect -79724 -80903 -79668 -80859
rect -79624 -80903 -79568 -80859
rect -79524 -80903 -79468 -80859
rect -79424 -80903 -78968 -80859
rect -78924 -80903 -78868 -80859
rect -78824 -80903 -78768 -80859
rect -78724 -80903 -78668 -80859
rect -78624 -80903 -78568 -80859
rect -78524 -80903 -78468 -80859
rect -78424 -80903 -78368 -80859
rect -78324 -80903 -78268 -80859
rect -78224 -80903 -78168 -80859
rect -78124 -80903 -78068 -80859
rect -78024 -80903 -77968 -80859
rect -77924 -80903 -77868 -80859
rect -77824 -80903 -77768 -80859
rect -77724 -80903 -77668 -80859
rect -77624 -80903 -77568 -80859
rect -77524 -80903 -77468 -80859
rect -77424 -80903 -76968 -80859
rect -76924 -80903 -76868 -80859
rect -76824 -80903 -76768 -80859
rect -76724 -80903 -76668 -80859
rect -76624 -80903 -76568 -80859
rect -76524 -80903 -76468 -80859
rect -76424 -80903 -76368 -80859
rect -76324 -80903 -76268 -80859
rect -76224 -80903 -76168 -80859
rect -76124 -80903 -76068 -80859
rect -76024 -80903 -75968 -80859
rect -75924 -80903 -75868 -80859
rect -75824 -80903 -75768 -80859
rect -75724 -80903 -75668 -80859
rect -75624 -80903 -75568 -80859
rect -75524 -80903 -75468 -80859
rect -75424 -80903 -71799 -80859
rect -87194 -80959 -71799 -80903
rect -87194 -81003 -82968 -80959
rect -82924 -81003 -82868 -80959
rect -82824 -81003 -82768 -80959
rect -82724 -81003 -82668 -80959
rect -82624 -81003 -82568 -80959
rect -82524 -81003 -82468 -80959
rect -82424 -81003 -82368 -80959
rect -82324 -81003 -82268 -80959
rect -82224 -81003 -82168 -80959
rect -82124 -81003 -82068 -80959
rect -82024 -81003 -81968 -80959
rect -81924 -81003 -81868 -80959
rect -81824 -81003 -81768 -80959
rect -81724 -81003 -81668 -80959
rect -81624 -81003 -81568 -80959
rect -81524 -81003 -81468 -80959
rect -81424 -81003 -80968 -80959
rect -80924 -81003 -80868 -80959
rect -80824 -81003 -80768 -80959
rect -80724 -81003 -80668 -80959
rect -80624 -81003 -80568 -80959
rect -80524 -81003 -80468 -80959
rect -80424 -81003 -80368 -80959
rect -80324 -81003 -80268 -80959
rect -80224 -81003 -80168 -80959
rect -80124 -81003 -80068 -80959
rect -80024 -81003 -79968 -80959
rect -79924 -81003 -79868 -80959
rect -79824 -81003 -79768 -80959
rect -79724 -81003 -79668 -80959
rect -79624 -81003 -79568 -80959
rect -79524 -81003 -79468 -80959
rect -79424 -81003 -78968 -80959
rect -78924 -81003 -78868 -80959
rect -78824 -81003 -78768 -80959
rect -78724 -81003 -78668 -80959
rect -78624 -81003 -78568 -80959
rect -78524 -81003 -78468 -80959
rect -78424 -81003 -78368 -80959
rect -78324 -81003 -78268 -80959
rect -78224 -81003 -78168 -80959
rect -78124 -81003 -78068 -80959
rect -78024 -81003 -77968 -80959
rect -77924 -81003 -77868 -80959
rect -77824 -81003 -77768 -80959
rect -77724 -81003 -77668 -80959
rect -77624 -81003 -77568 -80959
rect -77524 -81003 -77468 -80959
rect -77424 -81003 -76968 -80959
rect -76924 -81003 -76868 -80959
rect -76824 -81003 -76768 -80959
rect -76724 -81003 -76668 -80959
rect -76624 -81003 -76568 -80959
rect -76524 -81003 -76468 -80959
rect -76424 -81003 -76368 -80959
rect -76324 -81003 -76268 -80959
rect -76224 -81003 -76168 -80959
rect -76124 -81003 -76068 -80959
rect -76024 -81003 -75968 -80959
rect -75924 -81003 -75868 -80959
rect -75824 -81003 -75768 -80959
rect -75724 -81003 -75668 -80959
rect -75624 -81003 -75568 -80959
rect -75524 -81003 -75468 -80959
rect -75424 -81003 -71799 -80959
rect -87194 -81059 -71799 -81003
rect -87194 -81103 -82968 -81059
rect -82924 -81103 -82868 -81059
rect -82824 -81103 -82768 -81059
rect -82724 -81103 -82668 -81059
rect -82624 -81103 -82568 -81059
rect -82524 -81103 -82468 -81059
rect -82424 -81103 -82368 -81059
rect -82324 -81103 -82268 -81059
rect -82224 -81103 -82168 -81059
rect -82124 -81103 -82068 -81059
rect -82024 -81103 -81968 -81059
rect -81924 -81103 -81868 -81059
rect -81824 -81103 -81768 -81059
rect -81724 -81103 -81668 -81059
rect -81624 -81103 -81568 -81059
rect -81524 -81103 -81468 -81059
rect -81424 -81103 -80968 -81059
rect -80924 -81103 -80868 -81059
rect -80824 -81103 -80768 -81059
rect -80724 -81103 -80668 -81059
rect -80624 -81103 -80568 -81059
rect -80524 -81103 -80468 -81059
rect -80424 -81103 -80368 -81059
rect -80324 -81103 -80268 -81059
rect -80224 -81103 -80168 -81059
rect -80124 -81103 -80068 -81059
rect -80024 -81103 -79968 -81059
rect -79924 -81103 -79868 -81059
rect -79824 -81103 -79768 -81059
rect -79724 -81103 -79668 -81059
rect -79624 -81103 -79568 -81059
rect -79524 -81103 -79468 -81059
rect -79424 -81103 -78968 -81059
rect -78924 -81103 -78868 -81059
rect -78824 -81103 -78768 -81059
rect -78724 -81103 -78668 -81059
rect -78624 -81103 -78568 -81059
rect -78524 -81103 -78468 -81059
rect -78424 -81103 -78368 -81059
rect -78324 -81103 -78268 -81059
rect -78224 -81103 -78168 -81059
rect -78124 -81103 -78068 -81059
rect -78024 -81103 -77968 -81059
rect -77924 -81103 -77868 -81059
rect -77824 -81103 -77768 -81059
rect -77724 -81103 -77668 -81059
rect -77624 -81103 -77568 -81059
rect -77524 -81103 -77468 -81059
rect -77424 -81103 -76968 -81059
rect -76924 -81103 -76868 -81059
rect -76824 -81103 -76768 -81059
rect -76724 -81103 -76668 -81059
rect -76624 -81103 -76568 -81059
rect -76524 -81103 -76468 -81059
rect -76424 -81103 -76368 -81059
rect -76324 -81103 -76268 -81059
rect -76224 -81103 -76168 -81059
rect -76124 -81103 -76068 -81059
rect -76024 -81103 -75968 -81059
rect -75924 -81103 -75868 -81059
rect -75824 -81103 -75768 -81059
rect -75724 -81103 -75668 -81059
rect -75624 -81103 -75568 -81059
rect -75524 -81103 -75468 -81059
rect -75424 -81103 -71799 -81059
rect -87194 -81159 -71799 -81103
rect -87194 -81203 -82968 -81159
rect -82924 -81203 -82868 -81159
rect -82824 -81203 -82768 -81159
rect -82724 -81203 -82668 -81159
rect -82624 -81203 -82568 -81159
rect -82524 -81203 -82468 -81159
rect -82424 -81203 -82368 -81159
rect -82324 -81203 -82268 -81159
rect -82224 -81203 -82168 -81159
rect -82124 -81203 -82068 -81159
rect -82024 -81203 -81968 -81159
rect -81924 -81203 -81868 -81159
rect -81824 -81203 -81768 -81159
rect -81724 -81203 -81668 -81159
rect -81624 -81203 -81568 -81159
rect -81524 -81203 -81468 -81159
rect -81424 -81203 -80968 -81159
rect -80924 -81203 -80868 -81159
rect -80824 -81203 -80768 -81159
rect -80724 -81203 -80668 -81159
rect -80624 -81203 -80568 -81159
rect -80524 -81203 -80468 -81159
rect -80424 -81203 -80368 -81159
rect -80324 -81203 -80268 -81159
rect -80224 -81203 -80168 -81159
rect -80124 -81203 -80068 -81159
rect -80024 -81203 -79968 -81159
rect -79924 -81203 -79868 -81159
rect -79824 -81203 -79768 -81159
rect -79724 -81203 -79668 -81159
rect -79624 -81203 -79568 -81159
rect -79524 -81203 -79468 -81159
rect -79424 -81203 -78968 -81159
rect -78924 -81203 -78868 -81159
rect -78824 -81203 -78768 -81159
rect -78724 -81203 -78668 -81159
rect -78624 -81203 -78568 -81159
rect -78524 -81203 -78468 -81159
rect -78424 -81203 -78368 -81159
rect -78324 -81203 -78268 -81159
rect -78224 -81203 -78168 -81159
rect -78124 -81203 -78068 -81159
rect -78024 -81203 -77968 -81159
rect -77924 -81203 -77868 -81159
rect -77824 -81203 -77768 -81159
rect -77724 -81203 -77668 -81159
rect -77624 -81203 -77568 -81159
rect -77524 -81203 -77468 -81159
rect -77424 -81203 -76968 -81159
rect -76924 -81203 -76868 -81159
rect -76824 -81203 -76768 -81159
rect -76724 -81203 -76668 -81159
rect -76624 -81203 -76568 -81159
rect -76524 -81203 -76468 -81159
rect -76424 -81203 -76368 -81159
rect -76324 -81203 -76268 -81159
rect -76224 -81203 -76168 -81159
rect -76124 -81203 -76068 -81159
rect -76024 -81203 -75968 -81159
rect -75924 -81203 -75868 -81159
rect -75824 -81203 -75768 -81159
rect -75724 -81203 -75668 -81159
rect -75624 -81203 -75568 -81159
rect -75524 -81203 -75468 -81159
rect -75424 -81203 -71799 -81159
rect -87194 -81259 -71799 -81203
rect -87194 -81303 -82968 -81259
rect -82924 -81303 -82868 -81259
rect -82824 -81303 -82768 -81259
rect -82724 -81303 -82668 -81259
rect -82624 -81303 -82568 -81259
rect -82524 -81303 -82468 -81259
rect -82424 -81303 -82368 -81259
rect -82324 -81303 -82268 -81259
rect -82224 -81303 -82168 -81259
rect -82124 -81303 -82068 -81259
rect -82024 -81303 -81968 -81259
rect -81924 -81303 -81868 -81259
rect -81824 -81303 -81768 -81259
rect -81724 -81303 -81668 -81259
rect -81624 -81303 -81568 -81259
rect -81524 -81303 -81468 -81259
rect -81424 -81303 -80968 -81259
rect -80924 -81303 -80868 -81259
rect -80824 -81303 -80768 -81259
rect -80724 -81303 -80668 -81259
rect -80624 -81303 -80568 -81259
rect -80524 -81303 -80468 -81259
rect -80424 -81303 -80368 -81259
rect -80324 -81303 -80268 -81259
rect -80224 -81303 -80168 -81259
rect -80124 -81303 -80068 -81259
rect -80024 -81303 -79968 -81259
rect -79924 -81303 -79868 -81259
rect -79824 -81303 -79768 -81259
rect -79724 -81303 -79668 -81259
rect -79624 -81303 -79568 -81259
rect -79524 -81303 -79468 -81259
rect -79424 -81303 -78968 -81259
rect -78924 -81303 -78868 -81259
rect -78824 -81303 -78768 -81259
rect -78724 -81303 -78668 -81259
rect -78624 -81303 -78568 -81259
rect -78524 -81303 -78468 -81259
rect -78424 -81303 -78368 -81259
rect -78324 -81303 -78268 -81259
rect -78224 -81303 -78168 -81259
rect -78124 -81303 -78068 -81259
rect -78024 -81303 -77968 -81259
rect -77924 -81303 -77868 -81259
rect -77824 -81303 -77768 -81259
rect -77724 -81303 -77668 -81259
rect -77624 -81303 -77568 -81259
rect -77524 -81303 -77468 -81259
rect -77424 -81303 -76968 -81259
rect -76924 -81303 -76868 -81259
rect -76824 -81303 -76768 -81259
rect -76724 -81303 -76668 -81259
rect -76624 -81303 -76568 -81259
rect -76524 -81303 -76468 -81259
rect -76424 -81303 -76368 -81259
rect -76324 -81303 -76268 -81259
rect -76224 -81303 -76168 -81259
rect -76124 -81303 -76068 -81259
rect -76024 -81303 -75968 -81259
rect -75924 -81303 -75868 -81259
rect -75824 -81303 -75768 -81259
rect -75724 -81303 -75668 -81259
rect -75624 -81303 -75568 -81259
rect -75524 -81303 -75468 -81259
rect -75424 -81303 -71799 -81259
rect -87194 -81359 -71799 -81303
rect -87194 -81403 -82968 -81359
rect -82924 -81403 -82868 -81359
rect -82824 -81403 -82768 -81359
rect -82724 -81403 -82668 -81359
rect -82624 -81403 -82568 -81359
rect -82524 -81403 -82468 -81359
rect -82424 -81403 -82368 -81359
rect -82324 -81403 -82268 -81359
rect -82224 -81403 -82168 -81359
rect -82124 -81403 -82068 -81359
rect -82024 -81403 -81968 -81359
rect -81924 -81403 -81868 -81359
rect -81824 -81403 -81768 -81359
rect -81724 -81403 -81668 -81359
rect -81624 -81403 -81568 -81359
rect -81524 -81403 -81468 -81359
rect -81424 -81403 -80968 -81359
rect -80924 -81403 -80868 -81359
rect -80824 -81403 -80768 -81359
rect -80724 -81403 -80668 -81359
rect -80624 -81403 -80568 -81359
rect -80524 -81403 -80468 -81359
rect -80424 -81403 -80368 -81359
rect -80324 -81403 -80268 -81359
rect -80224 -81403 -80168 -81359
rect -80124 -81403 -80068 -81359
rect -80024 -81403 -79968 -81359
rect -79924 -81403 -79868 -81359
rect -79824 -81403 -79768 -81359
rect -79724 -81403 -79668 -81359
rect -79624 -81403 -79568 -81359
rect -79524 -81403 -79468 -81359
rect -79424 -81403 -78968 -81359
rect -78924 -81403 -78868 -81359
rect -78824 -81403 -78768 -81359
rect -78724 -81403 -78668 -81359
rect -78624 -81403 -78568 -81359
rect -78524 -81403 -78468 -81359
rect -78424 -81403 -78368 -81359
rect -78324 -81403 -78268 -81359
rect -78224 -81403 -78168 -81359
rect -78124 -81403 -78068 -81359
rect -78024 -81403 -77968 -81359
rect -77924 -81403 -77868 -81359
rect -77824 -81403 -77768 -81359
rect -77724 -81403 -77668 -81359
rect -77624 -81403 -77568 -81359
rect -77524 -81403 -77468 -81359
rect -77424 -81403 -76968 -81359
rect -76924 -81403 -76868 -81359
rect -76824 -81403 -76768 -81359
rect -76724 -81403 -76668 -81359
rect -76624 -81403 -76568 -81359
rect -76524 -81403 -76468 -81359
rect -76424 -81403 -76368 -81359
rect -76324 -81403 -76268 -81359
rect -76224 -81403 -76168 -81359
rect -76124 -81403 -76068 -81359
rect -76024 -81403 -75968 -81359
rect -75924 -81403 -75868 -81359
rect -75824 -81403 -75768 -81359
rect -75724 -81403 -75668 -81359
rect -75624 -81403 -75568 -81359
rect -75524 -81403 -75468 -81359
rect -75424 -81403 -71799 -81359
rect -87194 -81459 -71799 -81403
rect -87194 -81503 -82968 -81459
rect -82924 -81503 -82868 -81459
rect -82824 -81503 -82768 -81459
rect -82724 -81503 -82668 -81459
rect -82624 -81503 -82568 -81459
rect -82524 -81503 -82468 -81459
rect -82424 -81503 -82368 -81459
rect -82324 -81503 -82268 -81459
rect -82224 -81503 -82168 -81459
rect -82124 -81503 -82068 -81459
rect -82024 -81503 -81968 -81459
rect -81924 -81503 -81868 -81459
rect -81824 -81503 -81768 -81459
rect -81724 -81503 -81668 -81459
rect -81624 -81503 -81568 -81459
rect -81524 -81503 -81468 -81459
rect -81424 -81503 -80968 -81459
rect -80924 -81503 -80868 -81459
rect -80824 -81503 -80768 -81459
rect -80724 -81503 -80668 -81459
rect -80624 -81503 -80568 -81459
rect -80524 -81503 -80468 -81459
rect -80424 -81503 -80368 -81459
rect -80324 -81503 -80268 -81459
rect -80224 -81503 -80168 -81459
rect -80124 -81503 -80068 -81459
rect -80024 -81503 -79968 -81459
rect -79924 -81503 -79868 -81459
rect -79824 -81503 -79768 -81459
rect -79724 -81503 -79668 -81459
rect -79624 -81503 -79568 -81459
rect -79524 -81503 -79468 -81459
rect -79424 -81503 -78968 -81459
rect -78924 -81503 -78868 -81459
rect -78824 -81503 -78768 -81459
rect -78724 -81503 -78668 -81459
rect -78624 -81503 -78568 -81459
rect -78524 -81503 -78468 -81459
rect -78424 -81503 -78368 -81459
rect -78324 -81503 -78268 -81459
rect -78224 -81503 -78168 -81459
rect -78124 -81503 -78068 -81459
rect -78024 -81503 -77968 -81459
rect -77924 -81503 -77868 -81459
rect -77824 -81503 -77768 -81459
rect -77724 -81503 -77668 -81459
rect -77624 -81503 -77568 -81459
rect -77524 -81503 -77468 -81459
rect -77424 -81503 -76968 -81459
rect -76924 -81503 -76868 -81459
rect -76824 -81503 -76768 -81459
rect -76724 -81503 -76668 -81459
rect -76624 -81503 -76568 -81459
rect -76524 -81503 -76468 -81459
rect -76424 -81503 -76368 -81459
rect -76324 -81503 -76268 -81459
rect -76224 -81503 -76168 -81459
rect -76124 -81503 -76068 -81459
rect -76024 -81503 -75968 -81459
rect -75924 -81503 -75868 -81459
rect -75824 -81503 -75768 -81459
rect -75724 -81503 -75668 -81459
rect -75624 -81503 -75568 -81459
rect -75524 -81503 -75468 -81459
rect -75424 -81503 -71799 -81459
rect -87194 -81559 -71799 -81503
rect -87194 -81603 -82968 -81559
rect -82924 -81603 -82868 -81559
rect -82824 -81603 -82768 -81559
rect -82724 -81603 -82668 -81559
rect -82624 -81603 -82568 -81559
rect -82524 -81603 -82468 -81559
rect -82424 -81603 -82368 -81559
rect -82324 -81603 -82268 -81559
rect -82224 -81603 -82168 -81559
rect -82124 -81603 -82068 -81559
rect -82024 -81603 -81968 -81559
rect -81924 -81603 -81868 -81559
rect -81824 -81603 -81768 -81559
rect -81724 -81603 -81668 -81559
rect -81624 -81603 -81568 -81559
rect -81524 -81603 -81468 -81559
rect -81424 -81603 -80968 -81559
rect -80924 -81603 -80868 -81559
rect -80824 -81603 -80768 -81559
rect -80724 -81603 -80668 -81559
rect -80624 -81603 -80568 -81559
rect -80524 -81603 -80468 -81559
rect -80424 -81603 -80368 -81559
rect -80324 -81603 -80268 -81559
rect -80224 -81603 -80168 -81559
rect -80124 -81603 -80068 -81559
rect -80024 -81603 -79968 -81559
rect -79924 -81603 -79868 -81559
rect -79824 -81603 -79768 -81559
rect -79724 -81603 -79668 -81559
rect -79624 -81603 -79568 -81559
rect -79524 -81603 -79468 -81559
rect -79424 -81603 -78968 -81559
rect -78924 -81603 -78868 -81559
rect -78824 -81603 -78768 -81559
rect -78724 -81603 -78668 -81559
rect -78624 -81603 -78568 -81559
rect -78524 -81603 -78468 -81559
rect -78424 -81603 -78368 -81559
rect -78324 -81603 -78268 -81559
rect -78224 -81603 -78168 -81559
rect -78124 -81603 -78068 -81559
rect -78024 -81603 -77968 -81559
rect -77924 -81603 -77868 -81559
rect -77824 -81603 -77768 -81559
rect -77724 -81603 -77668 -81559
rect -77624 -81603 -77568 -81559
rect -77524 -81603 -77468 -81559
rect -77424 -81603 -76968 -81559
rect -76924 -81603 -76868 -81559
rect -76824 -81603 -76768 -81559
rect -76724 -81603 -76668 -81559
rect -76624 -81603 -76568 -81559
rect -76524 -81603 -76468 -81559
rect -76424 -81603 -76368 -81559
rect -76324 -81603 -76268 -81559
rect -76224 -81603 -76168 -81559
rect -76124 -81603 -76068 -81559
rect -76024 -81603 -75968 -81559
rect -75924 -81603 -75868 -81559
rect -75824 -81603 -75768 -81559
rect -75724 -81603 -75668 -81559
rect -75624 -81603 -75568 -81559
rect -75524 -81603 -75468 -81559
rect -75424 -81603 -71799 -81559
rect -87194 -81659 -71799 -81603
rect -87194 -81703 -82968 -81659
rect -82924 -81703 -82868 -81659
rect -82824 -81703 -82768 -81659
rect -82724 -81703 -82668 -81659
rect -82624 -81703 -82568 -81659
rect -82524 -81703 -82468 -81659
rect -82424 -81703 -82368 -81659
rect -82324 -81703 -82268 -81659
rect -82224 -81703 -82168 -81659
rect -82124 -81703 -82068 -81659
rect -82024 -81703 -81968 -81659
rect -81924 -81703 -81868 -81659
rect -81824 -81703 -81768 -81659
rect -81724 -81703 -81668 -81659
rect -81624 -81703 -81568 -81659
rect -81524 -81703 -81468 -81659
rect -81424 -81703 -80968 -81659
rect -80924 -81703 -80868 -81659
rect -80824 -81703 -80768 -81659
rect -80724 -81703 -80668 -81659
rect -80624 -81703 -80568 -81659
rect -80524 -81703 -80468 -81659
rect -80424 -81703 -80368 -81659
rect -80324 -81703 -80268 -81659
rect -80224 -81703 -80168 -81659
rect -80124 -81703 -80068 -81659
rect -80024 -81703 -79968 -81659
rect -79924 -81703 -79868 -81659
rect -79824 -81703 -79768 -81659
rect -79724 -81703 -79668 -81659
rect -79624 -81703 -79568 -81659
rect -79524 -81703 -79468 -81659
rect -79424 -81703 -78968 -81659
rect -78924 -81703 -78868 -81659
rect -78824 -81703 -78768 -81659
rect -78724 -81703 -78668 -81659
rect -78624 -81703 -78568 -81659
rect -78524 -81703 -78468 -81659
rect -78424 -81703 -78368 -81659
rect -78324 -81703 -78268 -81659
rect -78224 -81703 -78168 -81659
rect -78124 -81703 -78068 -81659
rect -78024 -81703 -77968 -81659
rect -77924 -81703 -77868 -81659
rect -77824 -81703 -77768 -81659
rect -77724 -81703 -77668 -81659
rect -77624 -81703 -77568 -81659
rect -77524 -81703 -77468 -81659
rect -77424 -81703 -76968 -81659
rect -76924 -81703 -76868 -81659
rect -76824 -81703 -76768 -81659
rect -76724 -81703 -76668 -81659
rect -76624 -81703 -76568 -81659
rect -76524 -81703 -76468 -81659
rect -76424 -81703 -76368 -81659
rect -76324 -81703 -76268 -81659
rect -76224 -81703 -76168 -81659
rect -76124 -81703 -76068 -81659
rect -76024 -81703 -75968 -81659
rect -75924 -81703 -75868 -81659
rect -75824 -81703 -75768 -81659
rect -75724 -81703 -75668 -81659
rect -75624 -81703 -75568 -81659
rect -75524 -81703 -75468 -81659
rect -75424 -81703 -71799 -81659
rect -87194 -81759 -71799 -81703
rect -87194 -81803 -82968 -81759
rect -82924 -81803 -82868 -81759
rect -82824 -81803 -82768 -81759
rect -82724 -81803 -82668 -81759
rect -82624 -81803 -82568 -81759
rect -82524 -81803 -82468 -81759
rect -82424 -81803 -82368 -81759
rect -82324 -81803 -82268 -81759
rect -82224 -81803 -82168 -81759
rect -82124 -81803 -82068 -81759
rect -82024 -81803 -81968 -81759
rect -81924 -81803 -81868 -81759
rect -81824 -81803 -81768 -81759
rect -81724 -81803 -81668 -81759
rect -81624 -81803 -81568 -81759
rect -81524 -81803 -81468 -81759
rect -81424 -81803 -80968 -81759
rect -80924 -81803 -80868 -81759
rect -80824 -81803 -80768 -81759
rect -80724 -81803 -80668 -81759
rect -80624 -81803 -80568 -81759
rect -80524 -81803 -80468 -81759
rect -80424 -81803 -80368 -81759
rect -80324 -81803 -80268 -81759
rect -80224 -81803 -80168 -81759
rect -80124 -81803 -80068 -81759
rect -80024 -81803 -79968 -81759
rect -79924 -81803 -79868 -81759
rect -79824 -81803 -79768 -81759
rect -79724 -81803 -79668 -81759
rect -79624 -81803 -79568 -81759
rect -79524 -81803 -79468 -81759
rect -79424 -81803 -78968 -81759
rect -78924 -81803 -78868 -81759
rect -78824 -81803 -78768 -81759
rect -78724 -81803 -78668 -81759
rect -78624 -81803 -78568 -81759
rect -78524 -81803 -78468 -81759
rect -78424 -81803 -78368 -81759
rect -78324 -81803 -78268 -81759
rect -78224 -81803 -78168 -81759
rect -78124 -81803 -78068 -81759
rect -78024 -81803 -77968 -81759
rect -77924 -81803 -77868 -81759
rect -77824 -81803 -77768 -81759
rect -77724 -81803 -77668 -81759
rect -77624 -81803 -77568 -81759
rect -77524 -81803 -77468 -81759
rect -77424 -81803 -76968 -81759
rect -76924 -81803 -76868 -81759
rect -76824 -81803 -76768 -81759
rect -76724 -81803 -76668 -81759
rect -76624 -81803 -76568 -81759
rect -76524 -81803 -76468 -81759
rect -76424 -81803 -76368 -81759
rect -76324 -81803 -76268 -81759
rect -76224 -81803 -76168 -81759
rect -76124 -81803 -76068 -81759
rect -76024 -81803 -75968 -81759
rect -75924 -81803 -75868 -81759
rect -75824 -81803 -75768 -81759
rect -75724 -81803 -75668 -81759
rect -75624 -81803 -75568 -81759
rect -75524 -81803 -75468 -81759
rect -75424 -81803 -71799 -81759
rect -87194 -81859 -71799 -81803
rect -87194 -81903 -82968 -81859
rect -82924 -81903 -82868 -81859
rect -82824 -81903 -82768 -81859
rect -82724 -81903 -82668 -81859
rect -82624 -81903 -82568 -81859
rect -82524 -81903 -82468 -81859
rect -82424 -81903 -82368 -81859
rect -82324 -81903 -82268 -81859
rect -82224 -81903 -82168 -81859
rect -82124 -81903 -82068 -81859
rect -82024 -81903 -81968 -81859
rect -81924 -81903 -81868 -81859
rect -81824 -81903 -81768 -81859
rect -81724 -81903 -81668 -81859
rect -81624 -81903 -81568 -81859
rect -81524 -81903 -81468 -81859
rect -81424 -81903 -80968 -81859
rect -80924 -81903 -80868 -81859
rect -80824 -81903 -80768 -81859
rect -80724 -81903 -80668 -81859
rect -80624 -81903 -80568 -81859
rect -80524 -81903 -80468 -81859
rect -80424 -81903 -80368 -81859
rect -80324 -81903 -80268 -81859
rect -80224 -81903 -80168 -81859
rect -80124 -81903 -80068 -81859
rect -80024 -81903 -79968 -81859
rect -79924 -81903 -79868 -81859
rect -79824 -81903 -79768 -81859
rect -79724 -81903 -79668 -81859
rect -79624 -81903 -79568 -81859
rect -79524 -81903 -79468 -81859
rect -79424 -81903 -78968 -81859
rect -78924 -81903 -78868 -81859
rect -78824 -81903 -78768 -81859
rect -78724 -81903 -78668 -81859
rect -78624 -81903 -78568 -81859
rect -78524 -81903 -78468 -81859
rect -78424 -81903 -78368 -81859
rect -78324 -81903 -78268 -81859
rect -78224 -81903 -78168 -81859
rect -78124 -81903 -78068 -81859
rect -78024 -81903 -77968 -81859
rect -77924 -81903 -77868 -81859
rect -77824 -81903 -77768 -81859
rect -77724 -81903 -77668 -81859
rect -77624 -81903 -77568 -81859
rect -77524 -81903 -77468 -81859
rect -77424 -81903 -76968 -81859
rect -76924 -81903 -76868 -81859
rect -76824 -81903 -76768 -81859
rect -76724 -81903 -76668 -81859
rect -76624 -81903 -76568 -81859
rect -76524 -81903 -76468 -81859
rect -76424 -81903 -76368 -81859
rect -76324 -81903 -76268 -81859
rect -76224 -81903 -76168 -81859
rect -76124 -81903 -76068 -81859
rect -76024 -81903 -75968 -81859
rect -75924 -81903 -75868 -81859
rect -75824 -81903 -75768 -81859
rect -75724 -81903 -75668 -81859
rect -75624 -81903 -75568 -81859
rect -75524 -81903 -75468 -81859
rect -75424 -81903 -71799 -81859
rect -87194 -81959 -71799 -81903
rect -87194 -82003 -82968 -81959
rect -82924 -82003 -82868 -81959
rect -82824 -82003 -82768 -81959
rect -82724 -82003 -82668 -81959
rect -82624 -82003 -82568 -81959
rect -82524 -82003 -82468 -81959
rect -82424 -82003 -82368 -81959
rect -82324 -82003 -82268 -81959
rect -82224 -82003 -82168 -81959
rect -82124 -82003 -82068 -81959
rect -82024 -82003 -81968 -81959
rect -81924 -82003 -81868 -81959
rect -81824 -82003 -81768 -81959
rect -81724 -82003 -81668 -81959
rect -81624 -82003 -81568 -81959
rect -81524 -82003 -81468 -81959
rect -81424 -82003 -80968 -81959
rect -80924 -82003 -80868 -81959
rect -80824 -82003 -80768 -81959
rect -80724 -82003 -80668 -81959
rect -80624 -82003 -80568 -81959
rect -80524 -82003 -80468 -81959
rect -80424 -82003 -80368 -81959
rect -80324 -82003 -80268 -81959
rect -80224 -82003 -80168 -81959
rect -80124 -82003 -80068 -81959
rect -80024 -82003 -79968 -81959
rect -79924 -82003 -79868 -81959
rect -79824 -82003 -79768 -81959
rect -79724 -82003 -79668 -81959
rect -79624 -82003 -79568 -81959
rect -79524 -82003 -79468 -81959
rect -79424 -82003 -78968 -81959
rect -78924 -82003 -78868 -81959
rect -78824 -82003 -78768 -81959
rect -78724 -82003 -78668 -81959
rect -78624 -82003 -78568 -81959
rect -78524 -82003 -78468 -81959
rect -78424 -82003 -78368 -81959
rect -78324 -82003 -78268 -81959
rect -78224 -82003 -78168 -81959
rect -78124 -82003 -78068 -81959
rect -78024 -82003 -77968 -81959
rect -77924 -82003 -77868 -81959
rect -77824 -82003 -77768 -81959
rect -77724 -82003 -77668 -81959
rect -77624 -82003 -77568 -81959
rect -77524 -82003 -77468 -81959
rect -77424 -82003 -76968 -81959
rect -76924 -82003 -76868 -81959
rect -76824 -82003 -76768 -81959
rect -76724 -82003 -76668 -81959
rect -76624 -82003 -76568 -81959
rect -76524 -82003 -76468 -81959
rect -76424 -82003 -76368 -81959
rect -76324 -82003 -76268 -81959
rect -76224 -82003 -76168 -81959
rect -76124 -82003 -76068 -81959
rect -76024 -82003 -75968 -81959
rect -75924 -82003 -75868 -81959
rect -75824 -82003 -75768 -81959
rect -75724 -82003 -75668 -81959
rect -75624 -82003 -75568 -81959
rect -75524 -82003 -75468 -81959
rect -75424 -82003 -71799 -81959
rect -87194 -140231 -71799 -82003
rect -50768 -80461 -42000 -80270
rect -50768 -80505 -50017 -80461
rect -49973 -80505 -49917 -80461
rect -49873 -80505 -49817 -80461
rect -49773 -80505 -49717 -80461
rect -49673 -80505 -49617 -80461
rect -49573 -80505 -49517 -80461
rect -49473 -80505 -49417 -80461
rect -49373 -80505 -49317 -80461
rect -49273 -80505 -49217 -80461
rect -49173 -80505 -49117 -80461
rect -49073 -80505 -49017 -80461
rect -48973 -80505 -48917 -80461
rect -48873 -80505 -48817 -80461
rect -48773 -80505 -48717 -80461
rect -48673 -80505 -48617 -80461
rect -48573 -80505 -48517 -80461
rect -48473 -80505 -48017 -80461
rect -47973 -80505 -47917 -80461
rect -47873 -80505 -47817 -80461
rect -47773 -80505 -47717 -80461
rect -47673 -80505 -47617 -80461
rect -47573 -80505 -47517 -80461
rect -47473 -80505 -47417 -80461
rect -47373 -80505 -47317 -80461
rect -47273 -80505 -47217 -80461
rect -47173 -80505 -47117 -80461
rect -47073 -80505 -47017 -80461
rect -46973 -80505 -46917 -80461
rect -46873 -80505 -46817 -80461
rect -46773 -80505 -46717 -80461
rect -46673 -80505 -46617 -80461
rect -46573 -80505 -46517 -80461
rect -46473 -80505 -46017 -80461
rect -45973 -80505 -45917 -80461
rect -45873 -80505 -45817 -80461
rect -45773 -80505 -45717 -80461
rect -45673 -80505 -45617 -80461
rect -45573 -80505 -45517 -80461
rect -45473 -80505 -45417 -80461
rect -45373 -80505 -45317 -80461
rect -45273 -80505 -45217 -80461
rect -45173 -80505 -45117 -80461
rect -45073 -80505 -45017 -80461
rect -44973 -80505 -44917 -80461
rect -44873 -80505 -44817 -80461
rect -44773 -80505 -44717 -80461
rect -44673 -80505 -44617 -80461
rect -44573 -80505 -44517 -80461
rect -44473 -80505 -44017 -80461
rect -43973 -80505 -43917 -80461
rect -43873 -80505 -43817 -80461
rect -43773 -80505 -43717 -80461
rect -43673 -80505 -43617 -80461
rect -43573 -80505 -43517 -80461
rect -43473 -80505 -43417 -80461
rect -43373 -80505 -43317 -80461
rect -43273 -80505 -43217 -80461
rect -43173 -80505 -43117 -80461
rect -43073 -80505 -43017 -80461
rect -42973 -80505 -42917 -80461
rect -42873 -80505 -42817 -80461
rect -42773 -80505 -42717 -80461
rect -42673 -80505 -42617 -80461
rect -42573 -80505 -42517 -80461
rect -42473 -80505 -42000 -80461
rect -50768 -80561 -42000 -80505
rect -50768 -80605 -50017 -80561
rect -49973 -80605 -49917 -80561
rect -49873 -80605 -49817 -80561
rect -49773 -80605 -49717 -80561
rect -49673 -80605 -49617 -80561
rect -49573 -80605 -49517 -80561
rect -49473 -80605 -49417 -80561
rect -49373 -80605 -49317 -80561
rect -49273 -80605 -49217 -80561
rect -49173 -80605 -49117 -80561
rect -49073 -80605 -49017 -80561
rect -48973 -80605 -48917 -80561
rect -48873 -80605 -48817 -80561
rect -48773 -80605 -48717 -80561
rect -48673 -80605 -48617 -80561
rect -48573 -80605 -48517 -80561
rect -48473 -80605 -48017 -80561
rect -47973 -80605 -47917 -80561
rect -47873 -80605 -47817 -80561
rect -47773 -80605 -47717 -80561
rect -47673 -80605 -47617 -80561
rect -47573 -80605 -47517 -80561
rect -47473 -80605 -47417 -80561
rect -47373 -80605 -47317 -80561
rect -47273 -80605 -47217 -80561
rect -47173 -80605 -47117 -80561
rect -47073 -80605 -47017 -80561
rect -46973 -80605 -46917 -80561
rect -46873 -80605 -46817 -80561
rect -46773 -80605 -46717 -80561
rect -46673 -80605 -46617 -80561
rect -46573 -80605 -46517 -80561
rect -46473 -80605 -46017 -80561
rect -45973 -80605 -45917 -80561
rect -45873 -80605 -45817 -80561
rect -45773 -80605 -45717 -80561
rect -45673 -80605 -45617 -80561
rect -45573 -80605 -45517 -80561
rect -45473 -80605 -45417 -80561
rect -45373 -80605 -45317 -80561
rect -45273 -80605 -45217 -80561
rect -45173 -80605 -45117 -80561
rect -45073 -80605 -45017 -80561
rect -44973 -80605 -44917 -80561
rect -44873 -80605 -44817 -80561
rect -44773 -80605 -44717 -80561
rect -44673 -80605 -44617 -80561
rect -44573 -80605 -44517 -80561
rect -44473 -80605 -44017 -80561
rect -43973 -80605 -43917 -80561
rect -43873 -80605 -43817 -80561
rect -43773 -80605 -43717 -80561
rect -43673 -80605 -43617 -80561
rect -43573 -80605 -43517 -80561
rect -43473 -80605 -43417 -80561
rect -43373 -80605 -43317 -80561
rect -43273 -80605 -43217 -80561
rect -43173 -80605 -43117 -80561
rect -43073 -80605 -43017 -80561
rect -42973 -80605 -42917 -80561
rect -42873 -80605 -42817 -80561
rect -42773 -80605 -42717 -80561
rect -42673 -80605 -42617 -80561
rect -42573 -80605 -42517 -80561
rect -42473 -80605 -42000 -80561
rect -50768 -80661 -42000 -80605
rect -50768 -80705 -50017 -80661
rect -49973 -80705 -49917 -80661
rect -49873 -80705 -49817 -80661
rect -49773 -80705 -49717 -80661
rect -49673 -80705 -49617 -80661
rect -49573 -80705 -49517 -80661
rect -49473 -80705 -49417 -80661
rect -49373 -80705 -49317 -80661
rect -49273 -80705 -49217 -80661
rect -49173 -80705 -49117 -80661
rect -49073 -80705 -49017 -80661
rect -48973 -80705 -48917 -80661
rect -48873 -80705 -48817 -80661
rect -48773 -80705 -48717 -80661
rect -48673 -80705 -48617 -80661
rect -48573 -80705 -48517 -80661
rect -48473 -80705 -48017 -80661
rect -47973 -80705 -47917 -80661
rect -47873 -80705 -47817 -80661
rect -47773 -80705 -47717 -80661
rect -47673 -80705 -47617 -80661
rect -47573 -80705 -47517 -80661
rect -47473 -80705 -47417 -80661
rect -47373 -80705 -47317 -80661
rect -47273 -80705 -47217 -80661
rect -47173 -80705 -47117 -80661
rect -47073 -80705 -47017 -80661
rect -46973 -80705 -46917 -80661
rect -46873 -80705 -46817 -80661
rect -46773 -80705 -46717 -80661
rect -46673 -80705 -46617 -80661
rect -46573 -80705 -46517 -80661
rect -46473 -80705 -46017 -80661
rect -45973 -80705 -45917 -80661
rect -45873 -80705 -45817 -80661
rect -45773 -80705 -45717 -80661
rect -45673 -80705 -45617 -80661
rect -45573 -80705 -45517 -80661
rect -45473 -80705 -45417 -80661
rect -45373 -80705 -45317 -80661
rect -45273 -80705 -45217 -80661
rect -45173 -80705 -45117 -80661
rect -45073 -80705 -45017 -80661
rect -44973 -80705 -44917 -80661
rect -44873 -80705 -44817 -80661
rect -44773 -80705 -44717 -80661
rect -44673 -80705 -44617 -80661
rect -44573 -80705 -44517 -80661
rect -44473 -80705 -44017 -80661
rect -43973 -80705 -43917 -80661
rect -43873 -80705 -43817 -80661
rect -43773 -80705 -43717 -80661
rect -43673 -80705 -43617 -80661
rect -43573 -80705 -43517 -80661
rect -43473 -80705 -43417 -80661
rect -43373 -80705 -43317 -80661
rect -43273 -80705 -43217 -80661
rect -43173 -80705 -43117 -80661
rect -43073 -80705 -43017 -80661
rect -42973 -80705 -42917 -80661
rect -42873 -80705 -42817 -80661
rect -42773 -80705 -42717 -80661
rect -42673 -80705 -42617 -80661
rect -42573 -80705 -42517 -80661
rect -42473 -80705 -42000 -80661
rect -50768 -80761 -42000 -80705
rect -50768 -80805 -50017 -80761
rect -49973 -80805 -49917 -80761
rect -49873 -80805 -49817 -80761
rect -49773 -80805 -49717 -80761
rect -49673 -80805 -49617 -80761
rect -49573 -80805 -49517 -80761
rect -49473 -80805 -49417 -80761
rect -49373 -80805 -49317 -80761
rect -49273 -80805 -49217 -80761
rect -49173 -80805 -49117 -80761
rect -49073 -80805 -49017 -80761
rect -48973 -80805 -48917 -80761
rect -48873 -80805 -48817 -80761
rect -48773 -80805 -48717 -80761
rect -48673 -80805 -48617 -80761
rect -48573 -80805 -48517 -80761
rect -48473 -80805 -48017 -80761
rect -47973 -80805 -47917 -80761
rect -47873 -80805 -47817 -80761
rect -47773 -80805 -47717 -80761
rect -47673 -80805 -47617 -80761
rect -47573 -80805 -47517 -80761
rect -47473 -80805 -47417 -80761
rect -47373 -80805 -47317 -80761
rect -47273 -80805 -47217 -80761
rect -47173 -80805 -47117 -80761
rect -47073 -80805 -47017 -80761
rect -46973 -80805 -46917 -80761
rect -46873 -80805 -46817 -80761
rect -46773 -80805 -46717 -80761
rect -46673 -80805 -46617 -80761
rect -46573 -80805 -46517 -80761
rect -46473 -80805 -46017 -80761
rect -45973 -80805 -45917 -80761
rect -45873 -80805 -45817 -80761
rect -45773 -80805 -45717 -80761
rect -45673 -80805 -45617 -80761
rect -45573 -80805 -45517 -80761
rect -45473 -80805 -45417 -80761
rect -45373 -80805 -45317 -80761
rect -45273 -80805 -45217 -80761
rect -45173 -80805 -45117 -80761
rect -45073 -80805 -45017 -80761
rect -44973 -80805 -44917 -80761
rect -44873 -80805 -44817 -80761
rect -44773 -80805 -44717 -80761
rect -44673 -80805 -44617 -80761
rect -44573 -80805 -44517 -80761
rect -44473 -80805 -44017 -80761
rect -43973 -80805 -43917 -80761
rect -43873 -80805 -43817 -80761
rect -43773 -80805 -43717 -80761
rect -43673 -80805 -43617 -80761
rect -43573 -80805 -43517 -80761
rect -43473 -80805 -43417 -80761
rect -43373 -80805 -43317 -80761
rect -43273 -80805 -43217 -80761
rect -43173 -80805 -43117 -80761
rect -43073 -80805 -43017 -80761
rect -42973 -80805 -42917 -80761
rect -42873 -80805 -42817 -80761
rect -42773 -80805 -42717 -80761
rect -42673 -80805 -42617 -80761
rect -42573 -80805 -42517 -80761
rect -42473 -80805 -42000 -80761
rect -50768 -80861 -42000 -80805
rect -50768 -80905 -50017 -80861
rect -49973 -80905 -49917 -80861
rect -49873 -80905 -49817 -80861
rect -49773 -80905 -49717 -80861
rect -49673 -80905 -49617 -80861
rect -49573 -80905 -49517 -80861
rect -49473 -80905 -49417 -80861
rect -49373 -80905 -49317 -80861
rect -49273 -80905 -49217 -80861
rect -49173 -80905 -49117 -80861
rect -49073 -80905 -49017 -80861
rect -48973 -80905 -48917 -80861
rect -48873 -80905 -48817 -80861
rect -48773 -80905 -48717 -80861
rect -48673 -80905 -48617 -80861
rect -48573 -80905 -48517 -80861
rect -48473 -80905 -48017 -80861
rect -47973 -80905 -47917 -80861
rect -47873 -80905 -47817 -80861
rect -47773 -80905 -47717 -80861
rect -47673 -80905 -47617 -80861
rect -47573 -80905 -47517 -80861
rect -47473 -80905 -47417 -80861
rect -47373 -80905 -47317 -80861
rect -47273 -80905 -47217 -80861
rect -47173 -80905 -47117 -80861
rect -47073 -80905 -47017 -80861
rect -46973 -80905 -46917 -80861
rect -46873 -80905 -46817 -80861
rect -46773 -80905 -46717 -80861
rect -46673 -80905 -46617 -80861
rect -46573 -80905 -46517 -80861
rect -46473 -80905 -46017 -80861
rect -45973 -80905 -45917 -80861
rect -45873 -80905 -45817 -80861
rect -45773 -80905 -45717 -80861
rect -45673 -80905 -45617 -80861
rect -45573 -80905 -45517 -80861
rect -45473 -80905 -45417 -80861
rect -45373 -80905 -45317 -80861
rect -45273 -80905 -45217 -80861
rect -45173 -80905 -45117 -80861
rect -45073 -80905 -45017 -80861
rect -44973 -80905 -44917 -80861
rect -44873 -80905 -44817 -80861
rect -44773 -80905 -44717 -80861
rect -44673 -80905 -44617 -80861
rect -44573 -80905 -44517 -80861
rect -44473 -80905 -44017 -80861
rect -43973 -80905 -43917 -80861
rect -43873 -80905 -43817 -80861
rect -43773 -80905 -43717 -80861
rect -43673 -80905 -43617 -80861
rect -43573 -80905 -43517 -80861
rect -43473 -80905 -43417 -80861
rect -43373 -80905 -43317 -80861
rect -43273 -80905 -43217 -80861
rect -43173 -80905 -43117 -80861
rect -43073 -80905 -43017 -80861
rect -42973 -80905 -42917 -80861
rect -42873 -80905 -42817 -80861
rect -42773 -80905 -42717 -80861
rect -42673 -80905 -42617 -80861
rect -42573 -80905 -42517 -80861
rect -42473 -80905 -42000 -80861
rect -50768 -80961 -42000 -80905
rect -50768 -81005 -50017 -80961
rect -49973 -81005 -49917 -80961
rect -49873 -81005 -49817 -80961
rect -49773 -81005 -49717 -80961
rect -49673 -81005 -49617 -80961
rect -49573 -81005 -49517 -80961
rect -49473 -81005 -49417 -80961
rect -49373 -81005 -49317 -80961
rect -49273 -81005 -49217 -80961
rect -49173 -81005 -49117 -80961
rect -49073 -81005 -49017 -80961
rect -48973 -81005 -48917 -80961
rect -48873 -81005 -48817 -80961
rect -48773 -81005 -48717 -80961
rect -48673 -81005 -48617 -80961
rect -48573 -81005 -48517 -80961
rect -48473 -81005 -48017 -80961
rect -47973 -81005 -47917 -80961
rect -47873 -81005 -47817 -80961
rect -47773 -81005 -47717 -80961
rect -47673 -81005 -47617 -80961
rect -47573 -81005 -47517 -80961
rect -47473 -81005 -47417 -80961
rect -47373 -81005 -47317 -80961
rect -47273 -81005 -47217 -80961
rect -47173 -81005 -47117 -80961
rect -47073 -81005 -47017 -80961
rect -46973 -81005 -46917 -80961
rect -46873 -81005 -46817 -80961
rect -46773 -81005 -46717 -80961
rect -46673 -81005 -46617 -80961
rect -46573 -81005 -46517 -80961
rect -46473 -81005 -46017 -80961
rect -45973 -81005 -45917 -80961
rect -45873 -81005 -45817 -80961
rect -45773 -81005 -45717 -80961
rect -45673 -81005 -45617 -80961
rect -45573 -81005 -45517 -80961
rect -45473 -81005 -45417 -80961
rect -45373 -81005 -45317 -80961
rect -45273 -81005 -45217 -80961
rect -45173 -81005 -45117 -80961
rect -45073 -81005 -45017 -80961
rect -44973 -81005 -44917 -80961
rect -44873 -81005 -44817 -80961
rect -44773 -81005 -44717 -80961
rect -44673 -81005 -44617 -80961
rect -44573 -81005 -44517 -80961
rect -44473 -81005 -44017 -80961
rect -43973 -81005 -43917 -80961
rect -43873 -81005 -43817 -80961
rect -43773 -81005 -43717 -80961
rect -43673 -81005 -43617 -80961
rect -43573 -81005 -43517 -80961
rect -43473 -81005 -43417 -80961
rect -43373 -81005 -43317 -80961
rect -43273 -81005 -43217 -80961
rect -43173 -81005 -43117 -80961
rect -43073 -81005 -43017 -80961
rect -42973 -81005 -42917 -80961
rect -42873 -81005 -42817 -80961
rect -42773 -81005 -42717 -80961
rect -42673 -81005 -42617 -80961
rect -42573 -81005 -42517 -80961
rect -42473 -81005 -42000 -80961
rect -50768 -81061 -42000 -81005
rect -50768 -81105 -50017 -81061
rect -49973 -81105 -49917 -81061
rect -49873 -81105 -49817 -81061
rect -49773 -81105 -49717 -81061
rect -49673 -81105 -49617 -81061
rect -49573 -81105 -49517 -81061
rect -49473 -81105 -49417 -81061
rect -49373 -81105 -49317 -81061
rect -49273 -81105 -49217 -81061
rect -49173 -81105 -49117 -81061
rect -49073 -81105 -49017 -81061
rect -48973 -81105 -48917 -81061
rect -48873 -81105 -48817 -81061
rect -48773 -81105 -48717 -81061
rect -48673 -81105 -48617 -81061
rect -48573 -81105 -48517 -81061
rect -48473 -81105 -48017 -81061
rect -47973 -81105 -47917 -81061
rect -47873 -81105 -47817 -81061
rect -47773 -81105 -47717 -81061
rect -47673 -81105 -47617 -81061
rect -47573 -81105 -47517 -81061
rect -47473 -81105 -47417 -81061
rect -47373 -81105 -47317 -81061
rect -47273 -81105 -47217 -81061
rect -47173 -81105 -47117 -81061
rect -47073 -81105 -47017 -81061
rect -46973 -81105 -46917 -81061
rect -46873 -81105 -46817 -81061
rect -46773 -81105 -46717 -81061
rect -46673 -81105 -46617 -81061
rect -46573 -81105 -46517 -81061
rect -46473 -81105 -46017 -81061
rect -45973 -81105 -45917 -81061
rect -45873 -81105 -45817 -81061
rect -45773 -81105 -45717 -81061
rect -45673 -81105 -45617 -81061
rect -45573 -81105 -45517 -81061
rect -45473 -81105 -45417 -81061
rect -45373 -81105 -45317 -81061
rect -45273 -81105 -45217 -81061
rect -45173 -81105 -45117 -81061
rect -45073 -81105 -45017 -81061
rect -44973 -81105 -44917 -81061
rect -44873 -81105 -44817 -81061
rect -44773 -81105 -44717 -81061
rect -44673 -81105 -44617 -81061
rect -44573 -81105 -44517 -81061
rect -44473 -81105 -44017 -81061
rect -43973 -81105 -43917 -81061
rect -43873 -81105 -43817 -81061
rect -43773 -81105 -43717 -81061
rect -43673 -81105 -43617 -81061
rect -43573 -81105 -43517 -81061
rect -43473 -81105 -43417 -81061
rect -43373 -81105 -43317 -81061
rect -43273 -81105 -43217 -81061
rect -43173 -81105 -43117 -81061
rect -43073 -81105 -43017 -81061
rect -42973 -81105 -42917 -81061
rect -42873 -81105 -42817 -81061
rect -42773 -81105 -42717 -81061
rect -42673 -81105 -42617 -81061
rect -42573 -81105 -42517 -81061
rect -42473 -81105 -42000 -81061
rect -50768 -81161 -42000 -81105
rect -50768 -81205 -50017 -81161
rect -49973 -81205 -49917 -81161
rect -49873 -81205 -49817 -81161
rect -49773 -81205 -49717 -81161
rect -49673 -81205 -49617 -81161
rect -49573 -81205 -49517 -81161
rect -49473 -81205 -49417 -81161
rect -49373 -81205 -49317 -81161
rect -49273 -81205 -49217 -81161
rect -49173 -81205 -49117 -81161
rect -49073 -81205 -49017 -81161
rect -48973 -81205 -48917 -81161
rect -48873 -81205 -48817 -81161
rect -48773 -81205 -48717 -81161
rect -48673 -81205 -48617 -81161
rect -48573 -81205 -48517 -81161
rect -48473 -81205 -48017 -81161
rect -47973 -81205 -47917 -81161
rect -47873 -81205 -47817 -81161
rect -47773 -81205 -47717 -81161
rect -47673 -81205 -47617 -81161
rect -47573 -81205 -47517 -81161
rect -47473 -81205 -47417 -81161
rect -47373 -81205 -47317 -81161
rect -47273 -81205 -47217 -81161
rect -47173 -81205 -47117 -81161
rect -47073 -81205 -47017 -81161
rect -46973 -81205 -46917 -81161
rect -46873 -81205 -46817 -81161
rect -46773 -81205 -46717 -81161
rect -46673 -81205 -46617 -81161
rect -46573 -81205 -46517 -81161
rect -46473 -81205 -46017 -81161
rect -45973 -81205 -45917 -81161
rect -45873 -81205 -45817 -81161
rect -45773 -81205 -45717 -81161
rect -45673 -81205 -45617 -81161
rect -45573 -81205 -45517 -81161
rect -45473 -81205 -45417 -81161
rect -45373 -81205 -45317 -81161
rect -45273 -81205 -45217 -81161
rect -45173 -81205 -45117 -81161
rect -45073 -81205 -45017 -81161
rect -44973 -81205 -44917 -81161
rect -44873 -81205 -44817 -81161
rect -44773 -81205 -44717 -81161
rect -44673 -81205 -44617 -81161
rect -44573 -81205 -44517 -81161
rect -44473 -81205 -44017 -81161
rect -43973 -81205 -43917 -81161
rect -43873 -81205 -43817 -81161
rect -43773 -81205 -43717 -81161
rect -43673 -81205 -43617 -81161
rect -43573 -81205 -43517 -81161
rect -43473 -81205 -43417 -81161
rect -43373 -81205 -43317 -81161
rect -43273 -81205 -43217 -81161
rect -43173 -81205 -43117 -81161
rect -43073 -81205 -43017 -81161
rect -42973 -81205 -42917 -81161
rect -42873 -81205 -42817 -81161
rect -42773 -81205 -42717 -81161
rect -42673 -81205 -42617 -81161
rect -42573 -81205 -42517 -81161
rect -42473 -81205 -42000 -81161
rect -50768 -81261 -42000 -81205
rect -50768 -81305 -50017 -81261
rect -49973 -81305 -49917 -81261
rect -49873 -81305 -49817 -81261
rect -49773 -81305 -49717 -81261
rect -49673 -81305 -49617 -81261
rect -49573 -81305 -49517 -81261
rect -49473 -81305 -49417 -81261
rect -49373 -81305 -49317 -81261
rect -49273 -81305 -49217 -81261
rect -49173 -81305 -49117 -81261
rect -49073 -81305 -49017 -81261
rect -48973 -81305 -48917 -81261
rect -48873 -81305 -48817 -81261
rect -48773 -81305 -48717 -81261
rect -48673 -81305 -48617 -81261
rect -48573 -81305 -48517 -81261
rect -48473 -81305 -48017 -81261
rect -47973 -81305 -47917 -81261
rect -47873 -81305 -47817 -81261
rect -47773 -81305 -47717 -81261
rect -47673 -81305 -47617 -81261
rect -47573 -81305 -47517 -81261
rect -47473 -81305 -47417 -81261
rect -47373 -81305 -47317 -81261
rect -47273 -81305 -47217 -81261
rect -47173 -81305 -47117 -81261
rect -47073 -81305 -47017 -81261
rect -46973 -81305 -46917 -81261
rect -46873 -81305 -46817 -81261
rect -46773 -81305 -46717 -81261
rect -46673 -81305 -46617 -81261
rect -46573 -81305 -46517 -81261
rect -46473 -81305 -46017 -81261
rect -45973 -81305 -45917 -81261
rect -45873 -81305 -45817 -81261
rect -45773 -81305 -45717 -81261
rect -45673 -81305 -45617 -81261
rect -45573 -81305 -45517 -81261
rect -45473 -81305 -45417 -81261
rect -45373 -81305 -45317 -81261
rect -45273 -81305 -45217 -81261
rect -45173 -81305 -45117 -81261
rect -45073 -81305 -45017 -81261
rect -44973 -81305 -44917 -81261
rect -44873 -81305 -44817 -81261
rect -44773 -81305 -44717 -81261
rect -44673 -81305 -44617 -81261
rect -44573 -81305 -44517 -81261
rect -44473 -81305 -44017 -81261
rect -43973 -81305 -43917 -81261
rect -43873 -81305 -43817 -81261
rect -43773 -81305 -43717 -81261
rect -43673 -81305 -43617 -81261
rect -43573 -81305 -43517 -81261
rect -43473 -81305 -43417 -81261
rect -43373 -81305 -43317 -81261
rect -43273 -81305 -43217 -81261
rect -43173 -81305 -43117 -81261
rect -43073 -81305 -43017 -81261
rect -42973 -81305 -42917 -81261
rect -42873 -81305 -42817 -81261
rect -42773 -81305 -42717 -81261
rect -42673 -81305 -42617 -81261
rect -42573 -81305 -42517 -81261
rect -42473 -81305 -42000 -81261
rect -50768 -81361 -42000 -81305
rect -50768 -81405 -50017 -81361
rect -49973 -81405 -49917 -81361
rect -49873 -81405 -49817 -81361
rect -49773 -81405 -49717 -81361
rect -49673 -81405 -49617 -81361
rect -49573 -81405 -49517 -81361
rect -49473 -81405 -49417 -81361
rect -49373 -81405 -49317 -81361
rect -49273 -81405 -49217 -81361
rect -49173 -81405 -49117 -81361
rect -49073 -81405 -49017 -81361
rect -48973 -81405 -48917 -81361
rect -48873 -81405 -48817 -81361
rect -48773 -81405 -48717 -81361
rect -48673 -81405 -48617 -81361
rect -48573 -81405 -48517 -81361
rect -48473 -81405 -48017 -81361
rect -47973 -81405 -47917 -81361
rect -47873 -81405 -47817 -81361
rect -47773 -81405 -47717 -81361
rect -47673 -81405 -47617 -81361
rect -47573 -81405 -47517 -81361
rect -47473 -81405 -47417 -81361
rect -47373 -81405 -47317 -81361
rect -47273 -81405 -47217 -81361
rect -47173 -81405 -47117 -81361
rect -47073 -81405 -47017 -81361
rect -46973 -81405 -46917 -81361
rect -46873 -81405 -46817 -81361
rect -46773 -81405 -46717 -81361
rect -46673 -81405 -46617 -81361
rect -46573 -81405 -46517 -81361
rect -46473 -81405 -46017 -81361
rect -45973 -81405 -45917 -81361
rect -45873 -81405 -45817 -81361
rect -45773 -81405 -45717 -81361
rect -45673 -81405 -45617 -81361
rect -45573 -81405 -45517 -81361
rect -45473 -81405 -45417 -81361
rect -45373 -81405 -45317 -81361
rect -45273 -81405 -45217 -81361
rect -45173 -81405 -45117 -81361
rect -45073 -81405 -45017 -81361
rect -44973 -81405 -44917 -81361
rect -44873 -81405 -44817 -81361
rect -44773 -81405 -44717 -81361
rect -44673 -81405 -44617 -81361
rect -44573 -81405 -44517 -81361
rect -44473 -81405 -44017 -81361
rect -43973 -81405 -43917 -81361
rect -43873 -81405 -43817 -81361
rect -43773 -81405 -43717 -81361
rect -43673 -81405 -43617 -81361
rect -43573 -81405 -43517 -81361
rect -43473 -81405 -43417 -81361
rect -43373 -81405 -43317 -81361
rect -43273 -81405 -43217 -81361
rect -43173 -81405 -43117 -81361
rect -43073 -81405 -43017 -81361
rect -42973 -81405 -42917 -81361
rect -42873 -81405 -42817 -81361
rect -42773 -81405 -42717 -81361
rect -42673 -81405 -42617 -81361
rect -42573 -81405 -42517 -81361
rect -42473 -81405 -42000 -81361
rect -50768 -81461 -42000 -81405
rect -50768 -81505 -50017 -81461
rect -49973 -81505 -49917 -81461
rect -49873 -81505 -49817 -81461
rect -49773 -81505 -49717 -81461
rect -49673 -81505 -49617 -81461
rect -49573 -81505 -49517 -81461
rect -49473 -81505 -49417 -81461
rect -49373 -81505 -49317 -81461
rect -49273 -81505 -49217 -81461
rect -49173 -81505 -49117 -81461
rect -49073 -81505 -49017 -81461
rect -48973 -81505 -48917 -81461
rect -48873 -81505 -48817 -81461
rect -48773 -81505 -48717 -81461
rect -48673 -81505 -48617 -81461
rect -48573 -81505 -48517 -81461
rect -48473 -81505 -48017 -81461
rect -47973 -81505 -47917 -81461
rect -47873 -81505 -47817 -81461
rect -47773 -81505 -47717 -81461
rect -47673 -81505 -47617 -81461
rect -47573 -81505 -47517 -81461
rect -47473 -81505 -47417 -81461
rect -47373 -81505 -47317 -81461
rect -47273 -81505 -47217 -81461
rect -47173 -81505 -47117 -81461
rect -47073 -81505 -47017 -81461
rect -46973 -81505 -46917 -81461
rect -46873 -81505 -46817 -81461
rect -46773 -81505 -46717 -81461
rect -46673 -81505 -46617 -81461
rect -46573 -81505 -46517 -81461
rect -46473 -81505 -46017 -81461
rect -45973 -81505 -45917 -81461
rect -45873 -81505 -45817 -81461
rect -45773 -81505 -45717 -81461
rect -45673 -81505 -45617 -81461
rect -45573 -81505 -45517 -81461
rect -45473 -81505 -45417 -81461
rect -45373 -81505 -45317 -81461
rect -45273 -81505 -45217 -81461
rect -45173 -81505 -45117 -81461
rect -45073 -81505 -45017 -81461
rect -44973 -81505 -44917 -81461
rect -44873 -81505 -44817 -81461
rect -44773 -81505 -44717 -81461
rect -44673 -81505 -44617 -81461
rect -44573 -81505 -44517 -81461
rect -44473 -81505 -44017 -81461
rect -43973 -81505 -43917 -81461
rect -43873 -81505 -43817 -81461
rect -43773 -81505 -43717 -81461
rect -43673 -81505 -43617 -81461
rect -43573 -81505 -43517 -81461
rect -43473 -81505 -43417 -81461
rect -43373 -81505 -43317 -81461
rect -43273 -81505 -43217 -81461
rect -43173 -81505 -43117 -81461
rect -43073 -81505 -43017 -81461
rect -42973 -81505 -42917 -81461
rect -42873 -81505 -42817 -81461
rect -42773 -81505 -42717 -81461
rect -42673 -81505 -42617 -81461
rect -42573 -81505 -42517 -81461
rect -42473 -81505 -42000 -81461
rect -50768 -81561 -42000 -81505
rect -50768 -81605 -50017 -81561
rect -49973 -81605 -49917 -81561
rect -49873 -81605 -49817 -81561
rect -49773 -81605 -49717 -81561
rect -49673 -81605 -49617 -81561
rect -49573 -81605 -49517 -81561
rect -49473 -81605 -49417 -81561
rect -49373 -81605 -49317 -81561
rect -49273 -81605 -49217 -81561
rect -49173 -81605 -49117 -81561
rect -49073 -81605 -49017 -81561
rect -48973 -81605 -48917 -81561
rect -48873 -81605 -48817 -81561
rect -48773 -81605 -48717 -81561
rect -48673 -81605 -48617 -81561
rect -48573 -81605 -48517 -81561
rect -48473 -81605 -48017 -81561
rect -47973 -81605 -47917 -81561
rect -47873 -81605 -47817 -81561
rect -47773 -81605 -47717 -81561
rect -47673 -81605 -47617 -81561
rect -47573 -81605 -47517 -81561
rect -47473 -81605 -47417 -81561
rect -47373 -81605 -47317 -81561
rect -47273 -81605 -47217 -81561
rect -47173 -81605 -47117 -81561
rect -47073 -81605 -47017 -81561
rect -46973 -81605 -46917 -81561
rect -46873 -81605 -46817 -81561
rect -46773 -81605 -46717 -81561
rect -46673 -81605 -46617 -81561
rect -46573 -81605 -46517 -81561
rect -46473 -81605 -46017 -81561
rect -45973 -81605 -45917 -81561
rect -45873 -81605 -45817 -81561
rect -45773 -81605 -45717 -81561
rect -45673 -81605 -45617 -81561
rect -45573 -81605 -45517 -81561
rect -45473 -81605 -45417 -81561
rect -45373 -81605 -45317 -81561
rect -45273 -81605 -45217 -81561
rect -45173 -81605 -45117 -81561
rect -45073 -81605 -45017 -81561
rect -44973 -81605 -44917 -81561
rect -44873 -81605 -44817 -81561
rect -44773 -81605 -44717 -81561
rect -44673 -81605 -44617 -81561
rect -44573 -81605 -44517 -81561
rect -44473 -81605 -44017 -81561
rect -43973 -81605 -43917 -81561
rect -43873 -81605 -43817 -81561
rect -43773 -81605 -43717 -81561
rect -43673 -81605 -43617 -81561
rect -43573 -81605 -43517 -81561
rect -43473 -81605 -43417 -81561
rect -43373 -81605 -43317 -81561
rect -43273 -81605 -43217 -81561
rect -43173 -81605 -43117 -81561
rect -43073 -81605 -43017 -81561
rect -42973 -81605 -42917 -81561
rect -42873 -81605 -42817 -81561
rect -42773 -81605 -42717 -81561
rect -42673 -81605 -42617 -81561
rect -42573 -81605 -42517 -81561
rect -42473 -81605 -42000 -81561
rect -50768 -81661 -42000 -81605
rect -50768 -81705 -50017 -81661
rect -49973 -81705 -49917 -81661
rect -49873 -81705 -49817 -81661
rect -49773 -81705 -49717 -81661
rect -49673 -81705 -49617 -81661
rect -49573 -81705 -49517 -81661
rect -49473 -81705 -49417 -81661
rect -49373 -81705 -49317 -81661
rect -49273 -81705 -49217 -81661
rect -49173 -81705 -49117 -81661
rect -49073 -81705 -49017 -81661
rect -48973 -81705 -48917 -81661
rect -48873 -81705 -48817 -81661
rect -48773 -81705 -48717 -81661
rect -48673 -81705 -48617 -81661
rect -48573 -81705 -48517 -81661
rect -48473 -81705 -48017 -81661
rect -47973 -81705 -47917 -81661
rect -47873 -81705 -47817 -81661
rect -47773 -81705 -47717 -81661
rect -47673 -81705 -47617 -81661
rect -47573 -81705 -47517 -81661
rect -47473 -81705 -47417 -81661
rect -47373 -81705 -47317 -81661
rect -47273 -81705 -47217 -81661
rect -47173 -81705 -47117 -81661
rect -47073 -81705 -47017 -81661
rect -46973 -81705 -46917 -81661
rect -46873 -81705 -46817 -81661
rect -46773 -81705 -46717 -81661
rect -46673 -81705 -46617 -81661
rect -46573 -81705 -46517 -81661
rect -46473 -81705 -46017 -81661
rect -45973 -81705 -45917 -81661
rect -45873 -81705 -45817 -81661
rect -45773 -81705 -45717 -81661
rect -45673 -81705 -45617 -81661
rect -45573 -81705 -45517 -81661
rect -45473 -81705 -45417 -81661
rect -45373 -81705 -45317 -81661
rect -45273 -81705 -45217 -81661
rect -45173 -81705 -45117 -81661
rect -45073 -81705 -45017 -81661
rect -44973 -81705 -44917 -81661
rect -44873 -81705 -44817 -81661
rect -44773 -81705 -44717 -81661
rect -44673 -81705 -44617 -81661
rect -44573 -81705 -44517 -81661
rect -44473 -81705 -44017 -81661
rect -43973 -81705 -43917 -81661
rect -43873 -81705 -43817 -81661
rect -43773 -81705 -43717 -81661
rect -43673 -81705 -43617 -81661
rect -43573 -81705 -43517 -81661
rect -43473 -81705 -43417 -81661
rect -43373 -81705 -43317 -81661
rect -43273 -81705 -43217 -81661
rect -43173 -81705 -43117 -81661
rect -43073 -81705 -43017 -81661
rect -42973 -81705 -42917 -81661
rect -42873 -81705 -42817 -81661
rect -42773 -81705 -42717 -81661
rect -42673 -81705 -42617 -81661
rect -42573 -81705 -42517 -81661
rect -42473 -81705 -42000 -81661
rect -50768 -81761 -42000 -81705
rect -50768 -81805 -50017 -81761
rect -49973 -81805 -49917 -81761
rect -49873 -81805 -49817 -81761
rect -49773 -81805 -49717 -81761
rect -49673 -81805 -49617 -81761
rect -49573 -81805 -49517 -81761
rect -49473 -81805 -49417 -81761
rect -49373 -81805 -49317 -81761
rect -49273 -81805 -49217 -81761
rect -49173 -81805 -49117 -81761
rect -49073 -81805 -49017 -81761
rect -48973 -81805 -48917 -81761
rect -48873 -81805 -48817 -81761
rect -48773 -81805 -48717 -81761
rect -48673 -81805 -48617 -81761
rect -48573 -81805 -48517 -81761
rect -48473 -81805 -48017 -81761
rect -47973 -81805 -47917 -81761
rect -47873 -81805 -47817 -81761
rect -47773 -81805 -47717 -81761
rect -47673 -81805 -47617 -81761
rect -47573 -81805 -47517 -81761
rect -47473 -81805 -47417 -81761
rect -47373 -81805 -47317 -81761
rect -47273 -81805 -47217 -81761
rect -47173 -81805 -47117 -81761
rect -47073 -81805 -47017 -81761
rect -46973 -81805 -46917 -81761
rect -46873 -81805 -46817 -81761
rect -46773 -81805 -46717 -81761
rect -46673 -81805 -46617 -81761
rect -46573 -81805 -46517 -81761
rect -46473 -81805 -46017 -81761
rect -45973 -81805 -45917 -81761
rect -45873 -81805 -45817 -81761
rect -45773 -81805 -45717 -81761
rect -45673 -81805 -45617 -81761
rect -45573 -81805 -45517 -81761
rect -45473 -81805 -45417 -81761
rect -45373 -81805 -45317 -81761
rect -45273 -81805 -45217 -81761
rect -45173 -81805 -45117 -81761
rect -45073 -81805 -45017 -81761
rect -44973 -81805 -44917 -81761
rect -44873 -81805 -44817 -81761
rect -44773 -81805 -44717 -81761
rect -44673 -81805 -44617 -81761
rect -44573 -81805 -44517 -81761
rect -44473 -81805 -44017 -81761
rect -43973 -81805 -43917 -81761
rect -43873 -81805 -43817 -81761
rect -43773 -81805 -43717 -81761
rect -43673 -81805 -43617 -81761
rect -43573 -81805 -43517 -81761
rect -43473 -81805 -43417 -81761
rect -43373 -81805 -43317 -81761
rect -43273 -81805 -43217 -81761
rect -43173 -81805 -43117 -81761
rect -43073 -81805 -43017 -81761
rect -42973 -81805 -42917 -81761
rect -42873 -81805 -42817 -81761
rect -42773 -81805 -42717 -81761
rect -42673 -81805 -42617 -81761
rect -42573 -81805 -42517 -81761
rect -42473 -81805 -42000 -81761
rect -50768 -81861 -42000 -81805
rect -50768 -81905 -50017 -81861
rect -49973 -81905 -49917 -81861
rect -49873 -81905 -49817 -81861
rect -49773 -81905 -49717 -81861
rect -49673 -81905 -49617 -81861
rect -49573 -81905 -49517 -81861
rect -49473 -81905 -49417 -81861
rect -49373 -81905 -49317 -81861
rect -49273 -81905 -49217 -81861
rect -49173 -81905 -49117 -81861
rect -49073 -81905 -49017 -81861
rect -48973 -81905 -48917 -81861
rect -48873 -81905 -48817 -81861
rect -48773 -81905 -48717 -81861
rect -48673 -81905 -48617 -81861
rect -48573 -81905 -48517 -81861
rect -48473 -81905 -48017 -81861
rect -47973 -81905 -47917 -81861
rect -47873 -81905 -47817 -81861
rect -47773 -81905 -47717 -81861
rect -47673 -81905 -47617 -81861
rect -47573 -81905 -47517 -81861
rect -47473 -81905 -47417 -81861
rect -47373 -81905 -47317 -81861
rect -47273 -81905 -47217 -81861
rect -47173 -81905 -47117 -81861
rect -47073 -81905 -47017 -81861
rect -46973 -81905 -46917 -81861
rect -46873 -81905 -46817 -81861
rect -46773 -81905 -46717 -81861
rect -46673 -81905 -46617 -81861
rect -46573 -81905 -46517 -81861
rect -46473 -81905 -46017 -81861
rect -45973 -81905 -45917 -81861
rect -45873 -81905 -45817 -81861
rect -45773 -81905 -45717 -81861
rect -45673 -81905 -45617 -81861
rect -45573 -81905 -45517 -81861
rect -45473 -81905 -45417 -81861
rect -45373 -81905 -45317 -81861
rect -45273 -81905 -45217 -81861
rect -45173 -81905 -45117 -81861
rect -45073 -81905 -45017 -81861
rect -44973 -81905 -44917 -81861
rect -44873 -81905 -44817 -81861
rect -44773 -81905 -44717 -81861
rect -44673 -81905 -44617 -81861
rect -44573 -81905 -44517 -81861
rect -44473 -81905 -44017 -81861
rect -43973 -81905 -43917 -81861
rect -43873 -81905 -43817 -81861
rect -43773 -81905 -43717 -81861
rect -43673 -81905 -43617 -81861
rect -43573 -81905 -43517 -81861
rect -43473 -81905 -43417 -81861
rect -43373 -81905 -43317 -81861
rect -43273 -81905 -43217 -81861
rect -43173 -81905 -43117 -81861
rect -43073 -81905 -43017 -81861
rect -42973 -81905 -42917 -81861
rect -42873 -81905 -42817 -81861
rect -42773 -81905 -42717 -81861
rect -42673 -81905 -42617 -81861
rect -42573 -81905 -42517 -81861
rect -42473 -81905 -42000 -81861
rect -50768 -81961 -42000 -81905
rect -50768 -82005 -50017 -81961
rect -49973 -82005 -49917 -81961
rect -49873 -82005 -49817 -81961
rect -49773 -82005 -49717 -81961
rect -49673 -82005 -49617 -81961
rect -49573 -82005 -49517 -81961
rect -49473 -82005 -49417 -81961
rect -49373 -82005 -49317 -81961
rect -49273 -82005 -49217 -81961
rect -49173 -82005 -49117 -81961
rect -49073 -82005 -49017 -81961
rect -48973 -82005 -48917 -81961
rect -48873 -82005 -48817 -81961
rect -48773 -82005 -48717 -81961
rect -48673 -82005 -48617 -81961
rect -48573 -82005 -48517 -81961
rect -48473 -82005 -48017 -81961
rect -47973 -82005 -47917 -81961
rect -47873 -82005 -47817 -81961
rect -47773 -82005 -47717 -81961
rect -47673 -82005 -47617 -81961
rect -47573 -82005 -47517 -81961
rect -47473 -82005 -47417 -81961
rect -47373 -82005 -47317 -81961
rect -47273 -82005 -47217 -81961
rect -47173 -82005 -47117 -81961
rect -47073 -82005 -47017 -81961
rect -46973 -82005 -46917 -81961
rect -46873 -82005 -46817 -81961
rect -46773 -82005 -46717 -81961
rect -46673 -82005 -46617 -81961
rect -46573 -82005 -46517 -81961
rect -46473 -82005 -46017 -81961
rect -45973 -82005 -45917 -81961
rect -45873 -82005 -45817 -81961
rect -45773 -82005 -45717 -81961
rect -45673 -82005 -45617 -81961
rect -45573 -82005 -45517 -81961
rect -45473 -82005 -45417 -81961
rect -45373 -82005 -45317 -81961
rect -45273 -82005 -45217 -81961
rect -45173 -82005 -45117 -81961
rect -45073 -82005 -45017 -81961
rect -44973 -82005 -44917 -81961
rect -44873 -82005 -44817 -81961
rect -44773 -82005 -44717 -81961
rect -44673 -82005 -44617 -81961
rect -44573 -82005 -44517 -81961
rect -44473 -82005 -44017 -81961
rect -43973 -82005 -43917 -81961
rect -43873 -82005 -43817 -81961
rect -43773 -82005 -43717 -81961
rect -43673 -82005 -43617 -81961
rect -43573 -82005 -43517 -81961
rect -43473 -82005 -43417 -81961
rect -43373 -82005 -43317 -81961
rect -43273 -82005 -43217 -81961
rect -43173 -82005 -43117 -81961
rect -43073 -82005 -43017 -81961
rect -42973 -82005 -42917 -81961
rect -42873 -82005 -42817 -81961
rect -42773 -82005 -42717 -81961
rect -42673 -82005 -42617 -81961
rect -42573 -82005 -42517 -81961
rect -42473 -82005 -42000 -81961
rect -50768 -106193 -42000 -82005
rect -50768 -106237 -50075 -106193
rect -50031 -106237 -49975 -106193
rect -49931 -106237 -49875 -106193
rect -49831 -106237 -49775 -106193
rect -49731 -106237 -49675 -106193
rect -49631 -106237 -49575 -106193
rect -49531 -106237 -49475 -106193
rect -49431 -106237 -49375 -106193
rect -49331 -106237 -49275 -106193
rect -49231 -106237 -49175 -106193
rect -49131 -106237 -49075 -106193
rect -49031 -106237 -48975 -106193
rect -48931 -106237 -48875 -106193
rect -48831 -106237 -48775 -106193
rect -48731 -106237 -48675 -106193
rect -48631 -106237 -48575 -106193
rect -48531 -106237 -48075 -106193
rect -48031 -106237 -47975 -106193
rect -47931 -106237 -47875 -106193
rect -47831 -106237 -47775 -106193
rect -47731 -106237 -47675 -106193
rect -47631 -106237 -47575 -106193
rect -47531 -106237 -47475 -106193
rect -47431 -106237 -47375 -106193
rect -47331 -106237 -47275 -106193
rect -47231 -106237 -47175 -106193
rect -47131 -106237 -47075 -106193
rect -47031 -106237 -46975 -106193
rect -46931 -106237 -46875 -106193
rect -46831 -106237 -46775 -106193
rect -46731 -106237 -46675 -106193
rect -46631 -106237 -46575 -106193
rect -46531 -106237 -46075 -106193
rect -46031 -106237 -45975 -106193
rect -45931 -106237 -45875 -106193
rect -45831 -106237 -45775 -106193
rect -45731 -106237 -45675 -106193
rect -45631 -106237 -45575 -106193
rect -45531 -106237 -45475 -106193
rect -45431 -106237 -45375 -106193
rect -45331 -106237 -45275 -106193
rect -45231 -106237 -45175 -106193
rect -45131 -106237 -45075 -106193
rect -45031 -106237 -44975 -106193
rect -44931 -106237 -44875 -106193
rect -44831 -106237 -44775 -106193
rect -44731 -106237 -44675 -106193
rect -44631 -106237 -44575 -106193
rect -44531 -106237 -44075 -106193
rect -44031 -106237 -43975 -106193
rect -43931 -106237 -43875 -106193
rect -43831 -106237 -43775 -106193
rect -43731 -106237 -43675 -106193
rect -43631 -106237 -43575 -106193
rect -43531 -106237 -43475 -106193
rect -43431 -106237 -43375 -106193
rect -43331 -106237 -43275 -106193
rect -43231 -106237 -43175 -106193
rect -43131 -106237 -43075 -106193
rect -43031 -106237 -42975 -106193
rect -42931 -106237 -42875 -106193
rect -42831 -106237 -42775 -106193
rect -42731 -106237 -42675 -106193
rect -42631 -106237 -42575 -106193
rect -42531 -106237 -42000 -106193
rect -50768 -106293 -42000 -106237
rect -50768 -106337 -50075 -106293
rect -50031 -106337 -49975 -106293
rect -49931 -106337 -49875 -106293
rect -49831 -106337 -49775 -106293
rect -49731 -106337 -49675 -106293
rect -49631 -106337 -49575 -106293
rect -49531 -106337 -49475 -106293
rect -49431 -106337 -49375 -106293
rect -49331 -106337 -49275 -106293
rect -49231 -106337 -49175 -106293
rect -49131 -106337 -49075 -106293
rect -49031 -106337 -48975 -106293
rect -48931 -106337 -48875 -106293
rect -48831 -106337 -48775 -106293
rect -48731 -106337 -48675 -106293
rect -48631 -106337 -48575 -106293
rect -48531 -106337 -48075 -106293
rect -48031 -106337 -47975 -106293
rect -47931 -106337 -47875 -106293
rect -47831 -106337 -47775 -106293
rect -47731 -106337 -47675 -106293
rect -47631 -106337 -47575 -106293
rect -47531 -106337 -47475 -106293
rect -47431 -106337 -47375 -106293
rect -47331 -106337 -47275 -106293
rect -47231 -106337 -47175 -106293
rect -47131 -106337 -47075 -106293
rect -47031 -106337 -46975 -106293
rect -46931 -106337 -46875 -106293
rect -46831 -106337 -46775 -106293
rect -46731 -106337 -46675 -106293
rect -46631 -106337 -46575 -106293
rect -46531 -106337 -46075 -106293
rect -46031 -106337 -45975 -106293
rect -45931 -106337 -45875 -106293
rect -45831 -106337 -45775 -106293
rect -45731 -106337 -45675 -106293
rect -45631 -106337 -45575 -106293
rect -45531 -106337 -45475 -106293
rect -45431 -106337 -45375 -106293
rect -45331 -106337 -45275 -106293
rect -45231 -106337 -45175 -106293
rect -45131 -106337 -45075 -106293
rect -45031 -106337 -44975 -106293
rect -44931 -106337 -44875 -106293
rect -44831 -106337 -44775 -106293
rect -44731 -106337 -44675 -106293
rect -44631 -106337 -44575 -106293
rect -44531 -106337 -44075 -106293
rect -44031 -106337 -43975 -106293
rect -43931 -106337 -43875 -106293
rect -43831 -106337 -43775 -106293
rect -43731 -106337 -43675 -106293
rect -43631 -106337 -43575 -106293
rect -43531 -106337 -43475 -106293
rect -43431 -106337 -43375 -106293
rect -43331 -106337 -43275 -106293
rect -43231 -106337 -43175 -106293
rect -43131 -106337 -43075 -106293
rect -43031 -106337 -42975 -106293
rect -42931 -106337 -42875 -106293
rect -42831 -106337 -42775 -106293
rect -42731 -106337 -42675 -106293
rect -42631 -106337 -42575 -106293
rect -42531 -106337 -42000 -106293
rect -50768 -106393 -42000 -106337
rect -50768 -106437 -50075 -106393
rect -50031 -106437 -49975 -106393
rect -49931 -106437 -49875 -106393
rect -49831 -106437 -49775 -106393
rect -49731 -106437 -49675 -106393
rect -49631 -106437 -49575 -106393
rect -49531 -106437 -49475 -106393
rect -49431 -106437 -49375 -106393
rect -49331 -106437 -49275 -106393
rect -49231 -106437 -49175 -106393
rect -49131 -106437 -49075 -106393
rect -49031 -106437 -48975 -106393
rect -48931 -106437 -48875 -106393
rect -48831 -106437 -48775 -106393
rect -48731 -106437 -48675 -106393
rect -48631 -106437 -48575 -106393
rect -48531 -106437 -48075 -106393
rect -48031 -106437 -47975 -106393
rect -47931 -106437 -47875 -106393
rect -47831 -106437 -47775 -106393
rect -47731 -106437 -47675 -106393
rect -47631 -106437 -47575 -106393
rect -47531 -106437 -47475 -106393
rect -47431 -106437 -47375 -106393
rect -47331 -106437 -47275 -106393
rect -47231 -106437 -47175 -106393
rect -47131 -106437 -47075 -106393
rect -47031 -106437 -46975 -106393
rect -46931 -106437 -46875 -106393
rect -46831 -106437 -46775 -106393
rect -46731 -106437 -46675 -106393
rect -46631 -106437 -46575 -106393
rect -46531 -106437 -46075 -106393
rect -46031 -106437 -45975 -106393
rect -45931 -106437 -45875 -106393
rect -45831 -106437 -45775 -106393
rect -45731 -106437 -45675 -106393
rect -45631 -106437 -45575 -106393
rect -45531 -106437 -45475 -106393
rect -45431 -106437 -45375 -106393
rect -45331 -106437 -45275 -106393
rect -45231 -106437 -45175 -106393
rect -45131 -106437 -45075 -106393
rect -45031 -106437 -44975 -106393
rect -44931 -106437 -44875 -106393
rect -44831 -106437 -44775 -106393
rect -44731 -106437 -44675 -106393
rect -44631 -106437 -44575 -106393
rect -44531 -106437 -44075 -106393
rect -44031 -106437 -43975 -106393
rect -43931 -106437 -43875 -106393
rect -43831 -106437 -43775 -106393
rect -43731 -106437 -43675 -106393
rect -43631 -106437 -43575 -106393
rect -43531 -106437 -43475 -106393
rect -43431 -106437 -43375 -106393
rect -43331 -106437 -43275 -106393
rect -43231 -106437 -43175 -106393
rect -43131 -106437 -43075 -106393
rect -43031 -106437 -42975 -106393
rect -42931 -106437 -42875 -106393
rect -42831 -106437 -42775 -106393
rect -42731 -106437 -42675 -106393
rect -42631 -106437 -42575 -106393
rect -42531 -106437 -42000 -106393
rect -50768 -106493 -42000 -106437
rect -50768 -106537 -50075 -106493
rect -50031 -106537 -49975 -106493
rect -49931 -106537 -49875 -106493
rect -49831 -106537 -49775 -106493
rect -49731 -106537 -49675 -106493
rect -49631 -106537 -49575 -106493
rect -49531 -106537 -49475 -106493
rect -49431 -106537 -49375 -106493
rect -49331 -106537 -49275 -106493
rect -49231 -106537 -49175 -106493
rect -49131 -106537 -49075 -106493
rect -49031 -106537 -48975 -106493
rect -48931 -106537 -48875 -106493
rect -48831 -106537 -48775 -106493
rect -48731 -106537 -48675 -106493
rect -48631 -106537 -48575 -106493
rect -48531 -106537 -48075 -106493
rect -48031 -106537 -47975 -106493
rect -47931 -106537 -47875 -106493
rect -47831 -106537 -47775 -106493
rect -47731 -106537 -47675 -106493
rect -47631 -106537 -47575 -106493
rect -47531 -106537 -47475 -106493
rect -47431 -106537 -47375 -106493
rect -47331 -106537 -47275 -106493
rect -47231 -106537 -47175 -106493
rect -47131 -106537 -47075 -106493
rect -47031 -106537 -46975 -106493
rect -46931 -106537 -46875 -106493
rect -46831 -106537 -46775 -106493
rect -46731 -106537 -46675 -106493
rect -46631 -106537 -46575 -106493
rect -46531 -106537 -46075 -106493
rect -46031 -106537 -45975 -106493
rect -45931 -106537 -45875 -106493
rect -45831 -106537 -45775 -106493
rect -45731 -106537 -45675 -106493
rect -45631 -106537 -45575 -106493
rect -45531 -106537 -45475 -106493
rect -45431 -106537 -45375 -106493
rect -45331 -106537 -45275 -106493
rect -45231 -106537 -45175 -106493
rect -45131 -106537 -45075 -106493
rect -45031 -106537 -44975 -106493
rect -44931 -106537 -44875 -106493
rect -44831 -106537 -44775 -106493
rect -44731 -106537 -44675 -106493
rect -44631 -106537 -44575 -106493
rect -44531 -106537 -44075 -106493
rect -44031 -106537 -43975 -106493
rect -43931 -106537 -43875 -106493
rect -43831 -106537 -43775 -106493
rect -43731 -106537 -43675 -106493
rect -43631 -106537 -43575 -106493
rect -43531 -106537 -43475 -106493
rect -43431 -106537 -43375 -106493
rect -43331 -106537 -43275 -106493
rect -43231 -106537 -43175 -106493
rect -43131 -106537 -43075 -106493
rect -43031 -106537 -42975 -106493
rect -42931 -106537 -42875 -106493
rect -42831 -106537 -42775 -106493
rect -42731 -106537 -42675 -106493
rect -42631 -106537 -42575 -106493
rect -42531 -106537 -42000 -106493
rect -50768 -106593 -42000 -106537
rect -50768 -106637 -50075 -106593
rect -50031 -106637 -49975 -106593
rect -49931 -106637 -49875 -106593
rect -49831 -106637 -49775 -106593
rect -49731 -106637 -49675 -106593
rect -49631 -106637 -49575 -106593
rect -49531 -106637 -49475 -106593
rect -49431 -106637 -49375 -106593
rect -49331 -106637 -49275 -106593
rect -49231 -106637 -49175 -106593
rect -49131 -106637 -49075 -106593
rect -49031 -106637 -48975 -106593
rect -48931 -106637 -48875 -106593
rect -48831 -106637 -48775 -106593
rect -48731 -106637 -48675 -106593
rect -48631 -106637 -48575 -106593
rect -48531 -106637 -48075 -106593
rect -48031 -106637 -47975 -106593
rect -47931 -106637 -47875 -106593
rect -47831 -106637 -47775 -106593
rect -47731 -106637 -47675 -106593
rect -47631 -106637 -47575 -106593
rect -47531 -106637 -47475 -106593
rect -47431 -106637 -47375 -106593
rect -47331 -106637 -47275 -106593
rect -47231 -106637 -47175 -106593
rect -47131 -106637 -47075 -106593
rect -47031 -106637 -46975 -106593
rect -46931 -106637 -46875 -106593
rect -46831 -106637 -46775 -106593
rect -46731 -106637 -46675 -106593
rect -46631 -106637 -46575 -106593
rect -46531 -106637 -46075 -106593
rect -46031 -106637 -45975 -106593
rect -45931 -106637 -45875 -106593
rect -45831 -106637 -45775 -106593
rect -45731 -106637 -45675 -106593
rect -45631 -106637 -45575 -106593
rect -45531 -106637 -45475 -106593
rect -45431 -106637 -45375 -106593
rect -45331 -106637 -45275 -106593
rect -45231 -106637 -45175 -106593
rect -45131 -106637 -45075 -106593
rect -45031 -106637 -44975 -106593
rect -44931 -106637 -44875 -106593
rect -44831 -106637 -44775 -106593
rect -44731 -106637 -44675 -106593
rect -44631 -106637 -44575 -106593
rect -44531 -106637 -44075 -106593
rect -44031 -106637 -43975 -106593
rect -43931 -106637 -43875 -106593
rect -43831 -106637 -43775 -106593
rect -43731 -106637 -43675 -106593
rect -43631 -106637 -43575 -106593
rect -43531 -106637 -43475 -106593
rect -43431 -106637 -43375 -106593
rect -43331 -106637 -43275 -106593
rect -43231 -106637 -43175 -106593
rect -43131 -106637 -43075 -106593
rect -43031 -106637 -42975 -106593
rect -42931 -106637 -42875 -106593
rect -42831 -106637 -42775 -106593
rect -42731 -106637 -42675 -106593
rect -42631 -106637 -42575 -106593
rect -42531 -106637 -42000 -106593
rect -50768 -106693 -42000 -106637
rect -50768 -106737 -50075 -106693
rect -50031 -106737 -49975 -106693
rect -49931 -106737 -49875 -106693
rect -49831 -106737 -49775 -106693
rect -49731 -106737 -49675 -106693
rect -49631 -106737 -49575 -106693
rect -49531 -106737 -49475 -106693
rect -49431 -106737 -49375 -106693
rect -49331 -106737 -49275 -106693
rect -49231 -106737 -49175 -106693
rect -49131 -106737 -49075 -106693
rect -49031 -106737 -48975 -106693
rect -48931 -106737 -48875 -106693
rect -48831 -106737 -48775 -106693
rect -48731 -106737 -48675 -106693
rect -48631 -106737 -48575 -106693
rect -48531 -106737 -48075 -106693
rect -48031 -106737 -47975 -106693
rect -47931 -106737 -47875 -106693
rect -47831 -106737 -47775 -106693
rect -47731 -106737 -47675 -106693
rect -47631 -106737 -47575 -106693
rect -47531 -106737 -47475 -106693
rect -47431 -106737 -47375 -106693
rect -47331 -106737 -47275 -106693
rect -47231 -106737 -47175 -106693
rect -47131 -106737 -47075 -106693
rect -47031 -106737 -46975 -106693
rect -46931 -106737 -46875 -106693
rect -46831 -106737 -46775 -106693
rect -46731 -106737 -46675 -106693
rect -46631 -106737 -46575 -106693
rect -46531 -106737 -46075 -106693
rect -46031 -106737 -45975 -106693
rect -45931 -106737 -45875 -106693
rect -45831 -106737 -45775 -106693
rect -45731 -106737 -45675 -106693
rect -45631 -106737 -45575 -106693
rect -45531 -106737 -45475 -106693
rect -45431 -106737 -45375 -106693
rect -45331 -106737 -45275 -106693
rect -45231 -106737 -45175 -106693
rect -45131 -106737 -45075 -106693
rect -45031 -106737 -44975 -106693
rect -44931 -106737 -44875 -106693
rect -44831 -106737 -44775 -106693
rect -44731 -106737 -44675 -106693
rect -44631 -106737 -44575 -106693
rect -44531 -106737 -44075 -106693
rect -44031 -106737 -43975 -106693
rect -43931 -106737 -43875 -106693
rect -43831 -106737 -43775 -106693
rect -43731 -106737 -43675 -106693
rect -43631 -106737 -43575 -106693
rect -43531 -106737 -43475 -106693
rect -43431 -106737 -43375 -106693
rect -43331 -106737 -43275 -106693
rect -43231 -106737 -43175 -106693
rect -43131 -106737 -43075 -106693
rect -43031 -106737 -42975 -106693
rect -42931 -106737 -42875 -106693
rect -42831 -106737 -42775 -106693
rect -42731 -106737 -42675 -106693
rect -42631 -106737 -42575 -106693
rect -42531 -106737 -42000 -106693
rect -50768 -106793 -42000 -106737
rect -50768 -106837 -50075 -106793
rect -50031 -106837 -49975 -106793
rect -49931 -106837 -49875 -106793
rect -49831 -106837 -49775 -106793
rect -49731 -106837 -49675 -106793
rect -49631 -106837 -49575 -106793
rect -49531 -106837 -49475 -106793
rect -49431 -106837 -49375 -106793
rect -49331 -106837 -49275 -106793
rect -49231 -106837 -49175 -106793
rect -49131 -106837 -49075 -106793
rect -49031 -106837 -48975 -106793
rect -48931 -106837 -48875 -106793
rect -48831 -106837 -48775 -106793
rect -48731 -106837 -48675 -106793
rect -48631 -106837 -48575 -106793
rect -48531 -106837 -48075 -106793
rect -48031 -106837 -47975 -106793
rect -47931 -106837 -47875 -106793
rect -47831 -106837 -47775 -106793
rect -47731 -106837 -47675 -106793
rect -47631 -106837 -47575 -106793
rect -47531 -106837 -47475 -106793
rect -47431 -106837 -47375 -106793
rect -47331 -106837 -47275 -106793
rect -47231 -106837 -47175 -106793
rect -47131 -106837 -47075 -106793
rect -47031 -106837 -46975 -106793
rect -46931 -106837 -46875 -106793
rect -46831 -106837 -46775 -106793
rect -46731 -106837 -46675 -106793
rect -46631 -106837 -46575 -106793
rect -46531 -106837 -46075 -106793
rect -46031 -106837 -45975 -106793
rect -45931 -106837 -45875 -106793
rect -45831 -106837 -45775 -106793
rect -45731 -106837 -45675 -106793
rect -45631 -106837 -45575 -106793
rect -45531 -106837 -45475 -106793
rect -45431 -106837 -45375 -106793
rect -45331 -106837 -45275 -106793
rect -45231 -106837 -45175 -106793
rect -45131 -106837 -45075 -106793
rect -45031 -106837 -44975 -106793
rect -44931 -106837 -44875 -106793
rect -44831 -106837 -44775 -106793
rect -44731 -106837 -44675 -106793
rect -44631 -106837 -44575 -106793
rect -44531 -106837 -44075 -106793
rect -44031 -106837 -43975 -106793
rect -43931 -106837 -43875 -106793
rect -43831 -106837 -43775 -106793
rect -43731 -106837 -43675 -106793
rect -43631 -106837 -43575 -106793
rect -43531 -106837 -43475 -106793
rect -43431 -106837 -43375 -106793
rect -43331 -106837 -43275 -106793
rect -43231 -106837 -43175 -106793
rect -43131 -106837 -43075 -106793
rect -43031 -106837 -42975 -106793
rect -42931 -106837 -42875 -106793
rect -42831 -106837 -42775 -106793
rect -42731 -106837 -42675 -106793
rect -42631 -106837 -42575 -106793
rect -42531 -106837 -42000 -106793
rect -50768 -106893 -42000 -106837
rect -50768 -106937 -50075 -106893
rect -50031 -106937 -49975 -106893
rect -49931 -106937 -49875 -106893
rect -49831 -106937 -49775 -106893
rect -49731 -106937 -49675 -106893
rect -49631 -106937 -49575 -106893
rect -49531 -106937 -49475 -106893
rect -49431 -106937 -49375 -106893
rect -49331 -106937 -49275 -106893
rect -49231 -106937 -49175 -106893
rect -49131 -106937 -49075 -106893
rect -49031 -106937 -48975 -106893
rect -48931 -106937 -48875 -106893
rect -48831 -106937 -48775 -106893
rect -48731 -106937 -48675 -106893
rect -48631 -106937 -48575 -106893
rect -48531 -106937 -48075 -106893
rect -48031 -106937 -47975 -106893
rect -47931 -106937 -47875 -106893
rect -47831 -106937 -47775 -106893
rect -47731 -106937 -47675 -106893
rect -47631 -106937 -47575 -106893
rect -47531 -106937 -47475 -106893
rect -47431 -106937 -47375 -106893
rect -47331 -106937 -47275 -106893
rect -47231 -106937 -47175 -106893
rect -47131 -106937 -47075 -106893
rect -47031 -106937 -46975 -106893
rect -46931 -106937 -46875 -106893
rect -46831 -106937 -46775 -106893
rect -46731 -106937 -46675 -106893
rect -46631 -106937 -46575 -106893
rect -46531 -106937 -46075 -106893
rect -46031 -106937 -45975 -106893
rect -45931 -106937 -45875 -106893
rect -45831 -106937 -45775 -106893
rect -45731 -106937 -45675 -106893
rect -45631 -106937 -45575 -106893
rect -45531 -106937 -45475 -106893
rect -45431 -106937 -45375 -106893
rect -45331 -106937 -45275 -106893
rect -45231 -106937 -45175 -106893
rect -45131 -106937 -45075 -106893
rect -45031 -106937 -44975 -106893
rect -44931 -106937 -44875 -106893
rect -44831 -106937 -44775 -106893
rect -44731 -106937 -44675 -106893
rect -44631 -106937 -44575 -106893
rect -44531 -106937 -44075 -106893
rect -44031 -106937 -43975 -106893
rect -43931 -106937 -43875 -106893
rect -43831 -106937 -43775 -106893
rect -43731 -106937 -43675 -106893
rect -43631 -106937 -43575 -106893
rect -43531 -106937 -43475 -106893
rect -43431 -106937 -43375 -106893
rect -43331 -106937 -43275 -106893
rect -43231 -106937 -43175 -106893
rect -43131 -106937 -43075 -106893
rect -43031 -106937 -42975 -106893
rect -42931 -106937 -42875 -106893
rect -42831 -106937 -42775 -106893
rect -42731 -106937 -42675 -106893
rect -42631 -106937 -42575 -106893
rect -42531 -106937 -42000 -106893
rect -50768 -106993 -42000 -106937
rect -50768 -107037 -50075 -106993
rect -50031 -107037 -49975 -106993
rect -49931 -107037 -49875 -106993
rect -49831 -107037 -49775 -106993
rect -49731 -107037 -49675 -106993
rect -49631 -107037 -49575 -106993
rect -49531 -107037 -49475 -106993
rect -49431 -107037 -49375 -106993
rect -49331 -107037 -49275 -106993
rect -49231 -107037 -49175 -106993
rect -49131 -107037 -49075 -106993
rect -49031 -107037 -48975 -106993
rect -48931 -107037 -48875 -106993
rect -48831 -107037 -48775 -106993
rect -48731 -107037 -48675 -106993
rect -48631 -107037 -48575 -106993
rect -48531 -107037 -48075 -106993
rect -48031 -107037 -47975 -106993
rect -47931 -107037 -47875 -106993
rect -47831 -107037 -47775 -106993
rect -47731 -107037 -47675 -106993
rect -47631 -107037 -47575 -106993
rect -47531 -107037 -47475 -106993
rect -47431 -107037 -47375 -106993
rect -47331 -107037 -47275 -106993
rect -47231 -107037 -47175 -106993
rect -47131 -107037 -47075 -106993
rect -47031 -107037 -46975 -106993
rect -46931 -107037 -46875 -106993
rect -46831 -107037 -46775 -106993
rect -46731 -107037 -46675 -106993
rect -46631 -107037 -46575 -106993
rect -46531 -107037 -46075 -106993
rect -46031 -107037 -45975 -106993
rect -45931 -107037 -45875 -106993
rect -45831 -107037 -45775 -106993
rect -45731 -107037 -45675 -106993
rect -45631 -107037 -45575 -106993
rect -45531 -107037 -45475 -106993
rect -45431 -107037 -45375 -106993
rect -45331 -107037 -45275 -106993
rect -45231 -107037 -45175 -106993
rect -45131 -107037 -45075 -106993
rect -45031 -107037 -44975 -106993
rect -44931 -107037 -44875 -106993
rect -44831 -107037 -44775 -106993
rect -44731 -107037 -44675 -106993
rect -44631 -107037 -44575 -106993
rect -44531 -107037 -44075 -106993
rect -44031 -107037 -43975 -106993
rect -43931 -107037 -43875 -106993
rect -43831 -107037 -43775 -106993
rect -43731 -107037 -43675 -106993
rect -43631 -107037 -43575 -106993
rect -43531 -107037 -43475 -106993
rect -43431 -107037 -43375 -106993
rect -43331 -107037 -43275 -106993
rect -43231 -107037 -43175 -106993
rect -43131 -107037 -43075 -106993
rect -43031 -107037 -42975 -106993
rect -42931 -107037 -42875 -106993
rect -42831 -107037 -42775 -106993
rect -42731 -107037 -42675 -106993
rect -42631 -107037 -42575 -106993
rect -42531 -107037 -42000 -106993
rect -50768 -107093 -42000 -107037
rect -50768 -107137 -50075 -107093
rect -50031 -107137 -49975 -107093
rect -49931 -107137 -49875 -107093
rect -49831 -107137 -49775 -107093
rect -49731 -107137 -49675 -107093
rect -49631 -107137 -49575 -107093
rect -49531 -107137 -49475 -107093
rect -49431 -107137 -49375 -107093
rect -49331 -107137 -49275 -107093
rect -49231 -107137 -49175 -107093
rect -49131 -107137 -49075 -107093
rect -49031 -107137 -48975 -107093
rect -48931 -107137 -48875 -107093
rect -48831 -107137 -48775 -107093
rect -48731 -107137 -48675 -107093
rect -48631 -107137 -48575 -107093
rect -48531 -107137 -48075 -107093
rect -48031 -107137 -47975 -107093
rect -47931 -107137 -47875 -107093
rect -47831 -107137 -47775 -107093
rect -47731 -107137 -47675 -107093
rect -47631 -107137 -47575 -107093
rect -47531 -107137 -47475 -107093
rect -47431 -107137 -47375 -107093
rect -47331 -107137 -47275 -107093
rect -47231 -107137 -47175 -107093
rect -47131 -107137 -47075 -107093
rect -47031 -107137 -46975 -107093
rect -46931 -107137 -46875 -107093
rect -46831 -107137 -46775 -107093
rect -46731 -107137 -46675 -107093
rect -46631 -107137 -46575 -107093
rect -46531 -107137 -46075 -107093
rect -46031 -107137 -45975 -107093
rect -45931 -107137 -45875 -107093
rect -45831 -107137 -45775 -107093
rect -45731 -107137 -45675 -107093
rect -45631 -107137 -45575 -107093
rect -45531 -107137 -45475 -107093
rect -45431 -107137 -45375 -107093
rect -45331 -107137 -45275 -107093
rect -45231 -107137 -45175 -107093
rect -45131 -107137 -45075 -107093
rect -45031 -107137 -44975 -107093
rect -44931 -107137 -44875 -107093
rect -44831 -107137 -44775 -107093
rect -44731 -107137 -44675 -107093
rect -44631 -107137 -44575 -107093
rect -44531 -107137 -44075 -107093
rect -44031 -107137 -43975 -107093
rect -43931 -107137 -43875 -107093
rect -43831 -107137 -43775 -107093
rect -43731 -107137 -43675 -107093
rect -43631 -107137 -43575 -107093
rect -43531 -107137 -43475 -107093
rect -43431 -107137 -43375 -107093
rect -43331 -107137 -43275 -107093
rect -43231 -107137 -43175 -107093
rect -43131 -107137 -43075 -107093
rect -43031 -107137 -42975 -107093
rect -42931 -107137 -42875 -107093
rect -42831 -107137 -42775 -107093
rect -42731 -107137 -42675 -107093
rect -42631 -107137 -42575 -107093
rect -42531 -107137 -42000 -107093
rect -50768 -107193 -42000 -107137
rect -50768 -107237 -50075 -107193
rect -50031 -107237 -49975 -107193
rect -49931 -107237 -49875 -107193
rect -49831 -107237 -49775 -107193
rect -49731 -107237 -49675 -107193
rect -49631 -107237 -49575 -107193
rect -49531 -107237 -49475 -107193
rect -49431 -107237 -49375 -107193
rect -49331 -107237 -49275 -107193
rect -49231 -107237 -49175 -107193
rect -49131 -107237 -49075 -107193
rect -49031 -107237 -48975 -107193
rect -48931 -107237 -48875 -107193
rect -48831 -107237 -48775 -107193
rect -48731 -107237 -48675 -107193
rect -48631 -107237 -48575 -107193
rect -48531 -107237 -48075 -107193
rect -48031 -107237 -47975 -107193
rect -47931 -107237 -47875 -107193
rect -47831 -107237 -47775 -107193
rect -47731 -107237 -47675 -107193
rect -47631 -107237 -47575 -107193
rect -47531 -107237 -47475 -107193
rect -47431 -107237 -47375 -107193
rect -47331 -107237 -47275 -107193
rect -47231 -107237 -47175 -107193
rect -47131 -107237 -47075 -107193
rect -47031 -107237 -46975 -107193
rect -46931 -107237 -46875 -107193
rect -46831 -107237 -46775 -107193
rect -46731 -107237 -46675 -107193
rect -46631 -107237 -46575 -107193
rect -46531 -107237 -46075 -107193
rect -46031 -107237 -45975 -107193
rect -45931 -107237 -45875 -107193
rect -45831 -107237 -45775 -107193
rect -45731 -107237 -45675 -107193
rect -45631 -107237 -45575 -107193
rect -45531 -107237 -45475 -107193
rect -45431 -107237 -45375 -107193
rect -45331 -107237 -45275 -107193
rect -45231 -107237 -45175 -107193
rect -45131 -107237 -45075 -107193
rect -45031 -107237 -44975 -107193
rect -44931 -107237 -44875 -107193
rect -44831 -107237 -44775 -107193
rect -44731 -107237 -44675 -107193
rect -44631 -107237 -44575 -107193
rect -44531 -107237 -44075 -107193
rect -44031 -107237 -43975 -107193
rect -43931 -107237 -43875 -107193
rect -43831 -107237 -43775 -107193
rect -43731 -107237 -43675 -107193
rect -43631 -107237 -43575 -107193
rect -43531 -107237 -43475 -107193
rect -43431 -107237 -43375 -107193
rect -43331 -107237 -43275 -107193
rect -43231 -107237 -43175 -107193
rect -43131 -107237 -43075 -107193
rect -43031 -107237 -42975 -107193
rect -42931 -107237 -42875 -107193
rect -42831 -107237 -42775 -107193
rect -42731 -107237 -42675 -107193
rect -42631 -107237 -42575 -107193
rect -42531 -107237 -42000 -107193
rect -50768 -107293 -42000 -107237
rect -50768 -107337 -50075 -107293
rect -50031 -107337 -49975 -107293
rect -49931 -107337 -49875 -107293
rect -49831 -107337 -49775 -107293
rect -49731 -107337 -49675 -107293
rect -49631 -107337 -49575 -107293
rect -49531 -107337 -49475 -107293
rect -49431 -107337 -49375 -107293
rect -49331 -107337 -49275 -107293
rect -49231 -107337 -49175 -107293
rect -49131 -107337 -49075 -107293
rect -49031 -107337 -48975 -107293
rect -48931 -107337 -48875 -107293
rect -48831 -107337 -48775 -107293
rect -48731 -107337 -48675 -107293
rect -48631 -107337 -48575 -107293
rect -48531 -107337 -48075 -107293
rect -48031 -107337 -47975 -107293
rect -47931 -107337 -47875 -107293
rect -47831 -107337 -47775 -107293
rect -47731 -107337 -47675 -107293
rect -47631 -107337 -47575 -107293
rect -47531 -107337 -47475 -107293
rect -47431 -107337 -47375 -107293
rect -47331 -107337 -47275 -107293
rect -47231 -107337 -47175 -107293
rect -47131 -107337 -47075 -107293
rect -47031 -107337 -46975 -107293
rect -46931 -107337 -46875 -107293
rect -46831 -107337 -46775 -107293
rect -46731 -107337 -46675 -107293
rect -46631 -107337 -46575 -107293
rect -46531 -107337 -46075 -107293
rect -46031 -107337 -45975 -107293
rect -45931 -107337 -45875 -107293
rect -45831 -107337 -45775 -107293
rect -45731 -107337 -45675 -107293
rect -45631 -107337 -45575 -107293
rect -45531 -107337 -45475 -107293
rect -45431 -107337 -45375 -107293
rect -45331 -107337 -45275 -107293
rect -45231 -107337 -45175 -107293
rect -45131 -107337 -45075 -107293
rect -45031 -107337 -44975 -107293
rect -44931 -107337 -44875 -107293
rect -44831 -107337 -44775 -107293
rect -44731 -107337 -44675 -107293
rect -44631 -107337 -44575 -107293
rect -44531 -107337 -44075 -107293
rect -44031 -107337 -43975 -107293
rect -43931 -107337 -43875 -107293
rect -43831 -107337 -43775 -107293
rect -43731 -107337 -43675 -107293
rect -43631 -107337 -43575 -107293
rect -43531 -107337 -43475 -107293
rect -43431 -107337 -43375 -107293
rect -43331 -107337 -43275 -107293
rect -43231 -107337 -43175 -107293
rect -43131 -107337 -43075 -107293
rect -43031 -107337 -42975 -107293
rect -42931 -107337 -42875 -107293
rect -42831 -107337 -42775 -107293
rect -42731 -107337 -42675 -107293
rect -42631 -107337 -42575 -107293
rect -42531 -107337 -42000 -107293
rect -50768 -107393 -42000 -107337
rect -50768 -107437 -50075 -107393
rect -50031 -107437 -49975 -107393
rect -49931 -107437 -49875 -107393
rect -49831 -107437 -49775 -107393
rect -49731 -107437 -49675 -107393
rect -49631 -107437 -49575 -107393
rect -49531 -107437 -49475 -107393
rect -49431 -107437 -49375 -107393
rect -49331 -107437 -49275 -107393
rect -49231 -107437 -49175 -107393
rect -49131 -107437 -49075 -107393
rect -49031 -107437 -48975 -107393
rect -48931 -107437 -48875 -107393
rect -48831 -107437 -48775 -107393
rect -48731 -107437 -48675 -107393
rect -48631 -107437 -48575 -107393
rect -48531 -107437 -48075 -107393
rect -48031 -107437 -47975 -107393
rect -47931 -107437 -47875 -107393
rect -47831 -107437 -47775 -107393
rect -47731 -107437 -47675 -107393
rect -47631 -107437 -47575 -107393
rect -47531 -107437 -47475 -107393
rect -47431 -107437 -47375 -107393
rect -47331 -107437 -47275 -107393
rect -47231 -107437 -47175 -107393
rect -47131 -107437 -47075 -107393
rect -47031 -107437 -46975 -107393
rect -46931 -107437 -46875 -107393
rect -46831 -107437 -46775 -107393
rect -46731 -107437 -46675 -107393
rect -46631 -107437 -46575 -107393
rect -46531 -107437 -46075 -107393
rect -46031 -107437 -45975 -107393
rect -45931 -107437 -45875 -107393
rect -45831 -107437 -45775 -107393
rect -45731 -107437 -45675 -107393
rect -45631 -107437 -45575 -107393
rect -45531 -107437 -45475 -107393
rect -45431 -107437 -45375 -107393
rect -45331 -107437 -45275 -107393
rect -45231 -107437 -45175 -107393
rect -45131 -107437 -45075 -107393
rect -45031 -107437 -44975 -107393
rect -44931 -107437 -44875 -107393
rect -44831 -107437 -44775 -107393
rect -44731 -107437 -44675 -107393
rect -44631 -107437 -44575 -107393
rect -44531 -107437 -44075 -107393
rect -44031 -107437 -43975 -107393
rect -43931 -107437 -43875 -107393
rect -43831 -107437 -43775 -107393
rect -43731 -107437 -43675 -107393
rect -43631 -107437 -43575 -107393
rect -43531 -107437 -43475 -107393
rect -43431 -107437 -43375 -107393
rect -43331 -107437 -43275 -107393
rect -43231 -107437 -43175 -107393
rect -43131 -107437 -43075 -107393
rect -43031 -107437 -42975 -107393
rect -42931 -107437 -42875 -107393
rect -42831 -107437 -42775 -107393
rect -42731 -107437 -42675 -107393
rect -42631 -107437 -42575 -107393
rect -42531 -107437 -42000 -107393
rect -50768 -107493 -42000 -107437
rect -50768 -107537 -50075 -107493
rect -50031 -107537 -49975 -107493
rect -49931 -107537 -49875 -107493
rect -49831 -107537 -49775 -107493
rect -49731 -107537 -49675 -107493
rect -49631 -107537 -49575 -107493
rect -49531 -107537 -49475 -107493
rect -49431 -107537 -49375 -107493
rect -49331 -107537 -49275 -107493
rect -49231 -107537 -49175 -107493
rect -49131 -107537 -49075 -107493
rect -49031 -107537 -48975 -107493
rect -48931 -107537 -48875 -107493
rect -48831 -107537 -48775 -107493
rect -48731 -107537 -48675 -107493
rect -48631 -107537 -48575 -107493
rect -48531 -107537 -48075 -107493
rect -48031 -107537 -47975 -107493
rect -47931 -107537 -47875 -107493
rect -47831 -107537 -47775 -107493
rect -47731 -107537 -47675 -107493
rect -47631 -107537 -47575 -107493
rect -47531 -107537 -47475 -107493
rect -47431 -107537 -47375 -107493
rect -47331 -107537 -47275 -107493
rect -47231 -107537 -47175 -107493
rect -47131 -107537 -47075 -107493
rect -47031 -107537 -46975 -107493
rect -46931 -107537 -46875 -107493
rect -46831 -107537 -46775 -107493
rect -46731 -107537 -46675 -107493
rect -46631 -107537 -46575 -107493
rect -46531 -107537 -46075 -107493
rect -46031 -107537 -45975 -107493
rect -45931 -107537 -45875 -107493
rect -45831 -107537 -45775 -107493
rect -45731 -107537 -45675 -107493
rect -45631 -107537 -45575 -107493
rect -45531 -107537 -45475 -107493
rect -45431 -107537 -45375 -107493
rect -45331 -107537 -45275 -107493
rect -45231 -107537 -45175 -107493
rect -45131 -107537 -45075 -107493
rect -45031 -107537 -44975 -107493
rect -44931 -107537 -44875 -107493
rect -44831 -107537 -44775 -107493
rect -44731 -107537 -44675 -107493
rect -44631 -107537 -44575 -107493
rect -44531 -107537 -44075 -107493
rect -44031 -107537 -43975 -107493
rect -43931 -107537 -43875 -107493
rect -43831 -107537 -43775 -107493
rect -43731 -107537 -43675 -107493
rect -43631 -107537 -43575 -107493
rect -43531 -107537 -43475 -107493
rect -43431 -107537 -43375 -107493
rect -43331 -107537 -43275 -107493
rect -43231 -107537 -43175 -107493
rect -43131 -107537 -43075 -107493
rect -43031 -107537 -42975 -107493
rect -42931 -107537 -42875 -107493
rect -42831 -107537 -42775 -107493
rect -42731 -107537 -42675 -107493
rect -42631 -107537 -42575 -107493
rect -42531 -107537 -42000 -107493
rect -50768 -107593 -42000 -107537
rect -50768 -107637 -50075 -107593
rect -50031 -107637 -49975 -107593
rect -49931 -107637 -49875 -107593
rect -49831 -107637 -49775 -107593
rect -49731 -107637 -49675 -107593
rect -49631 -107637 -49575 -107593
rect -49531 -107637 -49475 -107593
rect -49431 -107637 -49375 -107593
rect -49331 -107637 -49275 -107593
rect -49231 -107637 -49175 -107593
rect -49131 -107637 -49075 -107593
rect -49031 -107637 -48975 -107593
rect -48931 -107637 -48875 -107593
rect -48831 -107637 -48775 -107593
rect -48731 -107637 -48675 -107593
rect -48631 -107637 -48575 -107593
rect -48531 -107637 -48075 -107593
rect -48031 -107637 -47975 -107593
rect -47931 -107637 -47875 -107593
rect -47831 -107637 -47775 -107593
rect -47731 -107637 -47675 -107593
rect -47631 -107637 -47575 -107593
rect -47531 -107637 -47475 -107593
rect -47431 -107637 -47375 -107593
rect -47331 -107637 -47275 -107593
rect -47231 -107637 -47175 -107593
rect -47131 -107637 -47075 -107593
rect -47031 -107637 -46975 -107593
rect -46931 -107637 -46875 -107593
rect -46831 -107637 -46775 -107593
rect -46731 -107637 -46675 -107593
rect -46631 -107637 -46575 -107593
rect -46531 -107637 -46075 -107593
rect -46031 -107637 -45975 -107593
rect -45931 -107637 -45875 -107593
rect -45831 -107637 -45775 -107593
rect -45731 -107637 -45675 -107593
rect -45631 -107637 -45575 -107593
rect -45531 -107637 -45475 -107593
rect -45431 -107637 -45375 -107593
rect -45331 -107637 -45275 -107593
rect -45231 -107637 -45175 -107593
rect -45131 -107637 -45075 -107593
rect -45031 -107637 -44975 -107593
rect -44931 -107637 -44875 -107593
rect -44831 -107637 -44775 -107593
rect -44731 -107637 -44675 -107593
rect -44631 -107637 -44575 -107593
rect -44531 -107637 -44075 -107593
rect -44031 -107637 -43975 -107593
rect -43931 -107637 -43875 -107593
rect -43831 -107637 -43775 -107593
rect -43731 -107637 -43675 -107593
rect -43631 -107637 -43575 -107593
rect -43531 -107637 -43475 -107593
rect -43431 -107637 -43375 -107593
rect -43331 -107637 -43275 -107593
rect -43231 -107637 -43175 -107593
rect -43131 -107637 -43075 -107593
rect -43031 -107637 -42975 -107593
rect -42931 -107637 -42875 -107593
rect -42831 -107637 -42775 -107593
rect -42731 -107637 -42675 -107593
rect -42631 -107637 -42575 -107593
rect -42531 -107637 -42000 -107593
rect -50768 -107693 -42000 -107637
rect -50768 -107737 -50075 -107693
rect -50031 -107737 -49975 -107693
rect -49931 -107737 -49875 -107693
rect -49831 -107737 -49775 -107693
rect -49731 -107737 -49675 -107693
rect -49631 -107737 -49575 -107693
rect -49531 -107737 -49475 -107693
rect -49431 -107737 -49375 -107693
rect -49331 -107737 -49275 -107693
rect -49231 -107737 -49175 -107693
rect -49131 -107737 -49075 -107693
rect -49031 -107737 -48975 -107693
rect -48931 -107737 -48875 -107693
rect -48831 -107737 -48775 -107693
rect -48731 -107737 -48675 -107693
rect -48631 -107737 -48575 -107693
rect -48531 -107737 -48075 -107693
rect -48031 -107737 -47975 -107693
rect -47931 -107737 -47875 -107693
rect -47831 -107737 -47775 -107693
rect -47731 -107737 -47675 -107693
rect -47631 -107737 -47575 -107693
rect -47531 -107737 -47475 -107693
rect -47431 -107737 -47375 -107693
rect -47331 -107737 -47275 -107693
rect -47231 -107737 -47175 -107693
rect -47131 -107737 -47075 -107693
rect -47031 -107737 -46975 -107693
rect -46931 -107737 -46875 -107693
rect -46831 -107737 -46775 -107693
rect -46731 -107737 -46675 -107693
rect -46631 -107737 -46575 -107693
rect -46531 -107737 -46075 -107693
rect -46031 -107737 -45975 -107693
rect -45931 -107737 -45875 -107693
rect -45831 -107737 -45775 -107693
rect -45731 -107737 -45675 -107693
rect -45631 -107737 -45575 -107693
rect -45531 -107737 -45475 -107693
rect -45431 -107737 -45375 -107693
rect -45331 -107737 -45275 -107693
rect -45231 -107737 -45175 -107693
rect -45131 -107737 -45075 -107693
rect -45031 -107737 -44975 -107693
rect -44931 -107737 -44875 -107693
rect -44831 -107737 -44775 -107693
rect -44731 -107737 -44675 -107693
rect -44631 -107737 -44575 -107693
rect -44531 -107737 -44075 -107693
rect -44031 -107737 -43975 -107693
rect -43931 -107737 -43875 -107693
rect -43831 -107737 -43775 -107693
rect -43731 -107737 -43675 -107693
rect -43631 -107737 -43575 -107693
rect -43531 -107737 -43475 -107693
rect -43431 -107737 -43375 -107693
rect -43331 -107737 -43275 -107693
rect -43231 -107737 -43175 -107693
rect -43131 -107737 -43075 -107693
rect -43031 -107737 -42975 -107693
rect -42931 -107737 -42875 -107693
rect -42831 -107737 -42775 -107693
rect -42731 -107737 -42675 -107693
rect -42631 -107737 -42575 -107693
rect -42531 -107737 -42000 -107693
rect -50768 -108598 -42000 -107737
rect -16409 -131251 -2893 -13656
rect 7194 -11056 18364 -11000
rect 7194 -11100 9195 -11056
rect 9239 -11100 9295 -11056
rect 9339 -11100 9395 -11056
rect 9439 -11100 9495 -11056
rect 9539 -11100 9595 -11056
rect 9639 -11100 9695 -11056
rect 9739 -11100 9795 -11056
rect 9839 -11100 9895 -11056
rect 9939 -11100 9995 -11056
rect 10039 -11100 10095 -11056
rect 10139 -11100 10195 -11056
rect 10239 -11100 10295 -11056
rect 10339 -11100 10395 -11056
rect 10439 -11100 10495 -11056
rect 10539 -11100 10595 -11056
rect 10639 -11100 10695 -11056
rect 10739 -11100 11195 -11056
rect 11239 -11100 11295 -11056
rect 11339 -11100 11395 -11056
rect 11439 -11100 11495 -11056
rect 11539 -11100 11595 -11056
rect 11639 -11100 11695 -11056
rect 11739 -11100 11795 -11056
rect 11839 -11100 11895 -11056
rect 11939 -11100 11995 -11056
rect 12039 -11100 12095 -11056
rect 12139 -11100 12195 -11056
rect 12239 -11100 12295 -11056
rect 12339 -11100 12395 -11056
rect 12439 -11100 12495 -11056
rect 12539 -11100 12595 -11056
rect 12639 -11100 12695 -11056
rect 12739 -11100 13195 -11056
rect 13239 -11100 13295 -11056
rect 13339 -11100 13395 -11056
rect 13439 -11100 13495 -11056
rect 13539 -11100 13595 -11056
rect 13639 -11100 13695 -11056
rect 13739 -11100 13795 -11056
rect 13839 -11100 13895 -11056
rect 13939 -11100 13995 -11056
rect 14039 -11100 14095 -11056
rect 14139 -11100 14195 -11056
rect 14239 -11100 14295 -11056
rect 14339 -11100 14395 -11056
rect 14439 -11100 14495 -11056
rect 14539 -11100 14595 -11056
rect 14639 -11100 14695 -11056
rect 14739 -11100 15195 -11056
rect 15239 -11100 15295 -11056
rect 15339 -11100 15395 -11056
rect 15439 -11100 15495 -11056
rect 15539 -11100 15595 -11056
rect 15639 -11100 15695 -11056
rect 15739 -11100 15795 -11056
rect 15839 -11100 15895 -11056
rect 15939 -11100 15995 -11056
rect 16039 -11100 16095 -11056
rect 16139 -11100 16195 -11056
rect 16239 -11100 16295 -11056
rect 16339 -11100 16395 -11056
rect 16439 -11100 16495 -11056
rect 16539 -11100 16595 -11056
rect 16639 -11100 16695 -11056
rect 16739 -11100 18364 -11056
rect 7194 -11156 18364 -11100
rect 7194 -11200 9195 -11156
rect 9239 -11200 9295 -11156
rect 9339 -11200 9395 -11156
rect 9439 -11200 9495 -11156
rect 9539 -11200 9595 -11156
rect 9639 -11200 9695 -11156
rect 9739 -11200 9795 -11156
rect 9839 -11200 9895 -11156
rect 9939 -11200 9995 -11156
rect 10039 -11200 10095 -11156
rect 10139 -11200 10195 -11156
rect 10239 -11200 10295 -11156
rect 10339 -11200 10395 -11156
rect 10439 -11200 10495 -11156
rect 10539 -11200 10595 -11156
rect 10639 -11200 10695 -11156
rect 10739 -11200 11195 -11156
rect 11239 -11200 11295 -11156
rect 11339 -11200 11395 -11156
rect 11439 -11200 11495 -11156
rect 11539 -11200 11595 -11156
rect 11639 -11200 11695 -11156
rect 11739 -11200 11795 -11156
rect 11839 -11200 11895 -11156
rect 11939 -11200 11995 -11156
rect 12039 -11200 12095 -11156
rect 12139 -11200 12195 -11156
rect 12239 -11200 12295 -11156
rect 12339 -11200 12395 -11156
rect 12439 -11200 12495 -11156
rect 12539 -11200 12595 -11156
rect 12639 -11200 12695 -11156
rect 12739 -11200 13195 -11156
rect 13239 -11200 13295 -11156
rect 13339 -11200 13395 -11156
rect 13439 -11200 13495 -11156
rect 13539 -11200 13595 -11156
rect 13639 -11200 13695 -11156
rect 13739 -11200 13795 -11156
rect 13839 -11200 13895 -11156
rect 13939 -11200 13995 -11156
rect 14039 -11200 14095 -11156
rect 14139 -11200 14195 -11156
rect 14239 -11200 14295 -11156
rect 14339 -11200 14395 -11156
rect 14439 -11200 14495 -11156
rect 14539 -11200 14595 -11156
rect 14639 -11200 14695 -11156
rect 14739 -11200 15195 -11156
rect 15239 -11200 15295 -11156
rect 15339 -11200 15395 -11156
rect 15439 -11200 15495 -11156
rect 15539 -11200 15595 -11156
rect 15639 -11200 15695 -11156
rect 15739 -11200 15795 -11156
rect 15839 -11200 15895 -11156
rect 15939 -11200 15995 -11156
rect 16039 -11200 16095 -11156
rect 16139 -11200 16195 -11156
rect 16239 -11200 16295 -11156
rect 16339 -11200 16395 -11156
rect 16439 -11200 16495 -11156
rect 16539 -11200 16595 -11156
rect 16639 -11200 16695 -11156
rect 16739 -11200 18364 -11156
rect 7194 -11256 18364 -11200
rect 7194 -11300 9195 -11256
rect 9239 -11300 9295 -11256
rect 9339 -11300 9395 -11256
rect 9439 -11300 9495 -11256
rect 9539 -11300 9595 -11256
rect 9639 -11300 9695 -11256
rect 9739 -11300 9795 -11256
rect 9839 -11300 9895 -11256
rect 9939 -11300 9995 -11256
rect 10039 -11300 10095 -11256
rect 10139 -11300 10195 -11256
rect 10239 -11300 10295 -11256
rect 10339 -11300 10395 -11256
rect 10439 -11300 10495 -11256
rect 10539 -11300 10595 -11256
rect 10639 -11300 10695 -11256
rect 10739 -11300 11195 -11256
rect 11239 -11300 11295 -11256
rect 11339 -11300 11395 -11256
rect 11439 -11300 11495 -11256
rect 11539 -11300 11595 -11256
rect 11639 -11300 11695 -11256
rect 11739 -11300 11795 -11256
rect 11839 -11300 11895 -11256
rect 11939 -11300 11995 -11256
rect 12039 -11300 12095 -11256
rect 12139 -11300 12195 -11256
rect 12239 -11300 12295 -11256
rect 12339 -11300 12395 -11256
rect 12439 -11300 12495 -11256
rect 12539 -11300 12595 -11256
rect 12639 -11300 12695 -11256
rect 12739 -11300 13195 -11256
rect 13239 -11300 13295 -11256
rect 13339 -11300 13395 -11256
rect 13439 -11300 13495 -11256
rect 13539 -11300 13595 -11256
rect 13639 -11300 13695 -11256
rect 13739 -11300 13795 -11256
rect 13839 -11300 13895 -11256
rect 13939 -11300 13995 -11256
rect 14039 -11300 14095 -11256
rect 14139 -11300 14195 -11256
rect 14239 -11300 14295 -11256
rect 14339 -11300 14395 -11256
rect 14439 -11300 14495 -11256
rect 14539 -11300 14595 -11256
rect 14639 -11300 14695 -11256
rect 14739 -11300 15195 -11256
rect 15239 -11300 15295 -11256
rect 15339 -11300 15395 -11256
rect 15439 -11300 15495 -11256
rect 15539 -11300 15595 -11256
rect 15639 -11300 15695 -11256
rect 15739 -11300 15795 -11256
rect 15839 -11300 15895 -11256
rect 15939 -11300 15995 -11256
rect 16039 -11300 16095 -11256
rect 16139 -11300 16195 -11256
rect 16239 -11300 16295 -11256
rect 16339 -11300 16395 -11256
rect 16439 -11300 16495 -11256
rect 16539 -11300 16595 -11256
rect 16639 -11300 16695 -11256
rect 16739 -11300 18364 -11256
rect 7194 -75188 18364 -11300
rect 7194 -75232 9236 -75188
rect 9280 -75232 9336 -75188
rect 9380 -75232 9436 -75188
rect 9480 -75232 9536 -75188
rect 9580 -75232 9636 -75188
rect 9680 -75232 9736 -75188
rect 9780 -75232 9836 -75188
rect 9880 -75232 9936 -75188
rect 9980 -75232 10036 -75188
rect 10080 -75232 10136 -75188
rect 10180 -75232 10236 -75188
rect 10280 -75232 10336 -75188
rect 10380 -75232 10436 -75188
rect 10480 -75232 10536 -75188
rect 10580 -75232 10636 -75188
rect 10680 -75232 10736 -75188
rect 10780 -75232 11236 -75188
rect 11280 -75232 11336 -75188
rect 11380 -75232 11436 -75188
rect 11480 -75232 11536 -75188
rect 11580 -75232 11636 -75188
rect 11680 -75232 11736 -75188
rect 11780 -75232 11836 -75188
rect 11880 -75232 11936 -75188
rect 11980 -75232 12036 -75188
rect 12080 -75232 12136 -75188
rect 12180 -75232 12236 -75188
rect 12280 -75232 12336 -75188
rect 12380 -75232 12436 -75188
rect 12480 -75232 12536 -75188
rect 12580 -75232 12636 -75188
rect 12680 -75232 12736 -75188
rect 12780 -75232 13236 -75188
rect 13280 -75232 13336 -75188
rect 13380 -75232 13436 -75188
rect 13480 -75232 13536 -75188
rect 13580 -75232 13636 -75188
rect 13680 -75232 13736 -75188
rect 13780 -75232 13836 -75188
rect 13880 -75232 13936 -75188
rect 13980 -75232 14036 -75188
rect 14080 -75232 14136 -75188
rect 14180 -75232 14236 -75188
rect 14280 -75232 14336 -75188
rect 14380 -75232 14436 -75188
rect 14480 -75232 14536 -75188
rect 14580 -75232 14636 -75188
rect 14680 -75232 14736 -75188
rect 14780 -75232 15236 -75188
rect 15280 -75232 15336 -75188
rect 15380 -75232 15436 -75188
rect 15480 -75232 15536 -75188
rect 15580 -75232 15636 -75188
rect 15680 -75232 15736 -75188
rect 15780 -75232 15836 -75188
rect 15880 -75232 15936 -75188
rect 15980 -75232 16036 -75188
rect 16080 -75232 16136 -75188
rect 16180 -75232 16236 -75188
rect 16280 -75232 16336 -75188
rect 16380 -75232 16436 -75188
rect 16480 -75232 16536 -75188
rect 16580 -75232 16636 -75188
rect 16680 -75232 16736 -75188
rect 16780 -75232 18364 -75188
rect 7194 -75288 18364 -75232
rect 7194 -75332 9236 -75288
rect 9280 -75332 9336 -75288
rect 9380 -75332 9436 -75288
rect 9480 -75332 9536 -75288
rect 9580 -75332 9636 -75288
rect 9680 -75332 9736 -75288
rect 9780 -75332 9836 -75288
rect 9880 -75332 9936 -75288
rect 9980 -75332 10036 -75288
rect 10080 -75332 10136 -75288
rect 10180 -75332 10236 -75288
rect 10280 -75332 10336 -75288
rect 10380 -75332 10436 -75288
rect 10480 -75332 10536 -75288
rect 10580 -75332 10636 -75288
rect 10680 -75332 10736 -75288
rect 10780 -75332 11236 -75288
rect 11280 -75332 11336 -75288
rect 11380 -75332 11436 -75288
rect 11480 -75332 11536 -75288
rect 11580 -75332 11636 -75288
rect 11680 -75332 11736 -75288
rect 11780 -75332 11836 -75288
rect 11880 -75332 11936 -75288
rect 11980 -75332 12036 -75288
rect 12080 -75332 12136 -75288
rect 12180 -75332 12236 -75288
rect 12280 -75332 12336 -75288
rect 12380 -75332 12436 -75288
rect 12480 -75332 12536 -75288
rect 12580 -75332 12636 -75288
rect 12680 -75332 12736 -75288
rect 12780 -75332 13236 -75288
rect 13280 -75332 13336 -75288
rect 13380 -75332 13436 -75288
rect 13480 -75332 13536 -75288
rect 13580 -75332 13636 -75288
rect 13680 -75332 13736 -75288
rect 13780 -75332 13836 -75288
rect 13880 -75332 13936 -75288
rect 13980 -75332 14036 -75288
rect 14080 -75332 14136 -75288
rect 14180 -75332 14236 -75288
rect 14280 -75332 14336 -75288
rect 14380 -75332 14436 -75288
rect 14480 -75332 14536 -75288
rect 14580 -75332 14636 -75288
rect 14680 -75332 14736 -75288
rect 14780 -75332 15236 -75288
rect 15280 -75332 15336 -75288
rect 15380 -75332 15436 -75288
rect 15480 -75332 15536 -75288
rect 15580 -75332 15636 -75288
rect 15680 -75332 15736 -75288
rect 15780 -75332 15836 -75288
rect 15880 -75332 15936 -75288
rect 15980 -75332 16036 -75288
rect 16080 -75332 16136 -75288
rect 16180 -75332 16236 -75288
rect 16280 -75332 16336 -75288
rect 16380 -75332 16436 -75288
rect 16480 -75332 16536 -75288
rect 16580 -75332 16636 -75288
rect 16680 -75332 16736 -75288
rect 16780 -75332 18364 -75288
rect 7194 -75388 18364 -75332
rect 7194 -75432 9236 -75388
rect 9280 -75432 9336 -75388
rect 9380 -75432 9436 -75388
rect 9480 -75432 9536 -75388
rect 9580 -75432 9636 -75388
rect 9680 -75432 9736 -75388
rect 9780 -75432 9836 -75388
rect 9880 -75432 9936 -75388
rect 9980 -75432 10036 -75388
rect 10080 -75432 10136 -75388
rect 10180 -75432 10236 -75388
rect 10280 -75432 10336 -75388
rect 10380 -75432 10436 -75388
rect 10480 -75432 10536 -75388
rect 10580 -75432 10636 -75388
rect 10680 -75432 10736 -75388
rect 10780 -75432 11236 -75388
rect 11280 -75432 11336 -75388
rect 11380 -75432 11436 -75388
rect 11480 -75432 11536 -75388
rect 11580 -75432 11636 -75388
rect 11680 -75432 11736 -75388
rect 11780 -75432 11836 -75388
rect 11880 -75432 11936 -75388
rect 11980 -75432 12036 -75388
rect 12080 -75432 12136 -75388
rect 12180 -75432 12236 -75388
rect 12280 -75432 12336 -75388
rect 12380 -75432 12436 -75388
rect 12480 -75432 12536 -75388
rect 12580 -75432 12636 -75388
rect 12680 -75432 12736 -75388
rect 12780 -75432 13236 -75388
rect 13280 -75432 13336 -75388
rect 13380 -75432 13436 -75388
rect 13480 -75432 13536 -75388
rect 13580 -75432 13636 -75388
rect 13680 -75432 13736 -75388
rect 13780 -75432 13836 -75388
rect 13880 -75432 13936 -75388
rect 13980 -75432 14036 -75388
rect 14080 -75432 14136 -75388
rect 14180 -75432 14236 -75388
rect 14280 -75432 14336 -75388
rect 14380 -75432 14436 -75388
rect 14480 -75432 14536 -75388
rect 14580 -75432 14636 -75388
rect 14680 -75432 14736 -75388
rect 14780 -75432 15236 -75388
rect 15280 -75432 15336 -75388
rect 15380 -75432 15436 -75388
rect 15480 -75432 15536 -75388
rect 15580 -75432 15636 -75388
rect 15680 -75432 15736 -75388
rect 15780 -75432 15836 -75388
rect 15880 -75432 15936 -75388
rect 15980 -75432 16036 -75388
rect 16080 -75432 16136 -75388
rect 16180 -75432 16236 -75388
rect 16280 -75432 16336 -75388
rect 16380 -75432 16436 -75388
rect 16480 -75432 16536 -75388
rect 16580 -75432 16636 -75388
rect 16680 -75432 16736 -75388
rect 16780 -75432 18364 -75388
rect 7194 -75488 18364 -75432
rect 7194 -75532 9236 -75488
rect 9280 -75532 9336 -75488
rect 9380 -75532 9436 -75488
rect 9480 -75532 9536 -75488
rect 9580 -75532 9636 -75488
rect 9680 -75532 9736 -75488
rect 9780 -75532 9836 -75488
rect 9880 -75532 9936 -75488
rect 9980 -75532 10036 -75488
rect 10080 -75532 10136 -75488
rect 10180 -75532 10236 -75488
rect 10280 -75532 10336 -75488
rect 10380 -75532 10436 -75488
rect 10480 -75532 10536 -75488
rect 10580 -75532 10636 -75488
rect 10680 -75532 10736 -75488
rect 10780 -75532 11236 -75488
rect 11280 -75532 11336 -75488
rect 11380 -75532 11436 -75488
rect 11480 -75532 11536 -75488
rect 11580 -75532 11636 -75488
rect 11680 -75532 11736 -75488
rect 11780 -75532 11836 -75488
rect 11880 -75532 11936 -75488
rect 11980 -75532 12036 -75488
rect 12080 -75532 12136 -75488
rect 12180 -75532 12236 -75488
rect 12280 -75532 12336 -75488
rect 12380 -75532 12436 -75488
rect 12480 -75532 12536 -75488
rect 12580 -75532 12636 -75488
rect 12680 -75532 12736 -75488
rect 12780 -75532 13236 -75488
rect 13280 -75532 13336 -75488
rect 13380 -75532 13436 -75488
rect 13480 -75532 13536 -75488
rect 13580 -75532 13636 -75488
rect 13680 -75532 13736 -75488
rect 13780 -75532 13836 -75488
rect 13880 -75532 13936 -75488
rect 13980 -75532 14036 -75488
rect 14080 -75532 14136 -75488
rect 14180 -75532 14236 -75488
rect 14280 -75532 14336 -75488
rect 14380 -75532 14436 -75488
rect 14480 -75532 14536 -75488
rect 14580 -75532 14636 -75488
rect 14680 -75532 14736 -75488
rect 14780 -75532 15236 -75488
rect 15280 -75532 15336 -75488
rect 15380 -75532 15436 -75488
rect 15480 -75532 15536 -75488
rect 15580 -75532 15636 -75488
rect 15680 -75532 15736 -75488
rect 15780 -75532 15836 -75488
rect 15880 -75532 15936 -75488
rect 15980 -75532 16036 -75488
rect 16080 -75532 16136 -75488
rect 16180 -75532 16236 -75488
rect 16280 -75532 16336 -75488
rect 16380 -75532 16436 -75488
rect 16480 -75532 16536 -75488
rect 16580 -75532 16636 -75488
rect 16680 -75532 16736 -75488
rect 16780 -75532 18364 -75488
rect 7194 -75588 18364 -75532
rect 7194 -75632 9236 -75588
rect 9280 -75632 9336 -75588
rect 9380 -75632 9436 -75588
rect 9480 -75632 9536 -75588
rect 9580 -75632 9636 -75588
rect 9680 -75632 9736 -75588
rect 9780 -75632 9836 -75588
rect 9880 -75632 9936 -75588
rect 9980 -75632 10036 -75588
rect 10080 -75632 10136 -75588
rect 10180 -75632 10236 -75588
rect 10280 -75632 10336 -75588
rect 10380 -75632 10436 -75588
rect 10480 -75632 10536 -75588
rect 10580 -75632 10636 -75588
rect 10680 -75632 10736 -75588
rect 10780 -75632 11236 -75588
rect 11280 -75632 11336 -75588
rect 11380 -75632 11436 -75588
rect 11480 -75632 11536 -75588
rect 11580 -75632 11636 -75588
rect 11680 -75632 11736 -75588
rect 11780 -75632 11836 -75588
rect 11880 -75632 11936 -75588
rect 11980 -75632 12036 -75588
rect 12080 -75632 12136 -75588
rect 12180 -75632 12236 -75588
rect 12280 -75632 12336 -75588
rect 12380 -75632 12436 -75588
rect 12480 -75632 12536 -75588
rect 12580 -75632 12636 -75588
rect 12680 -75632 12736 -75588
rect 12780 -75632 13236 -75588
rect 13280 -75632 13336 -75588
rect 13380 -75632 13436 -75588
rect 13480 -75632 13536 -75588
rect 13580 -75632 13636 -75588
rect 13680 -75632 13736 -75588
rect 13780 -75632 13836 -75588
rect 13880 -75632 13936 -75588
rect 13980 -75632 14036 -75588
rect 14080 -75632 14136 -75588
rect 14180 -75632 14236 -75588
rect 14280 -75632 14336 -75588
rect 14380 -75632 14436 -75588
rect 14480 -75632 14536 -75588
rect 14580 -75632 14636 -75588
rect 14680 -75632 14736 -75588
rect 14780 -75632 15236 -75588
rect 15280 -75632 15336 -75588
rect 15380 -75632 15436 -75588
rect 15480 -75632 15536 -75588
rect 15580 -75632 15636 -75588
rect 15680 -75632 15736 -75588
rect 15780 -75632 15836 -75588
rect 15880 -75632 15936 -75588
rect 15980 -75632 16036 -75588
rect 16080 -75632 16136 -75588
rect 16180 -75632 16236 -75588
rect 16280 -75632 16336 -75588
rect 16380 -75632 16436 -75588
rect 16480 -75632 16536 -75588
rect 16580 -75632 16636 -75588
rect 16680 -75632 16736 -75588
rect 16780 -75632 18364 -75588
rect 7194 -75688 18364 -75632
rect 7194 -75732 9236 -75688
rect 9280 -75732 9336 -75688
rect 9380 -75732 9436 -75688
rect 9480 -75732 9536 -75688
rect 9580 -75732 9636 -75688
rect 9680 -75732 9736 -75688
rect 9780 -75732 9836 -75688
rect 9880 -75732 9936 -75688
rect 9980 -75732 10036 -75688
rect 10080 -75732 10136 -75688
rect 10180 -75732 10236 -75688
rect 10280 -75732 10336 -75688
rect 10380 -75732 10436 -75688
rect 10480 -75732 10536 -75688
rect 10580 -75732 10636 -75688
rect 10680 -75732 10736 -75688
rect 10780 -75732 11236 -75688
rect 11280 -75732 11336 -75688
rect 11380 -75732 11436 -75688
rect 11480 -75732 11536 -75688
rect 11580 -75732 11636 -75688
rect 11680 -75732 11736 -75688
rect 11780 -75732 11836 -75688
rect 11880 -75732 11936 -75688
rect 11980 -75732 12036 -75688
rect 12080 -75732 12136 -75688
rect 12180 -75732 12236 -75688
rect 12280 -75732 12336 -75688
rect 12380 -75732 12436 -75688
rect 12480 -75732 12536 -75688
rect 12580 -75732 12636 -75688
rect 12680 -75732 12736 -75688
rect 12780 -75732 13236 -75688
rect 13280 -75732 13336 -75688
rect 13380 -75732 13436 -75688
rect 13480 -75732 13536 -75688
rect 13580 -75732 13636 -75688
rect 13680 -75732 13736 -75688
rect 13780 -75732 13836 -75688
rect 13880 -75732 13936 -75688
rect 13980 -75732 14036 -75688
rect 14080 -75732 14136 -75688
rect 14180 -75732 14236 -75688
rect 14280 -75732 14336 -75688
rect 14380 -75732 14436 -75688
rect 14480 -75732 14536 -75688
rect 14580 -75732 14636 -75688
rect 14680 -75732 14736 -75688
rect 14780 -75732 15236 -75688
rect 15280 -75732 15336 -75688
rect 15380 -75732 15436 -75688
rect 15480 -75732 15536 -75688
rect 15580 -75732 15636 -75688
rect 15680 -75732 15736 -75688
rect 15780 -75732 15836 -75688
rect 15880 -75732 15936 -75688
rect 15980 -75732 16036 -75688
rect 16080 -75732 16136 -75688
rect 16180 -75732 16236 -75688
rect 16280 -75732 16336 -75688
rect 16380 -75732 16436 -75688
rect 16480 -75732 16536 -75688
rect 16580 -75732 16636 -75688
rect 16680 -75732 16736 -75688
rect 16780 -75732 18364 -75688
rect 7194 -75788 18364 -75732
rect 7194 -75832 9236 -75788
rect 9280 -75832 9336 -75788
rect 9380 -75832 9436 -75788
rect 9480 -75832 9536 -75788
rect 9580 -75832 9636 -75788
rect 9680 -75832 9736 -75788
rect 9780 -75832 9836 -75788
rect 9880 -75832 9936 -75788
rect 9980 -75832 10036 -75788
rect 10080 -75832 10136 -75788
rect 10180 -75832 10236 -75788
rect 10280 -75832 10336 -75788
rect 10380 -75832 10436 -75788
rect 10480 -75832 10536 -75788
rect 10580 -75832 10636 -75788
rect 10680 -75832 10736 -75788
rect 10780 -75832 11236 -75788
rect 11280 -75832 11336 -75788
rect 11380 -75832 11436 -75788
rect 11480 -75832 11536 -75788
rect 11580 -75832 11636 -75788
rect 11680 -75832 11736 -75788
rect 11780 -75832 11836 -75788
rect 11880 -75832 11936 -75788
rect 11980 -75832 12036 -75788
rect 12080 -75832 12136 -75788
rect 12180 -75832 12236 -75788
rect 12280 -75832 12336 -75788
rect 12380 -75832 12436 -75788
rect 12480 -75832 12536 -75788
rect 12580 -75832 12636 -75788
rect 12680 -75832 12736 -75788
rect 12780 -75832 13236 -75788
rect 13280 -75832 13336 -75788
rect 13380 -75832 13436 -75788
rect 13480 -75832 13536 -75788
rect 13580 -75832 13636 -75788
rect 13680 -75832 13736 -75788
rect 13780 -75832 13836 -75788
rect 13880 -75832 13936 -75788
rect 13980 -75832 14036 -75788
rect 14080 -75832 14136 -75788
rect 14180 -75832 14236 -75788
rect 14280 -75832 14336 -75788
rect 14380 -75832 14436 -75788
rect 14480 -75832 14536 -75788
rect 14580 -75832 14636 -75788
rect 14680 -75832 14736 -75788
rect 14780 -75832 15236 -75788
rect 15280 -75832 15336 -75788
rect 15380 -75832 15436 -75788
rect 15480 -75832 15536 -75788
rect 15580 -75832 15636 -75788
rect 15680 -75832 15736 -75788
rect 15780 -75832 15836 -75788
rect 15880 -75832 15936 -75788
rect 15980 -75832 16036 -75788
rect 16080 -75832 16136 -75788
rect 16180 -75832 16236 -75788
rect 16280 -75832 16336 -75788
rect 16380 -75832 16436 -75788
rect 16480 -75832 16536 -75788
rect 16580 -75832 16636 -75788
rect 16680 -75832 16736 -75788
rect 16780 -75832 18364 -75788
rect 7194 -75888 18364 -75832
rect 7194 -75932 9236 -75888
rect 9280 -75932 9336 -75888
rect 9380 -75932 9436 -75888
rect 9480 -75932 9536 -75888
rect 9580 -75932 9636 -75888
rect 9680 -75932 9736 -75888
rect 9780 -75932 9836 -75888
rect 9880 -75932 9936 -75888
rect 9980 -75932 10036 -75888
rect 10080 -75932 10136 -75888
rect 10180 -75932 10236 -75888
rect 10280 -75932 10336 -75888
rect 10380 -75932 10436 -75888
rect 10480 -75932 10536 -75888
rect 10580 -75932 10636 -75888
rect 10680 -75932 10736 -75888
rect 10780 -75932 11236 -75888
rect 11280 -75932 11336 -75888
rect 11380 -75932 11436 -75888
rect 11480 -75932 11536 -75888
rect 11580 -75932 11636 -75888
rect 11680 -75932 11736 -75888
rect 11780 -75932 11836 -75888
rect 11880 -75932 11936 -75888
rect 11980 -75932 12036 -75888
rect 12080 -75932 12136 -75888
rect 12180 -75932 12236 -75888
rect 12280 -75932 12336 -75888
rect 12380 -75932 12436 -75888
rect 12480 -75932 12536 -75888
rect 12580 -75932 12636 -75888
rect 12680 -75932 12736 -75888
rect 12780 -75932 13236 -75888
rect 13280 -75932 13336 -75888
rect 13380 -75932 13436 -75888
rect 13480 -75932 13536 -75888
rect 13580 -75932 13636 -75888
rect 13680 -75932 13736 -75888
rect 13780 -75932 13836 -75888
rect 13880 -75932 13936 -75888
rect 13980 -75932 14036 -75888
rect 14080 -75932 14136 -75888
rect 14180 -75932 14236 -75888
rect 14280 -75932 14336 -75888
rect 14380 -75932 14436 -75888
rect 14480 -75932 14536 -75888
rect 14580 -75932 14636 -75888
rect 14680 -75932 14736 -75888
rect 14780 -75932 15236 -75888
rect 15280 -75932 15336 -75888
rect 15380 -75932 15436 -75888
rect 15480 -75932 15536 -75888
rect 15580 -75932 15636 -75888
rect 15680 -75932 15736 -75888
rect 15780 -75932 15836 -75888
rect 15880 -75932 15936 -75888
rect 15980 -75932 16036 -75888
rect 16080 -75932 16136 -75888
rect 16180 -75932 16236 -75888
rect 16280 -75932 16336 -75888
rect 16380 -75932 16436 -75888
rect 16480 -75932 16536 -75888
rect 16580 -75932 16636 -75888
rect 16680 -75932 16736 -75888
rect 16780 -75932 18364 -75888
rect 7194 -75988 18364 -75932
rect 7194 -76032 9236 -75988
rect 9280 -76032 9336 -75988
rect 9380 -76032 9436 -75988
rect 9480 -76032 9536 -75988
rect 9580 -76032 9636 -75988
rect 9680 -76032 9736 -75988
rect 9780 -76032 9836 -75988
rect 9880 -76032 9936 -75988
rect 9980 -76032 10036 -75988
rect 10080 -76032 10136 -75988
rect 10180 -76032 10236 -75988
rect 10280 -76032 10336 -75988
rect 10380 -76032 10436 -75988
rect 10480 -76032 10536 -75988
rect 10580 -76032 10636 -75988
rect 10680 -76032 10736 -75988
rect 10780 -76032 11236 -75988
rect 11280 -76032 11336 -75988
rect 11380 -76032 11436 -75988
rect 11480 -76032 11536 -75988
rect 11580 -76032 11636 -75988
rect 11680 -76032 11736 -75988
rect 11780 -76032 11836 -75988
rect 11880 -76032 11936 -75988
rect 11980 -76032 12036 -75988
rect 12080 -76032 12136 -75988
rect 12180 -76032 12236 -75988
rect 12280 -76032 12336 -75988
rect 12380 -76032 12436 -75988
rect 12480 -76032 12536 -75988
rect 12580 -76032 12636 -75988
rect 12680 -76032 12736 -75988
rect 12780 -76032 13236 -75988
rect 13280 -76032 13336 -75988
rect 13380 -76032 13436 -75988
rect 13480 -76032 13536 -75988
rect 13580 -76032 13636 -75988
rect 13680 -76032 13736 -75988
rect 13780 -76032 13836 -75988
rect 13880 -76032 13936 -75988
rect 13980 -76032 14036 -75988
rect 14080 -76032 14136 -75988
rect 14180 -76032 14236 -75988
rect 14280 -76032 14336 -75988
rect 14380 -76032 14436 -75988
rect 14480 -76032 14536 -75988
rect 14580 -76032 14636 -75988
rect 14680 -76032 14736 -75988
rect 14780 -76032 15236 -75988
rect 15280 -76032 15336 -75988
rect 15380 -76032 15436 -75988
rect 15480 -76032 15536 -75988
rect 15580 -76032 15636 -75988
rect 15680 -76032 15736 -75988
rect 15780 -76032 15836 -75988
rect 15880 -76032 15936 -75988
rect 15980 -76032 16036 -75988
rect 16080 -76032 16136 -75988
rect 16180 -76032 16236 -75988
rect 16280 -76032 16336 -75988
rect 16380 -76032 16436 -75988
rect 16480 -76032 16536 -75988
rect 16580 -76032 16636 -75988
rect 16680 -76032 16736 -75988
rect 16780 -76032 18364 -75988
rect 7194 -76088 18364 -76032
rect 7194 -76132 9236 -76088
rect 9280 -76132 9336 -76088
rect 9380 -76132 9436 -76088
rect 9480 -76132 9536 -76088
rect 9580 -76132 9636 -76088
rect 9680 -76132 9736 -76088
rect 9780 -76132 9836 -76088
rect 9880 -76132 9936 -76088
rect 9980 -76132 10036 -76088
rect 10080 -76132 10136 -76088
rect 10180 -76132 10236 -76088
rect 10280 -76132 10336 -76088
rect 10380 -76132 10436 -76088
rect 10480 -76132 10536 -76088
rect 10580 -76132 10636 -76088
rect 10680 -76132 10736 -76088
rect 10780 -76132 11236 -76088
rect 11280 -76132 11336 -76088
rect 11380 -76132 11436 -76088
rect 11480 -76132 11536 -76088
rect 11580 -76132 11636 -76088
rect 11680 -76132 11736 -76088
rect 11780 -76132 11836 -76088
rect 11880 -76132 11936 -76088
rect 11980 -76132 12036 -76088
rect 12080 -76132 12136 -76088
rect 12180 -76132 12236 -76088
rect 12280 -76132 12336 -76088
rect 12380 -76132 12436 -76088
rect 12480 -76132 12536 -76088
rect 12580 -76132 12636 -76088
rect 12680 -76132 12736 -76088
rect 12780 -76132 13236 -76088
rect 13280 -76132 13336 -76088
rect 13380 -76132 13436 -76088
rect 13480 -76132 13536 -76088
rect 13580 -76132 13636 -76088
rect 13680 -76132 13736 -76088
rect 13780 -76132 13836 -76088
rect 13880 -76132 13936 -76088
rect 13980 -76132 14036 -76088
rect 14080 -76132 14136 -76088
rect 14180 -76132 14236 -76088
rect 14280 -76132 14336 -76088
rect 14380 -76132 14436 -76088
rect 14480 -76132 14536 -76088
rect 14580 -76132 14636 -76088
rect 14680 -76132 14736 -76088
rect 14780 -76132 15236 -76088
rect 15280 -76132 15336 -76088
rect 15380 -76132 15436 -76088
rect 15480 -76132 15536 -76088
rect 15580 -76132 15636 -76088
rect 15680 -76132 15736 -76088
rect 15780 -76132 15836 -76088
rect 15880 -76132 15936 -76088
rect 15980 -76132 16036 -76088
rect 16080 -76132 16136 -76088
rect 16180 -76132 16236 -76088
rect 16280 -76132 16336 -76088
rect 16380 -76132 16436 -76088
rect 16480 -76132 16536 -76088
rect 16580 -76132 16636 -76088
rect 16680 -76132 16736 -76088
rect 16780 -76132 18364 -76088
rect 7194 -76188 18364 -76132
rect 7194 -76232 9236 -76188
rect 9280 -76232 9336 -76188
rect 9380 -76232 9436 -76188
rect 9480 -76232 9536 -76188
rect 9580 -76232 9636 -76188
rect 9680 -76232 9736 -76188
rect 9780 -76232 9836 -76188
rect 9880 -76232 9936 -76188
rect 9980 -76232 10036 -76188
rect 10080 -76232 10136 -76188
rect 10180 -76232 10236 -76188
rect 10280 -76232 10336 -76188
rect 10380 -76232 10436 -76188
rect 10480 -76232 10536 -76188
rect 10580 -76232 10636 -76188
rect 10680 -76232 10736 -76188
rect 10780 -76232 11236 -76188
rect 11280 -76232 11336 -76188
rect 11380 -76232 11436 -76188
rect 11480 -76232 11536 -76188
rect 11580 -76232 11636 -76188
rect 11680 -76232 11736 -76188
rect 11780 -76232 11836 -76188
rect 11880 -76232 11936 -76188
rect 11980 -76232 12036 -76188
rect 12080 -76232 12136 -76188
rect 12180 -76232 12236 -76188
rect 12280 -76232 12336 -76188
rect 12380 -76232 12436 -76188
rect 12480 -76232 12536 -76188
rect 12580 -76232 12636 -76188
rect 12680 -76232 12736 -76188
rect 12780 -76232 13236 -76188
rect 13280 -76232 13336 -76188
rect 13380 -76232 13436 -76188
rect 13480 -76232 13536 -76188
rect 13580 -76232 13636 -76188
rect 13680 -76232 13736 -76188
rect 13780 -76232 13836 -76188
rect 13880 -76232 13936 -76188
rect 13980 -76232 14036 -76188
rect 14080 -76232 14136 -76188
rect 14180 -76232 14236 -76188
rect 14280 -76232 14336 -76188
rect 14380 -76232 14436 -76188
rect 14480 -76232 14536 -76188
rect 14580 -76232 14636 -76188
rect 14680 -76232 14736 -76188
rect 14780 -76232 15236 -76188
rect 15280 -76232 15336 -76188
rect 15380 -76232 15436 -76188
rect 15480 -76232 15536 -76188
rect 15580 -76232 15636 -76188
rect 15680 -76232 15736 -76188
rect 15780 -76232 15836 -76188
rect 15880 -76232 15936 -76188
rect 15980 -76232 16036 -76188
rect 16080 -76232 16136 -76188
rect 16180 -76232 16236 -76188
rect 16280 -76232 16336 -76188
rect 16380 -76232 16436 -76188
rect 16480 -76232 16536 -76188
rect 16580 -76232 16636 -76188
rect 16680 -76232 16736 -76188
rect 16780 -76232 18364 -76188
rect 7194 -76288 18364 -76232
rect 7194 -76332 9236 -76288
rect 9280 -76332 9336 -76288
rect 9380 -76332 9436 -76288
rect 9480 -76332 9536 -76288
rect 9580 -76332 9636 -76288
rect 9680 -76332 9736 -76288
rect 9780 -76332 9836 -76288
rect 9880 -76332 9936 -76288
rect 9980 -76332 10036 -76288
rect 10080 -76332 10136 -76288
rect 10180 -76332 10236 -76288
rect 10280 -76332 10336 -76288
rect 10380 -76332 10436 -76288
rect 10480 -76332 10536 -76288
rect 10580 -76332 10636 -76288
rect 10680 -76332 10736 -76288
rect 10780 -76332 11236 -76288
rect 11280 -76332 11336 -76288
rect 11380 -76332 11436 -76288
rect 11480 -76332 11536 -76288
rect 11580 -76332 11636 -76288
rect 11680 -76332 11736 -76288
rect 11780 -76332 11836 -76288
rect 11880 -76332 11936 -76288
rect 11980 -76332 12036 -76288
rect 12080 -76332 12136 -76288
rect 12180 -76332 12236 -76288
rect 12280 -76332 12336 -76288
rect 12380 -76332 12436 -76288
rect 12480 -76332 12536 -76288
rect 12580 -76332 12636 -76288
rect 12680 -76332 12736 -76288
rect 12780 -76332 13236 -76288
rect 13280 -76332 13336 -76288
rect 13380 -76332 13436 -76288
rect 13480 -76332 13536 -76288
rect 13580 -76332 13636 -76288
rect 13680 -76332 13736 -76288
rect 13780 -76332 13836 -76288
rect 13880 -76332 13936 -76288
rect 13980 -76332 14036 -76288
rect 14080 -76332 14136 -76288
rect 14180 -76332 14236 -76288
rect 14280 -76332 14336 -76288
rect 14380 -76332 14436 -76288
rect 14480 -76332 14536 -76288
rect 14580 -76332 14636 -76288
rect 14680 -76332 14736 -76288
rect 14780 -76332 15236 -76288
rect 15280 -76332 15336 -76288
rect 15380 -76332 15436 -76288
rect 15480 -76332 15536 -76288
rect 15580 -76332 15636 -76288
rect 15680 -76332 15736 -76288
rect 15780 -76332 15836 -76288
rect 15880 -76332 15936 -76288
rect 15980 -76332 16036 -76288
rect 16080 -76332 16136 -76288
rect 16180 -76332 16236 -76288
rect 16280 -76332 16336 -76288
rect 16380 -76332 16436 -76288
rect 16480 -76332 16536 -76288
rect 16580 -76332 16636 -76288
rect 16680 -76332 16736 -76288
rect 16780 -76332 18364 -76288
rect 7194 -76388 18364 -76332
rect 7194 -76432 9236 -76388
rect 9280 -76432 9336 -76388
rect 9380 -76432 9436 -76388
rect 9480 -76432 9536 -76388
rect 9580 -76432 9636 -76388
rect 9680 -76432 9736 -76388
rect 9780 -76432 9836 -76388
rect 9880 -76432 9936 -76388
rect 9980 -76432 10036 -76388
rect 10080 -76432 10136 -76388
rect 10180 -76432 10236 -76388
rect 10280 -76432 10336 -76388
rect 10380 -76432 10436 -76388
rect 10480 -76432 10536 -76388
rect 10580 -76432 10636 -76388
rect 10680 -76432 10736 -76388
rect 10780 -76432 11236 -76388
rect 11280 -76432 11336 -76388
rect 11380 -76432 11436 -76388
rect 11480 -76432 11536 -76388
rect 11580 -76432 11636 -76388
rect 11680 -76432 11736 -76388
rect 11780 -76432 11836 -76388
rect 11880 -76432 11936 -76388
rect 11980 -76432 12036 -76388
rect 12080 -76432 12136 -76388
rect 12180 -76432 12236 -76388
rect 12280 -76432 12336 -76388
rect 12380 -76432 12436 -76388
rect 12480 -76432 12536 -76388
rect 12580 -76432 12636 -76388
rect 12680 -76432 12736 -76388
rect 12780 -76432 13236 -76388
rect 13280 -76432 13336 -76388
rect 13380 -76432 13436 -76388
rect 13480 -76432 13536 -76388
rect 13580 -76432 13636 -76388
rect 13680 -76432 13736 -76388
rect 13780 -76432 13836 -76388
rect 13880 -76432 13936 -76388
rect 13980 -76432 14036 -76388
rect 14080 -76432 14136 -76388
rect 14180 -76432 14236 -76388
rect 14280 -76432 14336 -76388
rect 14380 -76432 14436 -76388
rect 14480 -76432 14536 -76388
rect 14580 -76432 14636 -76388
rect 14680 -76432 14736 -76388
rect 14780 -76432 15236 -76388
rect 15280 -76432 15336 -76388
rect 15380 -76432 15436 -76388
rect 15480 -76432 15536 -76388
rect 15580 -76432 15636 -76388
rect 15680 -76432 15736 -76388
rect 15780 -76432 15836 -76388
rect 15880 -76432 15936 -76388
rect 15980 -76432 16036 -76388
rect 16080 -76432 16136 -76388
rect 16180 -76432 16236 -76388
rect 16280 -76432 16336 -76388
rect 16380 -76432 16436 -76388
rect 16480 -76432 16536 -76388
rect 16580 -76432 16636 -76388
rect 16680 -76432 16736 -76388
rect 16780 -76432 18364 -76388
rect 7194 -76488 18364 -76432
rect 7194 -76532 9236 -76488
rect 9280 -76532 9336 -76488
rect 9380 -76532 9436 -76488
rect 9480 -76532 9536 -76488
rect 9580 -76532 9636 -76488
rect 9680 -76532 9736 -76488
rect 9780 -76532 9836 -76488
rect 9880 -76532 9936 -76488
rect 9980 -76532 10036 -76488
rect 10080 -76532 10136 -76488
rect 10180 -76532 10236 -76488
rect 10280 -76532 10336 -76488
rect 10380 -76532 10436 -76488
rect 10480 -76532 10536 -76488
rect 10580 -76532 10636 -76488
rect 10680 -76532 10736 -76488
rect 10780 -76532 11236 -76488
rect 11280 -76532 11336 -76488
rect 11380 -76532 11436 -76488
rect 11480 -76532 11536 -76488
rect 11580 -76532 11636 -76488
rect 11680 -76532 11736 -76488
rect 11780 -76532 11836 -76488
rect 11880 -76532 11936 -76488
rect 11980 -76532 12036 -76488
rect 12080 -76532 12136 -76488
rect 12180 -76532 12236 -76488
rect 12280 -76532 12336 -76488
rect 12380 -76532 12436 -76488
rect 12480 -76532 12536 -76488
rect 12580 -76532 12636 -76488
rect 12680 -76532 12736 -76488
rect 12780 -76532 13236 -76488
rect 13280 -76532 13336 -76488
rect 13380 -76532 13436 -76488
rect 13480 -76532 13536 -76488
rect 13580 -76532 13636 -76488
rect 13680 -76532 13736 -76488
rect 13780 -76532 13836 -76488
rect 13880 -76532 13936 -76488
rect 13980 -76532 14036 -76488
rect 14080 -76532 14136 -76488
rect 14180 -76532 14236 -76488
rect 14280 -76532 14336 -76488
rect 14380 -76532 14436 -76488
rect 14480 -76532 14536 -76488
rect 14580 -76532 14636 -76488
rect 14680 -76532 14736 -76488
rect 14780 -76532 15236 -76488
rect 15280 -76532 15336 -76488
rect 15380 -76532 15436 -76488
rect 15480 -76532 15536 -76488
rect 15580 -76532 15636 -76488
rect 15680 -76532 15736 -76488
rect 15780 -76532 15836 -76488
rect 15880 -76532 15936 -76488
rect 15980 -76532 16036 -76488
rect 16080 -76532 16136 -76488
rect 16180 -76532 16236 -76488
rect 16280 -76532 16336 -76488
rect 16380 -76532 16436 -76488
rect 16480 -76532 16536 -76488
rect 16580 -76532 16636 -76488
rect 16680 -76532 16736 -76488
rect 16780 -76532 18364 -76488
rect 7194 -76588 18364 -76532
rect 7194 -76632 9236 -76588
rect 9280 -76632 9336 -76588
rect 9380 -76632 9436 -76588
rect 9480 -76632 9536 -76588
rect 9580 -76632 9636 -76588
rect 9680 -76632 9736 -76588
rect 9780 -76632 9836 -76588
rect 9880 -76632 9936 -76588
rect 9980 -76632 10036 -76588
rect 10080 -76632 10136 -76588
rect 10180 -76632 10236 -76588
rect 10280 -76632 10336 -76588
rect 10380 -76632 10436 -76588
rect 10480 -76632 10536 -76588
rect 10580 -76632 10636 -76588
rect 10680 -76632 10736 -76588
rect 10780 -76632 11236 -76588
rect 11280 -76632 11336 -76588
rect 11380 -76632 11436 -76588
rect 11480 -76632 11536 -76588
rect 11580 -76632 11636 -76588
rect 11680 -76632 11736 -76588
rect 11780 -76632 11836 -76588
rect 11880 -76632 11936 -76588
rect 11980 -76632 12036 -76588
rect 12080 -76632 12136 -76588
rect 12180 -76632 12236 -76588
rect 12280 -76632 12336 -76588
rect 12380 -76632 12436 -76588
rect 12480 -76632 12536 -76588
rect 12580 -76632 12636 -76588
rect 12680 -76632 12736 -76588
rect 12780 -76632 13236 -76588
rect 13280 -76632 13336 -76588
rect 13380 -76632 13436 -76588
rect 13480 -76632 13536 -76588
rect 13580 -76632 13636 -76588
rect 13680 -76632 13736 -76588
rect 13780 -76632 13836 -76588
rect 13880 -76632 13936 -76588
rect 13980 -76632 14036 -76588
rect 14080 -76632 14136 -76588
rect 14180 -76632 14236 -76588
rect 14280 -76632 14336 -76588
rect 14380 -76632 14436 -76588
rect 14480 -76632 14536 -76588
rect 14580 -76632 14636 -76588
rect 14680 -76632 14736 -76588
rect 14780 -76632 15236 -76588
rect 15280 -76632 15336 -76588
rect 15380 -76632 15436 -76588
rect 15480 -76632 15536 -76588
rect 15580 -76632 15636 -76588
rect 15680 -76632 15736 -76588
rect 15780 -76632 15836 -76588
rect 15880 -76632 15936 -76588
rect 15980 -76632 16036 -76588
rect 16080 -76632 16136 -76588
rect 16180 -76632 16236 -76588
rect 16280 -76632 16336 -76588
rect 16380 -76632 16436 -76588
rect 16480 -76632 16536 -76588
rect 16580 -76632 16636 -76588
rect 16680 -76632 16736 -76588
rect 16780 -76632 18364 -76588
rect 7194 -76688 18364 -76632
rect 7194 -76732 9236 -76688
rect 9280 -76732 9336 -76688
rect 9380 -76732 9436 -76688
rect 9480 -76732 9536 -76688
rect 9580 -76732 9636 -76688
rect 9680 -76732 9736 -76688
rect 9780 -76732 9836 -76688
rect 9880 -76732 9936 -76688
rect 9980 -76732 10036 -76688
rect 10080 -76732 10136 -76688
rect 10180 -76732 10236 -76688
rect 10280 -76732 10336 -76688
rect 10380 -76732 10436 -76688
rect 10480 -76732 10536 -76688
rect 10580 -76732 10636 -76688
rect 10680 -76732 10736 -76688
rect 10780 -76732 11236 -76688
rect 11280 -76732 11336 -76688
rect 11380 -76732 11436 -76688
rect 11480 -76732 11536 -76688
rect 11580 -76732 11636 -76688
rect 11680 -76732 11736 -76688
rect 11780 -76732 11836 -76688
rect 11880 -76732 11936 -76688
rect 11980 -76732 12036 -76688
rect 12080 -76732 12136 -76688
rect 12180 -76732 12236 -76688
rect 12280 -76732 12336 -76688
rect 12380 -76732 12436 -76688
rect 12480 -76732 12536 -76688
rect 12580 -76732 12636 -76688
rect 12680 -76732 12736 -76688
rect 12780 -76732 13236 -76688
rect 13280 -76732 13336 -76688
rect 13380 -76732 13436 -76688
rect 13480 -76732 13536 -76688
rect 13580 -76732 13636 -76688
rect 13680 -76732 13736 -76688
rect 13780 -76732 13836 -76688
rect 13880 -76732 13936 -76688
rect 13980 -76732 14036 -76688
rect 14080 -76732 14136 -76688
rect 14180 -76732 14236 -76688
rect 14280 -76732 14336 -76688
rect 14380 -76732 14436 -76688
rect 14480 -76732 14536 -76688
rect 14580 -76732 14636 -76688
rect 14680 -76732 14736 -76688
rect 14780 -76732 15236 -76688
rect 15280 -76732 15336 -76688
rect 15380 -76732 15436 -76688
rect 15480 -76732 15536 -76688
rect 15580 -76732 15636 -76688
rect 15680 -76732 15736 -76688
rect 15780 -76732 15836 -76688
rect 15880 -76732 15936 -76688
rect 15980 -76732 16036 -76688
rect 16080 -76732 16136 -76688
rect 16180 -76732 16236 -76688
rect 16280 -76732 16336 -76688
rect 16380 -76732 16436 -76688
rect 16480 -76732 16536 -76688
rect 16580 -76732 16636 -76688
rect 16680 -76732 16736 -76688
rect 16780 -76732 18364 -76688
rect 7194 -77475 18364 -76732
rect 34207 -9638 47953 -7485
rect 34207 -9682 37223 -9638
rect 37267 -9682 37323 -9638
rect 37367 -9682 37423 -9638
rect 37467 -9682 37523 -9638
rect 37567 -9682 37623 -9638
rect 37667 -9682 37723 -9638
rect 37767 -9682 37823 -9638
rect 37867 -9682 37923 -9638
rect 37967 -9682 38023 -9638
rect 38067 -9682 38123 -9638
rect 38167 -9682 38223 -9638
rect 38267 -9682 38323 -9638
rect 38367 -9682 38423 -9638
rect 38467 -9682 38523 -9638
rect 38567 -9682 38623 -9638
rect 38667 -9682 38723 -9638
rect 38767 -9682 39223 -9638
rect 39267 -9682 39323 -9638
rect 39367 -9682 39423 -9638
rect 39467 -9682 39523 -9638
rect 39567 -9682 39623 -9638
rect 39667 -9682 39723 -9638
rect 39767 -9682 39823 -9638
rect 39867 -9682 39923 -9638
rect 39967 -9682 40023 -9638
rect 40067 -9682 40123 -9638
rect 40167 -9682 40223 -9638
rect 40267 -9682 40323 -9638
rect 40367 -9682 40423 -9638
rect 40467 -9682 40523 -9638
rect 40567 -9682 40623 -9638
rect 40667 -9682 40723 -9638
rect 40767 -9682 41223 -9638
rect 41267 -9682 41323 -9638
rect 41367 -9682 41423 -9638
rect 41467 -9682 41523 -9638
rect 41567 -9682 41623 -9638
rect 41667 -9682 41723 -9638
rect 41767 -9682 41823 -9638
rect 41867 -9682 41923 -9638
rect 41967 -9682 42023 -9638
rect 42067 -9682 42123 -9638
rect 42167 -9682 42223 -9638
rect 42267 -9682 42323 -9638
rect 42367 -9682 42423 -9638
rect 42467 -9682 42523 -9638
rect 42567 -9682 42623 -9638
rect 42667 -9682 42723 -9638
rect 42767 -9682 43223 -9638
rect 43267 -9682 43323 -9638
rect 43367 -9682 43423 -9638
rect 43467 -9682 43523 -9638
rect 43567 -9682 43623 -9638
rect 43667 -9682 43723 -9638
rect 43767 -9682 43823 -9638
rect 43867 -9682 43923 -9638
rect 43967 -9682 44023 -9638
rect 44067 -9682 44123 -9638
rect 44167 -9682 44223 -9638
rect 44267 -9682 44323 -9638
rect 44367 -9682 44423 -9638
rect 44467 -9682 44523 -9638
rect 44567 -9682 44623 -9638
rect 44667 -9682 44723 -9638
rect 44767 -9682 47953 -9638
rect 34207 -9738 47953 -9682
rect 34207 -9782 37223 -9738
rect 37267 -9782 37323 -9738
rect 37367 -9782 37423 -9738
rect 37467 -9782 37523 -9738
rect 37567 -9782 37623 -9738
rect 37667 -9782 37723 -9738
rect 37767 -9782 37823 -9738
rect 37867 -9782 37923 -9738
rect 37967 -9782 38023 -9738
rect 38067 -9782 38123 -9738
rect 38167 -9782 38223 -9738
rect 38267 -9782 38323 -9738
rect 38367 -9782 38423 -9738
rect 38467 -9782 38523 -9738
rect 38567 -9782 38623 -9738
rect 38667 -9782 38723 -9738
rect 38767 -9782 39223 -9738
rect 39267 -9782 39323 -9738
rect 39367 -9782 39423 -9738
rect 39467 -9782 39523 -9738
rect 39567 -9782 39623 -9738
rect 39667 -9782 39723 -9738
rect 39767 -9782 39823 -9738
rect 39867 -9782 39923 -9738
rect 39967 -9782 40023 -9738
rect 40067 -9782 40123 -9738
rect 40167 -9782 40223 -9738
rect 40267 -9782 40323 -9738
rect 40367 -9782 40423 -9738
rect 40467 -9782 40523 -9738
rect 40567 -9782 40623 -9738
rect 40667 -9782 40723 -9738
rect 40767 -9782 41223 -9738
rect 41267 -9782 41323 -9738
rect 41367 -9782 41423 -9738
rect 41467 -9782 41523 -9738
rect 41567 -9782 41623 -9738
rect 41667 -9782 41723 -9738
rect 41767 -9782 41823 -9738
rect 41867 -9782 41923 -9738
rect 41967 -9782 42023 -9738
rect 42067 -9782 42123 -9738
rect 42167 -9782 42223 -9738
rect 42267 -9782 42323 -9738
rect 42367 -9782 42423 -9738
rect 42467 -9782 42523 -9738
rect 42567 -9782 42623 -9738
rect 42667 -9782 42723 -9738
rect 42767 -9782 43223 -9738
rect 43267 -9782 43323 -9738
rect 43367 -9782 43423 -9738
rect 43467 -9782 43523 -9738
rect 43567 -9782 43623 -9738
rect 43667 -9782 43723 -9738
rect 43767 -9782 43823 -9738
rect 43867 -9782 43923 -9738
rect 43967 -9782 44023 -9738
rect 44067 -9782 44123 -9738
rect 44167 -9782 44223 -9738
rect 44267 -9782 44323 -9738
rect 44367 -9782 44423 -9738
rect 44467 -9782 44523 -9738
rect 44567 -9782 44623 -9738
rect 44667 -9782 44723 -9738
rect 44767 -9782 47953 -9738
rect 34207 -9838 47953 -9782
rect 34207 -9882 37223 -9838
rect 37267 -9882 37323 -9838
rect 37367 -9882 37423 -9838
rect 37467 -9882 37523 -9838
rect 37567 -9882 37623 -9838
rect 37667 -9882 37723 -9838
rect 37767 -9882 37823 -9838
rect 37867 -9882 37923 -9838
rect 37967 -9882 38023 -9838
rect 38067 -9882 38123 -9838
rect 38167 -9882 38223 -9838
rect 38267 -9882 38323 -9838
rect 38367 -9882 38423 -9838
rect 38467 -9882 38523 -9838
rect 38567 -9882 38623 -9838
rect 38667 -9882 38723 -9838
rect 38767 -9882 39223 -9838
rect 39267 -9882 39323 -9838
rect 39367 -9882 39423 -9838
rect 39467 -9882 39523 -9838
rect 39567 -9882 39623 -9838
rect 39667 -9882 39723 -9838
rect 39767 -9882 39823 -9838
rect 39867 -9882 39923 -9838
rect 39967 -9882 40023 -9838
rect 40067 -9882 40123 -9838
rect 40167 -9882 40223 -9838
rect 40267 -9882 40323 -9838
rect 40367 -9882 40423 -9838
rect 40467 -9882 40523 -9838
rect 40567 -9882 40623 -9838
rect 40667 -9882 40723 -9838
rect 40767 -9882 41223 -9838
rect 41267 -9882 41323 -9838
rect 41367 -9882 41423 -9838
rect 41467 -9882 41523 -9838
rect 41567 -9882 41623 -9838
rect 41667 -9882 41723 -9838
rect 41767 -9882 41823 -9838
rect 41867 -9882 41923 -9838
rect 41967 -9882 42023 -9838
rect 42067 -9882 42123 -9838
rect 42167 -9882 42223 -9838
rect 42267 -9882 42323 -9838
rect 42367 -9882 42423 -9838
rect 42467 -9882 42523 -9838
rect 42567 -9882 42623 -9838
rect 42667 -9882 42723 -9838
rect 42767 -9882 43223 -9838
rect 43267 -9882 43323 -9838
rect 43367 -9882 43423 -9838
rect 43467 -9882 43523 -9838
rect 43567 -9882 43623 -9838
rect 43667 -9882 43723 -9838
rect 43767 -9882 43823 -9838
rect 43867 -9882 43923 -9838
rect 43967 -9882 44023 -9838
rect 44067 -9882 44123 -9838
rect 44167 -9882 44223 -9838
rect 44267 -9882 44323 -9838
rect 44367 -9882 44423 -9838
rect 44467 -9882 44523 -9838
rect 44567 -9882 44623 -9838
rect 44667 -9882 44723 -9838
rect 44767 -9882 47953 -9838
rect 34207 -9938 47953 -9882
rect 34207 -9982 37223 -9938
rect 37267 -9982 37323 -9938
rect 37367 -9982 37423 -9938
rect 37467 -9982 37523 -9938
rect 37567 -9982 37623 -9938
rect 37667 -9982 37723 -9938
rect 37767 -9982 37823 -9938
rect 37867 -9982 37923 -9938
rect 37967 -9982 38023 -9938
rect 38067 -9982 38123 -9938
rect 38167 -9982 38223 -9938
rect 38267 -9982 38323 -9938
rect 38367 -9982 38423 -9938
rect 38467 -9982 38523 -9938
rect 38567 -9982 38623 -9938
rect 38667 -9982 38723 -9938
rect 38767 -9982 39223 -9938
rect 39267 -9982 39323 -9938
rect 39367 -9982 39423 -9938
rect 39467 -9982 39523 -9938
rect 39567 -9982 39623 -9938
rect 39667 -9982 39723 -9938
rect 39767 -9982 39823 -9938
rect 39867 -9982 39923 -9938
rect 39967 -9982 40023 -9938
rect 40067 -9982 40123 -9938
rect 40167 -9982 40223 -9938
rect 40267 -9982 40323 -9938
rect 40367 -9982 40423 -9938
rect 40467 -9982 40523 -9938
rect 40567 -9982 40623 -9938
rect 40667 -9982 40723 -9938
rect 40767 -9982 41223 -9938
rect 41267 -9982 41323 -9938
rect 41367 -9982 41423 -9938
rect 41467 -9982 41523 -9938
rect 41567 -9982 41623 -9938
rect 41667 -9982 41723 -9938
rect 41767 -9982 41823 -9938
rect 41867 -9982 41923 -9938
rect 41967 -9982 42023 -9938
rect 42067 -9982 42123 -9938
rect 42167 -9982 42223 -9938
rect 42267 -9982 42323 -9938
rect 42367 -9982 42423 -9938
rect 42467 -9982 42523 -9938
rect 42567 -9982 42623 -9938
rect 42667 -9982 42723 -9938
rect 42767 -9982 43223 -9938
rect 43267 -9982 43323 -9938
rect 43367 -9982 43423 -9938
rect 43467 -9982 43523 -9938
rect 43567 -9982 43623 -9938
rect 43667 -9982 43723 -9938
rect 43767 -9982 43823 -9938
rect 43867 -9982 43923 -9938
rect 43967 -9982 44023 -9938
rect 44067 -9982 44123 -9938
rect 44167 -9982 44223 -9938
rect 44267 -9982 44323 -9938
rect 44367 -9982 44423 -9938
rect 44467 -9982 44523 -9938
rect 44567 -9982 44623 -9938
rect 44667 -9982 44723 -9938
rect 44767 -9982 47953 -9938
rect 34207 -10038 47953 -9982
rect 34207 -10082 37223 -10038
rect 37267 -10082 37323 -10038
rect 37367 -10082 37423 -10038
rect 37467 -10082 37523 -10038
rect 37567 -10082 37623 -10038
rect 37667 -10082 37723 -10038
rect 37767 -10082 37823 -10038
rect 37867 -10082 37923 -10038
rect 37967 -10082 38023 -10038
rect 38067 -10082 38123 -10038
rect 38167 -10082 38223 -10038
rect 38267 -10082 38323 -10038
rect 38367 -10082 38423 -10038
rect 38467 -10082 38523 -10038
rect 38567 -10082 38623 -10038
rect 38667 -10082 38723 -10038
rect 38767 -10082 39223 -10038
rect 39267 -10082 39323 -10038
rect 39367 -10082 39423 -10038
rect 39467 -10082 39523 -10038
rect 39567 -10082 39623 -10038
rect 39667 -10082 39723 -10038
rect 39767 -10082 39823 -10038
rect 39867 -10082 39923 -10038
rect 39967 -10082 40023 -10038
rect 40067 -10082 40123 -10038
rect 40167 -10082 40223 -10038
rect 40267 -10082 40323 -10038
rect 40367 -10082 40423 -10038
rect 40467 -10082 40523 -10038
rect 40567 -10082 40623 -10038
rect 40667 -10082 40723 -10038
rect 40767 -10082 41223 -10038
rect 41267 -10082 41323 -10038
rect 41367 -10082 41423 -10038
rect 41467 -10082 41523 -10038
rect 41567 -10082 41623 -10038
rect 41667 -10082 41723 -10038
rect 41767 -10082 41823 -10038
rect 41867 -10082 41923 -10038
rect 41967 -10082 42023 -10038
rect 42067 -10082 42123 -10038
rect 42167 -10082 42223 -10038
rect 42267 -10082 42323 -10038
rect 42367 -10082 42423 -10038
rect 42467 -10082 42523 -10038
rect 42567 -10082 42623 -10038
rect 42667 -10082 42723 -10038
rect 42767 -10082 43223 -10038
rect 43267 -10082 43323 -10038
rect 43367 -10082 43423 -10038
rect 43467 -10082 43523 -10038
rect 43567 -10082 43623 -10038
rect 43667 -10082 43723 -10038
rect 43767 -10082 43823 -10038
rect 43867 -10082 43923 -10038
rect 43967 -10082 44023 -10038
rect 44067 -10082 44123 -10038
rect 44167 -10082 44223 -10038
rect 44267 -10082 44323 -10038
rect 44367 -10082 44423 -10038
rect 44467 -10082 44523 -10038
rect 44567 -10082 44623 -10038
rect 44667 -10082 44723 -10038
rect 44767 -10082 47953 -10038
rect 34207 -10138 47953 -10082
rect 34207 -10182 37223 -10138
rect 37267 -10182 37323 -10138
rect 37367 -10182 37423 -10138
rect 37467 -10182 37523 -10138
rect 37567 -10182 37623 -10138
rect 37667 -10182 37723 -10138
rect 37767 -10182 37823 -10138
rect 37867 -10182 37923 -10138
rect 37967 -10182 38023 -10138
rect 38067 -10182 38123 -10138
rect 38167 -10182 38223 -10138
rect 38267 -10182 38323 -10138
rect 38367 -10182 38423 -10138
rect 38467 -10182 38523 -10138
rect 38567 -10182 38623 -10138
rect 38667 -10182 38723 -10138
rect 38767 -10182 39223 -10138
rect 39267 -10182 39323 -10138
rect 39367 -10182 39423 -10138
rect 39467 -10182 39523 -10138
rect 39567 -10182 39623 -10138
rect 39667 -10182 39723 -10138
rect 39767 -10182 39823 -10138
rect 39867 -10182 39923 -10138
rect 39967 -10182 40023 -10138
rect 40067 -10182 40123 -10138
rect 40167 -10182 40223 -10138
rect 40267 -10182 40323 -10138
rect 40367 -10182 40423 -10138
rect 40467 -10182 40523 -10138
rect 40567 -10182 40623 -10138
rect 40667 -10182 40723 -10138
rect 40767 -10182 41223 -10138
rect 41267 -10182 41323 -10138
rect 41367 -10182 41423 -10138
rect 41467 -10182 41523 -10138
rect 41567 -10182 41623 -10138
rect 41667 -10182 41723 -10138
rect 41767 -10182 41823 -10138
rect 41867 -10182 41923 -10138
rect 41967 -10182 42023 -10138
rect 42067 -10182 42123 -10138
rect 42167 -10182 42223 -10138
rect 42267 -10182 42323 -10138
rect 42367 -10182 42423 -10138
rect 42467 -10182 42523 -10138
rect 42567 -10182 42623 -10138
rect 42667 -10182 42723 -10138
rect 42767 -10182 43223 -10138
rect 43267 -10182 43323 -10138
rect 43367 -10182 43423 -10138
rect 43467 -10182 43523 -10138
rect 43567 -10182 43623 -10138
rect 43667 -10182 43723 -10138
rect 43767 -10182 43823 -10138
rect 43867 -10182 43923 -10138
rect 43967 -10182 44023 -10138
rect 44067 -10182 44123 -10138
rect 44167 -10182 44223 -10138
rect 44267 -10182 44323 -10138
rect 44367 -10182 44423 -10138
rect 44467 -10182 44523 -10138
rect 44567 -10182 44623 -10138
rect 44667 -10182 44723 -10138
rect 44767 -10182 47953 -10138
rect 34207 -10238 47953 -10182
rect 34207 -10282 37223 -10238
rect 37267 -10282 37323 -10238
rect 37367 -10282 37423 -10238
rect 37467 -10282 37523 -10238
rect 37567 -10282 37623 -10238
rect 37667 -10282 37723 -10238
rect 37767 -10282 37823 -10238
rect 37867 -10282 37923 -10238
rect 37967 -10282 38023 -10238
rect 38067 -10282 38123 -10238
rect 38167 -10282 38223 -10238
rect 38267 -10282 38323 -10238
rect 38367 -10282 38423 -10238
rect 38467 -10282 38523 -10238
rect 38567 -10282 38623 -10238
rect 38667 -10282 38723 -10238
rect 38767 -10282 39223 -10238
rect 39267 -10282 39323 -10238
rect 39367 -10282 39423 -10238
rect 39467 -10282 39523 -10238
rect 39567 -10282 39623 -10238
rect 39667 -10282 39723 -10238
rect 39767 -10282 39823 -10238
rect 39867 -10282 39923 -10238
rect 39967 -10282 40023 -10238
rect 40067 -10282 40123 -10238
rect 40167 -10282 40223 -10238
rect 40267 -10282 40323 -10238
rect 40367 -10282 40423 -10238
rect 40467 -10282 40523 -10238
rect 40567 -10282 40623 -10238
rect 40667 -10282 40723 -10238
rect 40767 -10282 41223 -10238
rect 41267 -10282 41323 -10238
rect 41367 -10282 41423 -10238
rect 41467 -10282 41523 -10238
rect 41567 -10282 41623 -10238
rect 41667 -10282 41723 -10238
rect 41767 -10282 41823 -10238
rect 41867 -10282 41923 -10238
rect 41967 -10282 42023 -10238
rect 42067 -10282 42123 -10238
rect 42167 -10282 42223 -10238
rect 42267 -10282 42323 -10238
rect 42367 -10282 42423 -10238
rect 42467 -10282 42523 -10238
rect 42567 -10282 42623 -10238
rect 42667 -10282 42723 -10238
rect 42767 -10282 43223 -10238
rect 43267 -10282 43323 -10238
rect 43367 -10282 43423 -10238
rect 43467 -10282 43523 -10238
rect 43567 -10282 43623 -10238
rect 43667 -10282 43723 -10238
rect 43767 -10282 43823 -10238
rect 43867 -10282 43923 -10238
rect 43967 -10282 44023 -10238
rect 44067 -10282 44123 -10238
rect 44167 -10282 44223 -10238
rect 44267 -10282 44323 -10238
rect 44367 -10282 44423 -10238
rect 44467 -10282 44523 -10238
rect 44567 -10282 44623 -10238
rect 44667 -10282 44723 -10238
rect 44767 -10282 47953 -10238
rect 34207 -10338 47953 -10282
rect 34207 -10382 37223 -10338
rect 37267 -10382 37323 -10338
rect 37367 -10382 37423 -10338
rect 37467 -10382 37523 -10338
rect 37567 -10382 37623 -10338
rect 37667 -10382 37723 -10338
rect 37767 -10382 37823 -10338
rect 37867 -10382 37923 -10338
rect 37967 -10382 38023 -10338
rect 38067 -10382 38123 -10338
rect 38167 -10382 38223 -10338
rect 38267 -10382 38323 -10338
rect 38367 -10382 38423 -10338
rect 38467 -10382 38523 -10338
rect 38567 -10382 38623 -10338
rect 38667 -10382 38723 -10338
rect 38767 -10382 39223 -10338
rect 39267 -10382 39323 -10338
rect 39367 -10382 39423 -10338
rect 39467 -10382 39523 -10338
rect 39567 -10382 39623 -10338
rect 39667 -10382 39723 -10338
rect 39767 -10382 39823 -10338
rect 39867 -10382 39923 -10338
rect 39967 -10382 40023 -10338
rect 40067 -10382 40123 -10338
rect 40167 -10382 40223 -10338
rect 40267 -10382 40323 -10338
rect 40367 -10382 40423 -10338
rect 40467 -10382 40523 -10338
rect 40567 -10382 40623 -10338
rect 40667 -10382 40723 -10338
rect 40767 -10382 41223 -10338
rect 41267 -10382 41323 -10338
rect 41367 -10382 41423 -10338
rect 41467 -10382 41523 -10338
rect 41567 -10382 41623 -10338
rect 41667 -10382 41723 -10338
rect 41767 -10382 41823 -10338
rect 41867 -10382 41923 -10338
rect 41967 -10382 42023 -10338
rect 42067 -10382 42123 -10338
rect 42167 -10382 42223 -10338
rect 42267 -10382 42323 -10338
rect 42367 -10382 42423 -10338
rect 42467 -10382 42523 -10338
rect 42567 -10382 42623 -10338
rect 42667 -10382 42723 -10338
rect 42767 -10382 43223 -10338
rect 43267 -10382 43323 -10338
rect 43367 -10382 43423 -10338
rect 43467 -10382 43523 -10338
rect 43567 -10382 43623 -10338
rect 43667 -10382 43723 -10338
rect 43767 -10382 43823 -10338
rect 43867 -10382 43923 -10338
rect 43967 -10382 44023 -10338
rect 44067 -10382 44123 -10338
rect 44167 -10382 44223 -10338
rect 44267 -10382 44323 -10338
rect 44367 -10382 44423 -10338
rect 44467 -10382 44523 -10338
rect 44567 -10382 44623 -10338
rect 44667 -10382 44723 -10338
rect 44767 -10382 47953 -10338
rect 34207 -10438 47953 -10382
rect 34207 -10482 37223 -10438
rect 37267 -10482 37323 -10438
rect 37367 -10482 37423 -10438
rect 37467 -10482 37523 -10438
rect 37567 -10482 37623 -10438
rect 37667 -10482 37723 -10438
rect 37767 -10482 37823 -10438
rect 37867 -10482 37923 -10438
rect 37967 -10482 38023 -10438
rect 38067 -10482 38123 -10438
rect 38167 -10482 38223 -10438
rect 38267 -10482 38323 -10438
rect 38367 -10482 38423 -10438
rect 38467 -10482 38523 -10438
rect 38567 -10482 38623 -10438
rect 38667 -10482 38723 -10438
rect 38767 -10482 39223 -10438
rect 39267 -10482 39323 -10438
rect 39367 -10482 39423 -10438
rect 39467 -10482 39523 -10438
rect 39567 -10482 39623 -10438
rect 39667 -10482 39723 -10438
rect 39767 -10482 39823 -10438
rect 39867 -10482 39923 -10438
rect 39967 -10482 40023 -10438
rect 40067 -10482 40123 -10438
rect 40167 -10482 40223 -10438
rect 40267 -10482 40323 -10438
rect 40367 -10482 40423 -10438
rect 40467 -10482 40523 -10438
rect 40567 -10482 40623 -10438
rect 40667 -10482 40723 -10438
rect 40767 -10482 41223 -10438
rect 41267 -10482 41323 -10438
rect 41367 -10482 41423 -10438
rect 41467 -10482 41523 -10438
rect 41567 -10482 41623 -10438
rect 41667 -10482 41723 -10438
rect 41767 -10482 41823 -10438
rect 41867 -10482 41923 -10438
rect 41967 -10482 42023 -10438
rect 42067 -10482 42123 -10438
rect 42167 -10482 42223 -10438
rect 42267 -10482 42323 -10438
rect 42367 -10482 42423 -10438
rect 42467 -10482 42523 -10438
rect 42567 -10482 42623 -10438
rect 42667 -10482 42723 -10438
rect 42767 -10482 43223 -10438
rect 43267 -10482 43323 -10438
rect 43367 -10482 43423 -10438
rect 43467 -10482 43523 -10438
rect 43567 -10482 43623 -10438
rect 43667 -10482 43723 -10438
rect 43767 -10482 43823 -10438
rect 43867 -10482 43923 -10438
rect 43967 -10482 44023 -10438
rect 44067 -10482 44123 -10438
rect 44167 -10482 44223 -10438
rect 44267 -10482 44323 -10438
rect 44367 -10482 44423 -10438
rect 44467 -10482 44523 -10438
rect 44567 -10482 44623 -10438
rect 44667 -10482 44723 -10438
rect 44767 -10482 47953 -10438
rect 34207 -10538 47953 -10482
rect 34207 -10582 37223 -10538
rect 37267 -10582 37323 -10538
rect 37367 -10582 37423 -10538
rect 37467 -10582 37523 -10538
rect 37567 -10582 37623 -10538
rect 37667 -10582 37723 -10538
rect 37767 -10582 37823 -10538
rect 37867 -10582 37923 -10538
rect 37967 -10582 38023 -10538
rect 38067 -10582 38123 -10538
rect 38167 -10582 38223 -10538
rect 38267 -10582 38323 -10538
rect 38367 -10582 38423 -10538
rect 38467 -10582 38523 -10538
rect 38567 -10582 38623 -10538
rect 38667 -10582 38723 -10538
rect 38767 -10582 39223 -10538
rect 39267 -10582 39323 -10538
rect 39367 -10582 39423 -10538
rect 39467 -10582 39523 -10538
rect 39567 -10582 39623 -10538
rect 39667 -10582 39723 -10538
rect 39767 -10582 39823 -10538
rect 39867 -10582 39923 -10538
rect 39967 -10582 40023 -10538
rect 40067 -10582 40123 -10538
rect 40167 -10582 40223 -10538
rect 40267 -10582 40323 -10538
rect 40367 -10582 40423 -10538
rect 40467 -10582 40523 -10538
rect 40567 -10582 40623 -10538
rect 40667 -10582 40723 -10538
rect 40767 -10582 41223 -10538
rect 41267 -10582 41323 -10538
rect 41367 -10582 41423 -10538
rect 41467 -10582 41523 -10538
rect 41567 -10582 41623 -10538
rect 41667 -10582 41723 -10538
rect 41767 -10582 41823 -10538
rect 41867 -10582 41923 -10538
rect 41967 -10582 42023 -10538
rect 42067 -10582 42123 -10538
rect 42167 -10582 42223 -10538
rect 42267 -10582 42323 -10538
rect 42367 -10582 42423 -10538
rect 42467 -10582 42523 -10538
rect 42567 -10582 42623 -10538
rect 42667 -10582 42723 -10538
rect 42767 -10582 43223 -10538
rect 43267 -10582 43323 -10538
rect 43367 -10582 43423 -10538
rect 43467 -10582 43523 -10538
rect 43567 -10582 43623 -10538
rect 43667 -10582 43723 -10538
rect 43767 -10582 43823 -10538
rect 43867 -10582 43923 -10538
rect 43967 -10582 44023 -10538
rect 44067 -10582 44123 -10538
rect 44167 -10582 44223 -10538
rect 44267 -10582 44323 -10538
rect 44367 -10582 44423 -10538
rect 44467 -10582 44523 -10538
rect 44567 -10582 44623 -10538
rect 44667 -10582 44723 -10538
rect 44767 -10582 47953 -10538
rect 34207 -10638 47953 -10582
rect 34207 -10682 37223 -10638
rect 37267 -10682 37323 -10638
rect 37367 -10682 37423 -10638
rect 37467 -10682 37523 -10638
rect 37567 -10682 37623 -10638
rect 37667 -10682 37723 -10638
rect 37767 -10682 37823 -10638
rect 37867 -10682 37923 -10638
rect 37967 -10682 38023 -10638
rect 38067 -10682 38123 -10638
rect 38167 -10682 38223 -10638
rect 38267 -10682 38323 -10638
rect 38367 -10682 38423 -10638
rect 38467 -10682 38523 -10638
rect 38567 -10682 38623 -10638
rect 38667 -10682 38723 -10638
rect 38767 -10682 39223 -10638
rect 39267 -10682 39323 -10638
rect 39367 -10682 39423 -10638
rect 39467 -10682 39523 -10638
rect 39567 -10682 39623 -10638
rect 39667 -10682 39723 -10638
rect 39767 -10682 39823 -10638
rect 39867 -10682 39923 -10638
rect 39967 -10682 40023 -10638
rect 40067 -10682 40123 -10638
rect 40167 -10682 40223 -10638
rect 40267 -10682 40323 -10638
rect 40367 -10682 40423 -10638
rect 40467 -10682 40523 -10638
rect 40567 -10682 40623 -10638
rect 40667 -10682 40723 -10638
rect 40767 -10682 41223 -10638
rect 41267 -10682 41323 -10638
rect 41367 -10682 41423 -10638
rect 41467 -10682 41523 -10638
rect 41567 -10682 41623 -10638
rect 41667 -10682 41723 -10638
rect 41767 -10682 41823 -10638
rect 41867 -10682 41923 -10638
rect 41967 -10682 42023 -10638
rect 42067 -10682 42123 -10638
rect 42167 -10682 42223 -10638
rect 42267 -10682 42323 -10638
rect 42367 -10682 42423 -10638
rect 42467 -10682 42523 -10638
rect 42567 -10682 42623 -10638
rect 42667 -10682 42723 -10638
rect 42767 -10682 43223 -10638
rect 43267 -10682 43323 -10638
rect 43367 -10682 43423 -10638
rect 43467 -10682 43523 -10638
rect 43567 -10682 43623 -10638
rect 43667 -10682 43723 -10638
rect 43767 -10682 43823 -10638
rect 43867 -10682 43923 -10638
rect 43967 -10682 44023 -10638
rect 44067 -10682 44123 -10638
rect 44167 -10682 44223 -10638
rect 44267 -10682 44323 -10638
rect 44367 -10682 44423 -10638
rect 44467 -10682 44523 -10638
rect 44567 -10682 44623 -10638
rect 44667 -10682 44723 -10638
rect 44767 -10682 47953 -10638
rect 34207 -10738 47953 -10682
rect 34207 -10782 37223 -10738
rect 37267 -10782 37323 -10738
rect 37367 -10782 37423 -10738
rect 37467 -10782 37523 -10738
rect 37567 -10782 37623 -10738
rect 37667 -10782 37723 -10738
rect 37767 -10782 37823 -10738
rect 37867 -10782 37923 -10738
rect 37967 -10782 38023 -10738
rect 38067 -10782 38123 -10738
rect 38167 -10782 38223 -10738
rect 38267 -10782 38323 -10738
rect 38367 -10782 38423 -10738
rect 38467 -10782 38523 -10738
rect 38567 -10782 38623 -10738
rect 38667 -10782 38723 -10738
rect 38767 -10782 39223 -10738
rect 39267 -10782 39323 -10738
rect 39367 -10782 39423 -10738
rect 39467 -10782 39523 -10738
rect 39567 -10782 39623 -10738
rect 39667 -10782 39723 -10738
rect 39767 -10782 39823 -10738
rect 39867 -10782 39923 -10738
rect 39967 -10782 40023 -10738
rect 40067 -10782 40123 -10738
rect 40167 -10782 40223 -10738
rect 40267 -10782 40323 -10738
rect 40367 -10782 40423 -10738
rect 40467 -10782 40523 -10738
rect 40567 -10782 40623 -10738
rect 40667 -10782 40723 -10738
rect 40767 -10782 41223 -10738
rect 41267 -10782 41323 -10738
rect 41367 -10782 41423 -10738
rect 41467 -10782 41523 -10738
rect 41567 -10782 41623 -10738
rect 41667 -10782 41723 -10738
rect 41767 -10782 41823 -10738
rect 41867 -10782 41923 -10738
rect 41967 -10782 42023 -10738
rect 42067 -10782 42123 -10738
rect 42167 -10782 42223 -10738
rect 42267 -10782 42323 -10738
rect 42367 -10782 42423 -10738
rect 42467 -10782 42523 -10738
rect 42567 -10782 42623 -10738
rect 42667 -10782 42723 -10738
rect 42767 -10782 43223 -10738
rect 43267 -10782 43323 -10738
rect 43367 -10782 43423 -10738
rect 43467 -10782 43523 -10738
rect 43567 -10782 43623 -10738
rect 43667 -10782 43723 -10738
rect 43767 -10782 43823 -10738
rect 43867 -10782 43923 -10738
rect 43967 -10782 44023 -10738
rect 44067 -10782 44123 -10738
rect 44167 -10782 44223 -10738
rect 44267 -10782 44323 -10738
rect 44367 -10782 44423 -10738
rect 44467 -10782 44523 -10738
rect 44567 -10782 44623 -10738
rect 44667 -10782 44723 -10738
rect 44767 -10782 47953 -10738
rect 34207 -10838 47953 -10782
rect 34207 -10882 37223 -10838
rect 37267 -10882 37323 -10838
rect 37367 -10882 37423 -10838
rect 37467 -10882 37523 -10838
rect 37567 -10882 37623 -10838
rect 37667 -10882 37723 -10838
rect 37767 -10882 37823 -10838
rect 37867 -10882 37923 -10838
rect 37967 -10882 38023 -10838
rect 38067 -10882 38123 -10838
rect 38167 -10882 38223 -10838
rect 38267 -10882 38323 -10838
rect 38367 -10882 38423 -10838
rect 38467 -10882 38523 -10838
rect 38567 -10882 38623 -10838
rect 38667 -10882 38723 -10838
rect 38767 -10882 39223 -10838
rect 39267 -10882 39323 -10838
rect 39367 -10882 39423 -10838
rect 39467 -10882 39523 -10838
rect 39567 -10882 39623 -10838
rect 39667 -10882 39723 -10838
rect 39767 -10882 39823 -10838
rect 39867 -10882 39923 -10838
rect 39967 -10882 40023 -10838
rect 40067 -10882 40123 -10838
rect 40167 -10882 40223 -10838
rect 40267 -10882 40323 -10838
rect 40367 -10882 40423 -10838
rect 40467 -10882 40523 -10838
rect 40567 -10882 40623 -10838
rect 40667 -10882 40723 -10838
rect 40767 -10882 41223 -10838
rect 41267 -10882 41323 -10838
rect 41367 -10882 41423 -10838
rect 41467 -10882 41523 -10838
rect 41567 -10882 41623 -10838
rect 41667 -10882 41723 -10838
rect 41767 -10882 41823 -10838
rect 41867 -10882 41923 -10838
rect 41967 -10882 42023 -10838
rect 42067 -10882 42123 -10838
rect 42167 -10882 42223 -10838
rect 42267 -10882 42323 -10838
rect 42367 -10882 42423 -10838
rect 42467 -10882 42523 -10838
rect 42567 -10882 42623 -10838
rect 42667 -10882 42723 -10838
rect 42767 -10882 43223 -10838
rect 43267 -10882 43323 -10838
rect 43367 -10882 43423 -10838
rect 43467 -10882 43523 -10838
rect 43567 -10882 43623 -10838
rect 43667 -10882 43723 -10838
rect 43767 -10882 43823 -10838
rect 43867 -10882 43923 -10838
rect 43967 -10882 44023 -10838
rect 44067 -10882 44123 -10838
rect 44167 -10882 44223 -10838
rect 44267 -10882 44323 -10838
rect 44367 -10882 44423 -10838
rect 44467 -10882 44523 -10838
rect 44567 -10882 44623 -10838
rect 44667 -10882 44723 -10838
rect 44767 -10882 47953 -10838
rect 34207 -10938 47953 -10882
rect 34207 -10982 37223 -10938
rect 37267 -10982 37323 -10938
rect 37367 -10982 37423 -10938
rect 37467 -10982 37523 -10938
rect 37567 -10982 37623 -10938
rect 37667 -10982 37723 -10938
rect 37767 -10982 37823 -10938
rect 37867 -10982 37923 -10938
rect 37967 -10982 38023 -10938
rect 38067 -10982 38123 -10938
rect 38167 -10982 38223 -10938
rect 38267 -10982 38323 -10938
rect 38367 -10982 38423 -10938
rect 38467 -10982 38523 -10938
rect 38567 -10982 38623 -10938
rect 38667 -10982 38723 -10938
rect 38767 -10982 39223 -10938
rect 39267 -10982 39323 -10938
rect 39367 -10982 39423 -10938
rect 39467 -10982 39523 -10938
rect 39567 -10982 39623 -10938
rect 39667 -10982 39723 -10938
rect 39767 -10982 39823 -10938
rect 39867 -10982 39923 -10938
rect 39967 -10982 40023 -10938
rect 40067 -10982 40123 -10938
rect 40167 -10982 40223 -10938
rect 40267 -10982 40323 -10938
rect 40367 -10982 40423 -10938
rect 40467 -10982 40523 -10938
rect 40567 -10982 40623 -10938
rect 40667 -10982 40723 -10938
rect 40767 -10982 41223 -10938
rect 41267 -10982 41323 -10938
rect 41367 -10982 41423 -10938
rect 41467 -10982 41523 -10938
rect 41567 -10982 41623 -10938
rect 41667 -10982 41723 -10938
rect 41767 -10982 41823 -10938
rect 41867 -10982 41923 -10938
rect 41967 -10982 42023 -10938
rect 42067 -10982 42123 -10938
rect 42167 -10982 42223 -10938
rect 42267 -10982 42323 -10938
rect 42367 -10982 42423 -10938
rect 42467 -10982 42523 -10938
rect 42567 -10982 42623 -10938
rect 42667 -10982 42723 -10938
rect 42767 -10982 43223 -10938
rect 43267 -10982 43323 -10938
rect 43367 -10982 43423 -10938
rect 43467 -10982 43523 -10938
rect 43567 -10982 43623 -10938
rect 43667 -10982 43723 -10938
rect 43767 -10982 43823 -10938
rect 43867 -10982 43923 -10938
rect 43967 -10982 44023 -10938
rect 44067 -10982 44123 -10938
rect 44167 -10982 44223 -10938
rect 44267 -10982 44323 -10938
rect 44367 -10982 44423 -10938
rect 44467 -10982 44523 -10938
rect 44567 -10982 44623 -10938
rect 44667 -10982 44723 -10938
rect 44767 -10982 47953 -10938
rect 34207 -11038 47953 -10982
rect 34207 -11082 37223 -11038
rect 37267 -11082 37323 -11038
rect 37367 -11082 37423 -11038
rect 37467 -11082 37523 -11038
rect 37567 -11082 37623 -11038
rect 37667 -11082 37723 -11038
rect 37767 -11082 37823 -11038
rect 37867 -11082 37923 -11038
rect 37967 -11082 38023 -11038
rect 38067 -11082 38123 -11038
rect 38167 -11082 38223 -11038
rect 38267 -11082 38323 -11038
rect 38367 -11082 38423 -11038
rect 38467 -11082 38523 -11038
rect 38567 -11082 38623 -11038
rect 38667 -11082 38723 -11038
rect 38767 -11082 39223 -11038
rect 39267 -11082 39323 -11038
rect 39367 -11082 39423 -11038
rect 39467 -11082 39523 -11038
rect 39567 -11082 39623 -11038
rect 39667 -11082 39723 -11038
rect 39767 -11082 39823 -11038
rect 39867 -11082 39923 -11038
rect 39967 -11082 40023 -11038
rect 40067 -11082 40123 -11038
rect 40167 -11082 40223 -11038
rect 40267 -11082 40323 -11038
rect 40367 -11082 40423 -11038
rect 40467 -11082 40523 -11038
rect 40567 -11082 40623 -11038
rect 40667 -11082 40723 -11038
rect 40767 -11082 41223 -11038
rect 41267 -11082 41323 -11038
rect 41367 -11082 41423 -11038
rect 41467 -11082 41523 -11038
rect 41567 -11082 41623 -11038
rect 41667 -11082 41723 -11038
rect 41767 -11082 41823 -11038
rect 41867 -11082 41923 -11038
rect 41967 -11082 42023 -11038
rect 42067 -11082 42123 -11038
rect 42167 -11082 42223 -11038
rect 42267 -11082 42323 -11038
rect 42367 -11082 42423 -11038
rect 42467 -11082 42523 -11038
rect 42567 -11082 42623 -11038
rect 42667 -11082 42723 -11038
rect 42767 -11082 43223 -11038
rect 43267 -11082 43323 -11038
rect 43367 -11082 43423 -11038
rect 43467 -11082 43523 -11038
rect 43567 -11082 43623 -11038
rect 43667 -11082 43723 -11038
rect 43767 -11082 43823 -11038
rect 43867 -11082 43923 -11038
rect 43967 -11082 44023 -11038
rect 44067 -11082 44123 -11038
rect 44167 -11082 44223 -11038
rect 44267 -11082 44323 -11038
rect 44367 -11082 44423 -11038
rect 44467 -11082 44523 -11038
rect 44567 -11082 44623 -11038
rect 44667 -11082 44723 -11038
rect 44767 -11082 47953 -11038
rect 34207 -11138 47953 -11082
rect 34207 -11182 37223 -11138
rect 37267 -11182 37323 -11138
rect 37367 -11182 37423 -11138
rect 37467 -11182 37523 -11138
rect 37567 -11182 37623 -11138
rect 37667 -11182 37723 -11138
rect 37767 -11182 37823 -11138
rect 37867 -11182 37923 -11138
rect 37967 -11182 38023 -11138
rect 38067 -11182 38123 -11138
rect 38167 -11182 38223 -11138
rect 38267 -11182 38323 -11138
rect 38367 -11182 38423 -11138
rect 38467 -11182 38523 -11138
rect 38567 -11182 38623 -11138
rect 38667 -11182 38723 -11138
rect 38767 -11182 39223 -11138
rect 39267 -11182 39323 -11138
rect 39367 -11182 39423 -11138
rect 39467 -11182 39523 -11138
rect 39567 -11182 39623 -11138
rect 39667 -11182 39723 -11138
rect 39767 -11182 39823 -11138
rect 39867 -11182 39923 -11138
rect 39967 -11182 40023 -11138
rect 40067 -11182 40123 -11138
rect 40167 -11182 40223 -11138
rect 40267 -11182 40323 -11138
rect 40367 -11182 40423 -11138
rect 40467 -11182 40523 -11138
rect 40567 -11182 40623 -11138
rect 40667 -11182 40723 -11138
rect 40767 -11182 41223 -11138
rect 41267 -11182 41323 -11138
rect 41367 -11182 41423 -11138
rect 41467 -11182 41523 -11138
rect 41567 -11182 41623 -11138
rect 41667 -11182 41723 -11138
rect 41767 -11182 41823 -11138
rect 41867 -11182 41923 -11138
rect 41967 -11182 42023 -11138
rect 42067 -11182 42123 -11138
rect 42167 -11182 42223 -11138
rect 42267 -11182 42323 -11138
rect 42367 -11182 42423 -11138
rect 42467 -11182 42523 -11138
rect 42567 -11182 42623 -11138
rect 42667 -11182 42723 -11138
rect 42767 -11182 43223 -11138
rect 43267 -11182 43323 -11138
rect 43367 -11182 43423 -11138
rect 43467 -11182 43523 -11138
rect 43567 -11182 43623 -11138
rect 43667 -11182 43723 -11138
rect 43767 -11182 43823 -11138
rect 43867 -11182 43923 -11138
rect 43967 -11182 44023 -11138
rect 44067 -11182 44123 -11138
rect 44167 -11182 44223 -11138
rect 44267 -11182 44323 -11138
rect 44367 -11182 44423 -11138
rect 44467 -11182 44523 -11138
rect 44567 -11182 44623 -11138
rect 44667 -11182 44723 -11138
rect 44767 -11182 47953 -11138
rect -16409 -131295 -13354 -131251
rect -13310 -131295 -13254 -131251
rect -13210 -131295 -13154 -131251
rect -13110 -131295 -13054 -131251
rect -13010 -131295 -12954 -131251
rect -12910 -131295 -12854 -131251
rect -12810 -131295 -12754 -131251
rect -12710 -131295 -12654 -131251
rect -12610 -131295 -12554 -131251
rect -12510 -131295 -12454 -131251
rect -12410 -131295 -12354 -131251
rect -12310 -131295 -12254 -131251
rect -12210 -131295 -12154 -131251
rect -12110 -131295 -12054 -131251
rect -12010 -131295 -11954 -131251
rect -11910 -131295 -11854 -131251
rect -11810 -131295 -11354 -131251
rect -11310 -131295 -11254 -131251
rect -11210 -131295 -11154 -131251
rect -11110 -131295 -11054 -131251
rect -11010 -131295 -10954 -131251
rect -10910 -131295 -10854 -131251
rect -10810 -131295 -10754 -131251
rect -10710 -131295 -10654 -131251
rect -10610 -131295 -10554 -131251
rect -10510 -131295 -10454 -131251
rect -10410 -131295 -10354 -131251
rect -10310 -131295 -10254 -131251
rect -10210 -131295 -10154 -131251
rect -10110 -131295 -10054 -131251
rect -10010 -131295 -9954 -131251
rect -9910 -131295 -9854 -131251
rect -9810 -131295 -9354 -131251
rect -9310 -131295 -9254 -131251
rect -9210 -131295 -9154 -131251
rect -9110 -131295 -9054 -131251
rect -9010 -131295 -8954 -131251
rect -8910 -131295 -8854 -131251
rect -8810 -131295 -8754 -131251
rect -8710 -131295 -8654 -131251
rect -8610 -131295 -8554 -131251
rect -8510 -131295 -8454 -131251
rect -8410 -131295 -8354 -131251
rect -8310 -131295 -8254 -131251
rect -8210 -131295 -8154 -131251
rect -8110 -131295 -8054 -131251
rect -8010 -131295 -7954 -131251
rect -7910 -131295 -7854 -131251
rect -7810 -131295 -7354 -131251
rect -7310 -131295 -7254 -131251
rect -7210 -131295 -7154 -131251
rect -7110 -131295 -7054 -131251
rect -7010 -131295 -6954 -131251
rect -6910 -131295 -6854 -131251
rect -6810 -131295 -6754 -131251
rect -6710 -131295 -6654 -131251
rect -6610 -131295 -6554 -131251
rect -6510 -131295 -6454 -131251
rect -6410 -131295 -6354 -131251
rect -6310 -131295 -6254 -131251
rect -6210 -131295 -6154 -131251
rect -6110 -131295 -6054 -131251
rect -6010 -131295 -5954 -131251
rect -5910 -131295 -5854 -131251
rect -5810 -131295 -2893 -131251
rect -16409 -131351 -2893 -131295
rect -16409 -131395 -13354 -131351
rect -13310 -131395 -13254 -131351
rect -13210 -131395 -13154 -131351
rect -13110 -131395 -13054 -131351
rect -13010 -131395 -12954 -131351
rect -12910 -131395 -12854 -131351
rect -12810 -131395 -12754 -131351
rect -12710 -131395 -12654 -131351
rect -12610 -131395 -12554 -131351
rect -12510 -131395 -12454 -131351
rect -12410 -131395 -12354 -131351
rect -12310 -131395 -12254 -131351
rect -12210 -131395 -12154 -131351
rect -12110 -131395 -12054 -131351
rect -12010 -131395 -11954 -131351
rect -11910 -131395 -11854 -131351
rect -11810 -131395 -11354 -131351
rect -11310 -131395 -11254 -131351
rect -11210 -131395 -11154 -131351
rect -11110 -131395 -11054 -131351
rect -11010 -131395 -10954 -131351
rect -10910 -131395 -10854 -131351
rect -10810 -131395 -10754 -131351
rect -10710 -131395 -10654 -131351
rect -10610 -131395 -10554 -131351
rect -10510 -131395 -10454 -131351
rect -10410 -131395 -10354 -131351
rect -10310 -131395 -10254 -131351
rect -10210 -131395 -10154 -131351
rect -10110 -131395 -10054 -131351
rect -10010 -131395 -9954 -131351
rect -9910 -131395 -9854 -131351
rect -9810 -131395 -9354 -131351
rect -9310 -131395 -9254 -131351
rect -9210 -131395 -9154 -131351
rect -9110 -131395 -9054 -131351
rect -9010 -131395 -8954 -131351
rect -8910 -131395 -8854 -131351
rect -8810 -131395 -8754 -131351
rect -8710 -131395 -8654 -131351
rect -8610 -131395 -8554 -131351
rect -8510 -131395 -8454 -131351
rect -8410 -131395 -8354 -131351
rect -8310 -131395 -8254 -131351
rect -8210 -131395 -8154 -131351
rect -8110 -131395 -8054 -131351
rect -8010 -131395 -7954 -131351
rect -7910 -131395 -7854 -131351
rect -7810 -131395 -7354 -131351
rect -7310 -131395 -7254 -131351
rect -7210 -131395 -7154 -131351
rect -7110 -131395 -7054 -131351
rect -7010 -131395 -6954 -131351
rect -6910 -131395 -6854 -131351
rect -6810 -131395 -6754 -131351
rect -6710 -131395 -6654 -131351
rect -6610 -131395 -6554 -131351
rect -6510 -131395 -6454 -131351
rect -6410 -131395 -6354 -131351
rect -6310 -131395 -6254 -131351
rect -6210 -131395 -6154 -131351
rect -6110 -131395 -6054 -131351
rect -6010 -131395 -5954 -131351
rect -5910 -131395 -5854 -131351
rect -5810 -131395 -2893 -131351
rect -16409 -131451 -2893 -131395
rect -16409 -131495 -13354 -131451
rect -13310 -131495 -13254 -131451
rect -13210 -131495 -13154 -131451
rect -13110 -131495 -13054 -131451
rect -13010 -131495 -12954 -131451
rect -12910 -131495 -12854 -131451
rect -12810 -131495 -12754 -131451
rect -12710 -131495 -12654 -131451
rect -12610 -131495 -12554 -131451
rect -12510 -131495 -12454 -131451
rect -12410 -131495 -12354 -131451
rect -12310 -131495 -12254 -131451
rect -12210 -131495 -12154 -131451
rect -12110 -131495 -12054 -131451
rect -12010 -131495 -11954 -131451
rect -11910 -131495 -11854 -131451
rect -11810 -131495 -11354 -131451
rect -11310 -131495 -11254 -131451
rect -11210 -131495 -11154 -131451
rect -11110 -131495 -11054 -131451
rect -11010 -131495 -10954 -131451
rect -10910 -131495 -10854 -131451
rect -10810 -131495 -10754 -131451
rect -10710 -131495 -10654 -131451
rect -10610 -131495 -10554 -131451
rect -10510 -131495 -10454 -131451
rect -10410 -131495 -10354 -131451
rect -10310 -131495 -10254 -131451
rect -10210 -131495 -10154 -131451
rect -10110 -131495 -10054 -131451
rect -10010 -131495 -9954 -131451
rect -9910 -131495 -9854 -131451
rect -9810 -131495 -9354 -131451
rect -9310 -131495 -9254 -131451
rect -9210 -131495 -9154 -131451
rect -9110 -131495 -9054 -131451
rect -9010 -131495 -8954 -131451
rect -8910 -131495 -8854 -131451
rect -8810 -131495 -8754 -131451
rect -8710 -131495 -8654 -131451
rect -8610 -131495 -8554 -131451
rect -8510 -131495 -8454 -131451
rect -8410 -131495 -8354 -131451
rect -8310 -131495 -8254 -131451
rect -8210 -131495 -8154 -131451
rect -8110 -131495 -8054 -131451
rect -8010 -131495 -7954 -131451
rect -7910 -131495 -7854 -131451
rect -7810 -131495 -7354 -131451
rect -7310 -131495 -7254 -131451
rect -7210 -131495 -7154 -131451
rect -7110 -131495 -7054 -131451
rect -7010 -131495 -6954 -131451
rect -6910 -131495 -6854 -131451
rect -6810 -131495 -6754 -131451
rect -6710 -131495 -6654 -131451
rect -6610 -131495 -6554 -131451
rect -6510 -131495 -6454 -131451
rect -6410 -131495 -6354 -131451
rect -6310 -131495 -6254 -131451
rect -6210 -131495 -6154 -131451
rect -6110 -131495 -6054 -131451
rect -6010 -131495 -5954 -131451
rect -5910 -131495 -5854 -131451
rect -5810 -131495 -2893 -131451
rect -16409 -131551 -2893 -131495
rect -16409 -131595 -13354 -131551
rect -13310 -131595 -13254 -131551
rect -13210 -131595 -13154 -131551
rect -13110 -131595 -13054 -131551
rect -13010 -131595 -12954 -131551
rect -12910 -131595 -12854 -131551
rect -12810 -131595 -12754 -131551
rect -12710 -131595 -12654 -131551
rect -12610 -131595 -12554 -131551
rect -12510 -131595 -12454 -131551
rect -12410 -131595 -12354 -131551
rect -12310 -131595 -12254 -131551
rect -12210 -131595 -12154 -131551
rect -12110 -131595 -12054 -131551
rect -12010 -131595 -11954 -131551
rect -11910 -131595 -11854 -131551
rect -11810 -131595 -11354 -131551
rect -11310 -131595 -11254 -131551
rect -11210 -131595 -11154 -131551
rect -11110 -131595 -11054 -131551
rect -11010 -131595 -10954 -131551
rect -10910 -131595 -10854 -131551
rect -10810 -131595 -10754 -131551
rect -10710 -131595 -10654 -131551
rect -10610 -131595 -10554 -131551
rect -10510 -131595 -10454 -131551
rect -10410 -131595 -10354 -131551
rect -10310 -131595 -10254 -131551
rect -10210 -131595 -10154 -131551
rect -10110 -131595 -10054 -131551
rect -10010 -131595 -9954 -131551
rect -9910 -131595 -9854 -131551
rect -9810 -131595 -9354 -131551
rect -9310 -131595 -9254 -131551
rect -9210 -131595 -9154 -131551
rect -9110 -131595 -9054 -131551
rect -9010 -131595 -8954 -131551
rect -8910 -131595 -8854 -131551
rect -8810 -131595 -8754 -131551
rect -8710 -131595 -8654 -131551
rect -8610 -131595 -8554 -131551
rect -8510 -131595 -8454 -131551
rect -8410 -131595 -8354 -131551
rect -8310 -131595 -8254 -131551
rect -8210 -131595 -8154 -131551
rect -8110 -131595 -8054 -131551
rect -8010 -131595 -7954 -131551
rect -7910 -131595 -7854 -131551
rect -7810 -131595 -7354 -131551
rect -7310 -131595 -7254 -131551
rect -7210 -131595 -7154 -131551
rect -7110 -131595 -7054 -131551
rect -7010 -131595 -6954 -131551
rect -6910 -131595 -6854 -131551
rect -6810 -131595 -6754 -131551
rect -6710 -131595 -6654 -131551
rect -6610 -131595 -6554 -131551
rect -6510 -131595 -6454 -131551
rect -6410 -131595 -6354 -131551
rect -6310 -131595 -6254 -131551
rect -6210 -131595 -6154 -131551
rect -6110 -131595 -6054 -131551
rect -6010 -131595 -5954 -131551
rect -5910 -131595 -5854 -131551
rect -5810 -131595 -2893 -131551
rect -16409 -131651 -2893 -131595
rect -16409 -131695 -13354 -131651
rect -13310 -131695 -13254 -131651
rect -13210 -131695 -13154 -131651
rect -13110 -131695 -13054 -131651
rect -13010 -131695 -12954 -131651
rect -12910 -131695 -12854 -131651
rect -12810 -131695 -12754 -131651
rect -12710 -131695 -12654 -131651
rect -12610 -131695 -12554 -131651
rect -12510 -131695 -12454 -131651
rect -12410 -131695 -12354 -131651
rect -12310 -131695 -12254 -131651
rect -12210 -131695 -12154 -131651
rect -12110 -131695 -12054 -131651
rect -12010 -131695 -11954 -131651
rect -11910 -131695 -11854 -131651
rect -11810 -131695 -11354 -131651
rect -11310 -131695 -11254 -131651
rect -11210 -131695 -11154 -131651
rect -11110 -131695 -11054 -131651
rect -11010 -131695 -10954 -131651
rect -10910 -131695 -10854 -131651
rect -10810 -131695 -10754 -131651
rect -10710 -131695 -10654 -131651
rect -10610 -131695 -10554 -131651
rect -10510 -131695 -10454 -131651
rect -10410 -131695 -10354 -131651
rect -10310 -131695 -10254 -131651
rect -10210 -131695 -10154 -131651
rect -10110 -131695 -10054 -131651
rect -10010 -131695 -9954 -131651
rect -9910 -131695 -9854 -131651
rect -9810 -131695 -9354 -131651
rect -9310 -131695 -9254 -131651
rect -9210 -131695 -9154 -131651
rect -9110 -131695 -9054 -131651
rect -9010 -131695 -8954 -131651
rect -8910 -131695 -8854 -131651
rect -8810 -131695 -8754 -131651
rect -8710 -131695 -8654 -131651
rect -8610 -131695 -8554 -131651
rect -8510 -131695 -8454 -131651
rect -8410 -131695 -8354 -131651
rect -8310 -131695 -8254 -131651
rect -8210 -131695 -8154 -131651
rect -8110 -131695 -8054 -131651
rect -8010 -131695 -7954 -131651
rect -7910 -131695 -7854 -131651
rect -7810 -131695 -7354 -131651
rect -7310 -131695 -7254 -131651
rect -7210 -131695 -7154 -131651
rect -7110 -131695 -7054 -131651
rect -7010 -131695 -6954 -131651
rect -6910 -131695 -6854 -131651
rect -6810 -131695 -6754 -131651
rect -6710 -131695 -6654 -131651
rect -6610 -131695 -6554 -131651
rect -6510 -131695 -6454 -131651
rect -6410 -131695 -6354 -131651
rect -6310 -131695 -6254 -131651
rect -6210 -131695 -6154 -131651
rect -6110 -131695 -6054 -131651
rect -6010 -131695 -5954 -131651
rect -5910 -131695 -5854 -131651
rect -5810 -131695 -2893 -131651
rect -16409 -131751 -2893 -131695
rect -16409 -131795 -13354 -131751
rect -13310 -131795 -13254 -131751
rect -13210 -131795 -13154 -131751
rect -13110 -131795 -13054 -131751
rect -13010 -131795 -12954 -131751
rect -12910 -131795 -12854 -131751
rect -12810 -131795 -12754 -131751
rect -12710 -131795 -12654 -131751
rect -12610 -131795 -12554 -131751
rect -12510 -131795 -12454 -131751
rect -12410 -131795 -12354 -131751
rect -12310 -131795 -12254 -131751
rect -12210 -131795 -12154 -131751
rect -12110 -131795 -12054 -131751
rect -12010 -131795 -11954 -131751
rect -11910 -131795 -11854 -131751
rect -11810 -131795 -11354 -131751
rect -11310 -131795 -11254 -131751
rect -11210 -131795 -11154 -131751
rect -11110 -131795 -11054 -131751
rect -11010 -131795 -10954 -131751
rect -10910 -131795 -10854 -131751
rect -10810 -131795 -10754 -131751
rect -10710 -131795 -10654 -131751
rect -10610 -131795 -10554 -131751
rect -10510 -131795 -10454 -131751
rect -10410 -131795 -10354 -131751
rect -10310 -131795 -10254 -131751
rect -10210 -131795 -10154 -131751
rect -10110 -131795 -10054 -131751
rect -10010 -131795 -9954 -131751
rect -9910 -131795 -9854 -131751
rect -9810 -131795 -9354 -131751
rect -9310 -131795 -9254 -131751
rect -9210 -131795 -9154 -131751
rect -9110 -131795 -9054 -131751
rect -9010 -131795 -8954 -131751
rect -8910 -131795 -8854 -131751
rect -8810 -131795 -8754 -131751
rect -8710 -131795 -8654 -131751
rect -8610 -131795 -8554 -131751
rect -8510 -131795 -8454 -131751
rect -8410 -131795 -8354 -131751
rect -8310 -131795 -8254 -131751
rect -8210 -131795 -8154 -131751
rect -8110 -131795 -8054 -131751
rect -8010 -131795 -7954 -131751
rect -7910 -131795 -7854 -131751
rect -7810 -131795 -7354 -131751
rect -7310 -131795 -7254 -131751
rect -7210 -131795 -7154 -131751
rect -7110 -131795 -7054 -131751
rect -7010 -131795 -6954 -131751
rect -6910 -131795 -6854 -131751
rect -6810 -131795 -6754 -131751
rect -6710 -131795 -6654 -131751
rect -6610 -131795 -6554 -131751
rect -6510 -131795 -6454 -131751
rect -6410 -131795 -6354 -131751
rect -6310 -131795 -6254 -131751
rect -6210 -131795 -6154 -131751
rect -6110 -131795 -6054 -131751
rect -6010 -131795 -5954 -131751
rect -5910 -131795 -5854 -131751
rect -5810 -131795 -2893 -131751
rect -16409 -131851 -2893 -131795
rect -16409 -131895 -13354 -131851
rect -13310 -131895 -13254 -131851
rect -13210 -131895 -13154 -131851
rect -13110 -131895 -13054 -131851
rect -13010 -131895 -12954 -131851
rect -12910 -131895 -12854 -131851
rect -12810 -131895 -12754 -131851
rect -12710 -131895 -12654 -131851
rect -12610 -131895 -12554 -131851
rect -12510 -131895 -12454 -131851
rect -12410 -131895 -12354 -131851
rect -12310 -131895 -12254 -131851
rect -12210 -131895 -12154 -131851
rect -12110 -131895 -12054 -131851
rect -12010 -131895 -11954 -131851
rect -11910 -131895 -11854 -131851
rect -11810 -131895 -11354 -131851
rect -11310 -131895 -11254 -131851
rect -11210 -131895 -11154 -131851
rect -11110 -131895 -11054 -131851
rect -11010 -131895 -10954 -131851
rect -10910 -131895 -10854 -131851
rect -10810 -131895 -10754 -131851
rect -10710 -131895 -10654 -131851
rect -10610 -131895 -10554 -131851
rect -10510 -131895 -10454 -131851
rect -10410 -131895 -10354 -131851
rect -10310 -131895 -10254 -131851
rect -10210 -131895 -10154 -131851
rect -10110 -131895 -10054 -131851
rect -10010 -131895 -9954 -131851
rect -9910 -131895 -9854 -131851
rect -9810 -131895 -9354 -131851
rect -9310 -131895 -9254 -131851
rect -9210 -131895 -9154 -131851
rect -9110 -131895 -9054 -131851
rect -9010 -131895 -8954 -131851
rect -8910 -131895 -8854 -131851
rect -8810 -131895 -8754 -131851
rect -8710 -131895 -8654 -131851
rect -8610 -131895 -8554 -131851
rect -8510 -131895 -8454 -131851
rect -8410 -131895 -8354 -131851
rect -8310 -131895 -8254 -131851
rect -8210 -131895 -8154 -131851
rect -8110 -131895 -8054 -131851
rect -8010 -131895 -7954 -131851
rect -7910 -131895 -7854 -131851
rect -7810 -131895 -7354 -131851
rect -7310 -131895 -7254 -131851
rect -7210 -131895 -7154 -131851
rect -7110 -131895 -7054 -131851
rect -7010 -131895 -6954 -131851
rect -6910 -131895 -6854 -131851
rect -6810 -131895 -6754 -131851
rect -6710 -131895 -6654 -131851
rect -6610 -131895 -6554 -131851
rect -6510 -131895 -6454 -131851
rect -6410 -131895 -6354 -131851
rect -6310 -131895 -6254 -131851
rect -6210 -131895 -6154 -131851
rect -6110 -131895 -6054 -131851
rect -6010 -131895 -5954 -131851
rect -5910 -131895 -5854 -131851
rect -5810 -131895 -2893 -131851
rect -16409 -131951 -2893 -131895
rect -16409 -131995 -13354 -131951
rect -13310 -131995 -13254 -131951
rect -13210 -131995 -13154 -131951
rect -13110 -131995 -13054 -131951
rect -13010 -131995 -12954 -131951
rect -12910 -131995 -12854 -131951
rect -12810 -131995 -12754 -131951
rect -12710 -131995 -12654 -131951
rect -12610 -131995 -12554 -131951
rect -12510 -131995 -12454 -131951
rect -12410 -131995 -12354 -131951
rect -12310 -131995 -12254 -131951
rect -12210 -131995 -12154 -131951
rect -12110 -131995 -12054 -131951
rect -12010 -131995 -11954 -131951
rect -11910 -131995 -11854 -131951
rect -11810 -131995 -11354 -131951
rect -11310 -131995 -11254 -131951
rect -11210 -131995 -11154 -131951
rect -11110 -131995 -11054 -131951
rect -11010 -131995 -10954 -131951
rect -10910 -131995 -10854 -131951
rect -10810 -131995 -10754 -131951
rect -10710 -131995 -10654 -131951
rect -10610 -131995 -10554 -131951
rect -10510 -131995 -10454 -131951
rect -10410 -131995 -10354 -131951
rect -10310 -131995 -10254 -131951
rect -10210 -131995 -10154 -131951
rect -10110 -131995 -10054 -131951
rect -10010 -131995 -9954 -131951
rect -9910 -131995 -9854 -131951
rect -9810 -131995 -9354 -131951
rect -9310 -131995 -9254 -131951
rect -9210 -131995 -9154 -131951
rect -9110 -131995 -9054 -131951
rect -9010 -131995 -8954 -131951
rect -8910 -131995 -8854 -131951
rect -8810 -131995 -8754 -131951
rect -8710 -131995 -8654 -131951
rect -8610 -131995 -8554 -131951
rect -8510 -131995 -8454 -131951
rect -8410 -131995 -8354 -131951
rect -8310 -131995 -8254 -131951
rect -8210 -131995 -8154 -131951
rect -8110 -131995 -8054 -131951
rect -8010 -131995 -7954 -131951
rect -7910 -131995 -7854 -131951
rect -7810 -131995 -7354 -131951
rect -7310 -131995 -7254 -131951
rect -7210 -131995 -7154 -131951
rect -7110 -131995 -7054 -131951
rect -7010 -131995 -6954 -131951
rect -6910 -131995 -6854 -131951
rect -6810 -131995 -6754 -131951
rect -6710 -131995 -6654 -131951
rect -6610 -131995 -6554 -131951
rect -6510 -131995 -6454 -131951
rect -6410 -131995 -6354 -131951
rect -6310 -131995 -6254 -131951
rect -6210 -131995 -6154 -131951
rect -6110 -131995 -6054 -131951
rect -6010 -131995 -5954 -131951
rect -5910 -131995 -5854 -131951
rect -5810 -131995 -2893 -131951
rect -16409 -132051 -2893 -131995
rect -16409 -132095 -13354 -132051
rect -13310 -132095 -13254 -132051
rect -13210 -132095 -13154 -132051
rect -13110 -132095 -13054 -132051
rect -13010 -132095 -12954 -132051
rect -12910 -132095 -12854 -132051
rect -12810 -132095 -12754 -132051
rect -12710 -132095 -12654 -132051
rect -12610 -132095 -12554 -132051
rect -12510 -132095 -12454 -132051
rect -12410 -132095 -12354 -132051
rect -12310 -132095 -12254 -132051
rect -12210 -132095 -12154 -132051
rect -12110 -132095 -12054 -132051
rect -12010 -132095 -11954 -132051
rect -11910 -132095 -11854 -132051
rect -11810 -132095 -11354 -132051
rect -11310 -132095 -11254 -132051
rect -11210 -132095 -11154 -132051
rect -11110 -132095 -11054 -132051
rect -11010 -132095 -10954 -132051
rect -10910 -132095 -10854 -132051
rect -10810 -132095 -10754 -132051
rect -10710 -132095 -10654 -132051
rect -10610 -132095 -10554 -132051
rect -10510 -132095 -10454 -132051
rect -10410 -132095 -10354 -132051
rect -10310 -132095 -10254 -132051
rect -10210 -132095 -10154 -132051
rect -10110 -132095 -10054 -132051
rect -10010 -132095 -9954 -132051
rect -9910 -132095 -9854 -132051
rect -9810 -132095 -9354 -132051
rect -9310 -132095 -9254 -132051
rect -9210 -132095 -9154 -132051
rect -9110 -132095 -9054 -132051
rect -9010 -132095 -8954 -132051
rect -8910 -132095 -8854 -132051
rect -8810 -132095 -8754 -132051
rect -8710 -132095 -8654 -132051
rect -8610 -132095 -8554 -132051
rect -8510 -132095 -8454 -132051
rect -8410 -132095 -8354 -132051
rect -8310 -132095 -8254 -132051
rect -8210 -132095 -8154 -132051
rect -8110 -132095 -8054 -132051
rect -8010 -132095 -7954 -132051
rect -7910 -132095 -7854 -132051
rect -7810 -132095 -7354 -132051
rect -7310 -132095 -7254 -132051
rect -7210 -132095 -7154 -132051
rect -7110 -132095 -7054 -132051
rect -7010 -132095 -6954 -132051
rect -6910 -132095 -6854 -132051
rect -6810 -132095 -6754 -132051
rect -6710 -132095 -6654 -132051
rect -6610 -132095 -6554 -132051
rect -6510 -132095 -6454 -132051
rect -6410 -132095 -6354 -132051
rect -6310 -132095 -6254 -132051
rect -6210 -132095 -6154 -132051
rect -6110 -132095 -6054 -132051
rect -6010 -132095 -5954 -132051
rect -5910 -132095 -5854 -132051
rect -5810 -132095 -2893 -132051
rect -16409 -132151 -2893 -132095
rect -16409 -132195 -13354 -132151
rect -13310 -132195 -13254 -132151
rect -13210 -132195 -13154 -132151
rect -13110 -132195 -13054 -132151
rect -13010 -132195 -12954 -132151
rect -12910 -132195 -12854 -132151
rect -12810 -132195 -12754 -132151
rect -12710 -132195 -12654 -132151
rect -12610 -132195 -12554 -132151
rect -12510 -132195 -12454 -132151
rect -12410 -132195 -12354 -132151
rect -12310 -132195 -12254 -132151
rect -12210 -132195 -12154 -132151
rect -12110 -132195 -12054 -132151
rect -12010 -132195 -11954 -132151
rect -11910 -132195 -11854 -132151
rect -11810 -132195 -11354 -132151
rect -11310 -132195 -11254 -132151
rect -11210 -132195 -11154 -132151
rect -11110 -132195 -11054 -132151
rect -11010 -132195 -10954 -132151
rect -10910 -132195 -10854 -132151
rect -10810 -132195 -10754 -132151
rect -10710 -132195 -10654 -132151
rect -10610 -132195 -10554 -132151
rect -10510 -132195 -10454 -132151
rect -10410 -132195 -10354 -132151
rect -10310 -132195 -10254 -132151
rect -10210 -132195 -10154 -132151
rect -10110 -132195 -10054 -132151
rect -10010 -132195 -9954 -132151
rect -9910 -132195 -9854 -132151
rect -9810 -132195 -9354 -132151
rect -9310 -132195 -9254 -132151
rect -9210 -132195 -9154 -132151
rect -9110 -132195 -9054 -132151
rect -9010 -132195 -8954 -132151
rect -8910 -132195 -8854 -132151
rect -8810 -132195 -8754 -132151
rect -8710 -132195 -8654 -132151
rect -8610 -132195 -8554 -132151
rect -8510 -132195 -8454 -132151
rect -8410 -132195 -8354 -132151
rect -8310 -132195 -8254 -132151
rect -8210 -132195 -8154 -132151
rect -8110 -132195 -8054 -132151
rect -8010 -132195 -7954 -132151
rect -7910 -132195 -7854 -132151
rect -7810 -132195 -7354 -132151
rect -7310 -132195 -7254 -132151
rect -7210 -132195 -7154 -132151
rect -7110 -132195 -7054 -132151
rect -7010 -132195 -6954 -132151
rect -6910 -132195 -6854 -132151
rect -6810 -132195 -6754 -132151
rect -6710 -132195 -6654 -132151
rect -6610 -132195 -6554 -132151
rect -6510 -132195 -6454 -132151
rect -6410 -132195 -6354 -132151
rect -6310 -132195 -6254 -132151
rect -6210 -132195 -6154 -132151
rect -6110 -132195 -6054 -132151
rect -6010 -132195 -5954 -132151
rect -5910 -132195 -5854 -132151
rect -5810 -132195 -2893 -132151
rect -16409 -132251 -2893 -132195
rect -16409 -132295 -13354 -132251
rect -13310 -132295 -13254 -132251
rect -13210 -132295 -13154 -132251
rect -13110 -132295 -13054 -132251
rect -13010 -132295 -12954 -132251
rect -12910 -132295 -12854 -132251
rect -12810 -132295 -12754 -132251
rect -12710 -132295 -12654 -132251
rect -12610 -132295 -12554 -132251
rect -12510 -132295 -12454 -132251
rect -12410 -132295 -12354 -132251
rect -12310 -132295 -12254 -132251
rect -12210 -132295 -12154 -132251
rect -12110 -132295 -12054 -132251
rect -12010 -132295 -11954 -132251
rect -11910 -132295 -11854 -132251
rect -11810 -132295 -11354 -132251
rect -11310 -132295 -11254 -132251
rect -11210 -132295 -11154 -132251
rect -11110 -132295 -11054 -132251
rect -11010 -132295 -10954 -132251
rect -10910 -132295 -10854 -132251
rect -10810 -132295 -10754 -132251
rect -10710 -132295 -10654 -132251
rect -10610 -132295 -10554 -132251
rect -10510 -132295 -10454 -132251
rect -10410 -132295 -10354 -132251
rect -10310 -132295 -10254 -132251
rect -10210 -132295 -10154 -132251
rect -10110 -132295 -10054 -132251
rect -10010 -132295 -9954 -132251
rect -9910 -132295 -9854 -132251
rect -9810 -132295 -9354 -132251
rect -9310 -132295 -9254 -132251
rect -9210 -132295 -9154 -132251
rect -9110 -132295 -9054 -132251
rect -9010 -132295 -8954 -132251
rect -8910 -132295 -8854 -132251
rect -8810 -132295 -8754 -132251
rect -8710 -132295 -8654 -132251
rect -8610 -132295 -8554 -132251
rect -8510 -132295 -8454 -132251
rect -8410 -132295 -8354 -132251
rect -8310 -132295 -8254 -132251
rect -8210 -132295 -8154 -132251
rect -8110 -132295 -8054 -132251
rect -8010 -132295 -7954 -132251
rect -7910 -132295 -7854 -132251
rect -7810 -132295 -7354 -132251
rect -7310 -132295 -7254 -132251
rect -7210 -132295 -7154 -132251
rect -7110 -132295 -7054 -132251
rect -7010 -132295 -6954 -132251
rect -6910 -132295 -6854 -132251
rect -6810 -132295 -6754 -132251
rect -6710 -132295 -6654 -132251
rect -6610 -132295 -6554 -132251
rect -6510 -132295 -6454 -132251
rect -6410 -132295 -6354 -132251
rect -6310 -132295 -6254 -132251
rect -6210 -132295 -6154 -132251
rect -6110 -132295 -6054 -132251
rect -6010 -132295 -5954 -132251
rect -5910 -132295 -5854 -132251
rect -5810 -132295 -2893 -132251
rect -16409 -132351 -2893 -132295
rect -16409 -132395 -13354 -132351
rect -13310 -132395 -13254 -132351
rect -13210 -132395 -13154 -132351
rect -13110 -132395 -13054 -132351
rect -13010 -132395 -12954 -132351
rect -12910 -132395 -12854 -132351
rect -12810 -132395 -12754 -132351
rect -12710 -132395 -12654 -132351
rect -12610 -132395 -12554 -132351
rect -12510 -132395 -12454 -132351
rect -12410 -132395 -12354 -132351
rect -12310 -132395 -12254 -132351
rect -12210 -132395 -12154 -132351
rect -12110 -132395 -12054 -132351
rect -12010 -132395 -11954 -132351
rect -11910 -132395 -11854 -132351
rect -11810 -132395 -11354 -132351
rect -11310 -132395 -11254 -132351
rect -11210 -132395 -11154 -132351
rect -11110 -132395 -11054 -132351
rect -11010 -132395 -10954 -132351
rect -10910 -132395 -10854 -132351
rect -10810 -132395 -10754 -132351
rect -10710 -132395 -10654 -132351
rect -10610 -132395 -10554 -132351
rect -10510 -132395 -10454 -132351
rect -10410 -132395 -10354 -132351
rect -10310 -132395 -10254 -132351
rect -10210 -132395 -10154 -132351
rect -10110 -132395 -10054 -132351
rect -10010 -132395 -9954 -132351
rect -9910 -132395 -9854 -132351
rect -9810 -132395 -9354 -132351
rect -9310 -132395 -9254 -132351
rect -9210 -132395 -9154 -132351
rect -9110 -132395 -9054 -132351
rect -9010 -132395 -8954 -132351
rect -8910 -132395 -8854 -132351
rect -8810 -132395 -8754 -132351
rect -8710 -132395 -8654 -132351
rect -8610 -132395 -8554 -132351
rect -8510 -132395 -8454 -132351
rect -8410 -132395 -8354 -132351
rect -8310 -132395 -8254 -132351
rect -8210 -132395 -8154 -132351
rect -8110 -132395 -8054 -132351
rect -8010 -132395 -7954 -132351
rect -7910 -132395 -7854 -132351
rect -7810 -132395 -7354 -132351
rect -7310 -132395 -7254 -132351
rect -7210 -132395 -7154 -132351
rect -7110 -132395 -7054 -132351
rect -7010 -132395 -6954 -132351
rect -6910 -132395 -6854 -132351
rect -6810 -132395 -6754 -132351
rect -6710 -132395 -6654 -132351
rect -6610 -132395 -6554 -132351
rect -6510 -132395 -6454 -132351
rect -6410 -132395 -6354 -132351
rect -6310 -132395 -6254 -132351
rect -6210 -132395 -6154 -132351
rect -6110 -132395 -6054 -132351
rect -6010 -132395 -5954 -132351
rect -5910 -132395 -5854 -132351
rect -5810 -132395 -2893 -132351
rect -16409 -132451 -2893 -132395
rect -16409 -132495 -13354 -132451
rect -13310 -132495 -13254 -132451
rect -13210 -132495 -13154 -132451
rect -13110 -132495 -13054 -132451
rect -13010 -132495 -12954 -132451
rect -12910 -132495 -12854 -132451
rect -12810 -132495 -12754 -132451
rect -12710 -132495 -12654 -132451
rect -12610 -132495 -12554 -132451
rect -12510 -132495 -12454 -132451
rect -12410 -132495 -12354 -132451
rect -12310 -132495 -12254 -132451
rect -12210 -132495 -12154 -132451
rect -12110 -132495 -12054 -132451
rect -12010 -132495 -11954 -132451
rect -11910 -132495 -11854 -132451
rect -11810 -132495 -11354 -132451
rect -11310 -132495 -11254 -132451
rect -11210 -132495 -11154 -132451
rect -11110 -132495 -11054 -132451
rect -11010 -132495 -10954 -132451
rect -10910 -132495 -10854 -132451
rect -10810 -132495 -10754 -132451
rect -10710 -132495 -10654 -132451
rect -10610 -132495 -10554 -132451
rect -10510 -132495 -10454 -132451
rect -10410 -132495 -10354 -132451
rect -10310 -132495 -10254 -132451
rect -10210 -132495 -10154 -132451
rect -10110 -132495 -10054 -132451
rect -10010 -132495 -9954 -132451
rect -9910 -132495 -9854 -132451
rect -9810 -132495 -9354 -132451
rect -9310 -132495 -9254 -132451
rect -9210 -132495 -9154 -132451
rect -9110 -132495 -9054 -132451
rect -9010 -132495 -8954 -132451
rect -8910 -132495 -8854 -132451
rect -8810 -132495 -8754 -132451
rect -8710 -132495 -8654 -132451
rect -8610 -132495 -8554 -132451
rect -8510 -132495 -8454 -132451
rect -8410 -132495 -8354 -132451
rect -8310 -132495 -8254 -132451
rect -8210 -132495 -8154 -132451
rect -8110 -132495 -8054 -132451
rect -8010 -132495 -7954 -132451
rect -7910 -132495 -7854 -132451
rect -7810 -132495 -7354 -132451
rect -7310 -132495 -7254 -132451
rect -7210 -132495 -7154 -132451
rect -7110 -132495 -7054 -132451
rect -7010 -132495 -6954 -132451
rect -6910 -132495 -6854 -132451
rect -6810 -132495 -6754 -132451
rect -6710 -132495 -6654 -132451
rect -6610 -132495 -6554 -132451
rect -6510 -132495 -6454 -132451
rect -6410 -132495 -6354 -132451
rect -6310 -132495 -6254 -132451
rect -6210 -132495 -6154 -132451
rect -6110 -132495 -6054 -132451
rect -6010 -132495 -5954 -132451
rect -5910 -132495 -5854 -132451
rect -5810 -132495 -2893 -132451
rect -16409 -132551 -2893 -132495
rect -16409 -132595 -13354 -132551
rect -13310 -132595 -13254 -132551
rect -13210 -132595 -13154 -132551
rect -13110 -132595 -13054 -132551
rect -13010 -132595 -12954 -132551
rect -12910 -132595 -12854 -132551
rect -12810 -132595 -12754 -132551
rect -12710 -132595 -12654 -132551
rect -12610 -132595 -12554 -132551
rect -12510 -132595 -12454 -132551
rect -12410 -132595 -12354 -132551
rect -12310 -132595 -12254 -132551
rect -12210 -132595 -12154 -132551
rect -12110 -132595 -12054 -132551
rect -12010 -132595 -11954 -132551
rect -11910 -132595 -11854 -132551
rect -11810 -132595 -11354 -132551
rect -11310 -132595 -11254 -132551
rect -11210 -132595 -11154 -132551
rect -11110 -132595 -11054 -132551
rect -11010 -132595 -10954 -132551
rect -10910 -132595 -10854 -132551
rect -10810 -132595 -10754 -132551
rect -10710 -132595 -10654 -132551
rect -10610 -132595 -10554 -132551
rect -10510 -132595 -10454 -132551
rect -10410 -132595 -10354 -132551
rect -10310 -132595 -10254 -132551
rect -10210 -132595 -10154 -132551
rect -10110 -132595 -10054 -132551
rect -10010 -132595 -9954 -132551
rect -9910 -132595 -9854 -132551
rect -9810 -132595 -9354 -132551
rect -9310 -132595 -9254 -132551
rect -9210 -132595 -9154 -132551
rect -9110 -132595 -9054 -132551
rect -9010 -132595 -8954 -132551
rect -8910 -132595 -8854 -132551
rect -8810 -132595 -8754 -132551
rect -8710 -132595 -8654 -132551
rect -8610 -132595 -8554 -132551
rect -8510 -132595 -8454 -132551
rect -8410 -132595 -8354 -132551
rect -8310 -132595 -8254 -132551
rect -8210 -132595 -8154 -132551
rect -8110 -132595 -8054 -132551
rect -8010 -132595 -7954 -132551
rect -7910 -132595 -7854 -132551
rect -7810 -132595 -7354 -132551
rect -7310 -132595 -7254 -132551
rect -7210 -132595 -7154 -132551
rect -7110 -132595 -7054 -132551
rect -7010 -132595 -6954 -132551
rect -6910 -132595 -6854 -132551
rect -6810 -132595 -6754 -132551
rect -6710 -132595 -6654 -132551
rect -6610 -132595 -6554 -132551
rect -6510 -132595 -6454 -132551
rect -6410 -132595 -6354 -132551
rect -6310 -132595 -6254 -132551
rect -6210 -132595 -6154 -132551
rect -6110 -132595 -6054 -132551
rect -6010 -132595 -5954 -132551
rect -5910 -132595 -5854 -132551
rect -5810 -132595 -2893 -132551
rect -16409 -132651 -2893 -132595
rect -16409 -132695 -13354 -132651
rect -13310 -132695 -13254 -132651
rect -13210 -132695 -13154 -132651
rect -13110 -132695 -13054 -132651
rect -13010 -132695 -12954 -132651
rect -12910 -132695 -12854 -132651
rect -12810 -132695 -12754 -132651
rect -12710 -132695 -12654 -132651
rect -12610 -132695 -12554 -132651
rect -12510 -132695 -12454 -132651
rect -12410 -132695 -12354 -132651
rect -12310 -132695 -12254 -132651
rect -12210 -132695 -12154 -132651
rect -12110 -132695 -12054 -132651
rect -12010 -132695 -11954 -132651
rect -11910 -132695 -11854 -132651
rect -11810 -132695 -11354 -132651
rect -11310 -132695 -11254 -132651
rect -11210 -132695 -11154 -132651
rect -11110 -132695 -11054 -132651
rect -11010 -132695 -10954 -132651
rect -10910 -132695 -10854 -132651
rect -10810 -132695 -10754 -132651
rect -10710 -132695 -10654 -132651
rect -10610 -132695 -10554 -132651
rect -10510 -132695 -10454 -132651
rect -10410 -132695 -10354 -132651
rect -10310 -132695 -10254 -132651
rect -10210 -132695 -10154 -132651
rect -10110 -132695 -10054 -132651
rect -10010 -132695 -9954 -132651
rect -9910 -132695 -9854 -132651
rect -9810 -132695 -9354 -132651
rect -9310 -132695 -9254 -132651
rect -9210 -132695 -9154 -132651
rect -9110 -132695 -9054 -132651
rect -9010 -132695 -8954 -132651
rect -8910 -132695 -8854 -132651
rect -8810 -132695 -8754 -132651
rect -8710 -132695 -8654 -132651
rect -8610 -132695 -8554 -132651
rect -8510 -132695 -8454 -132651
rect -8410 -132695 -8354 -132651
rect -8310 -132695 -8254 -132651
rect -8210 -132695 -8154 -132651
rect -8110 -132695 -8054 -132651
rect -8010 -132695 -7954 -132651
rect -7910 -132695 -7854 -132651
rect -7810 -132695 -7354 -132651
rect -7310 -132695 -7254 -132651
rect -7210 -132695 -7154 -132651
rect -7110 -132695 -7054 -132651
rect -7010 -132695 -6954 -132651
rect -6910 -132695 -6854 -132651
rect -6810 -132695 -6754 -132651
rect -6710 -132695 -6654 -132651
rect -6610 -132695 -6554 -132651
rect -6510 -132695 -6454 -132651
rect -6410 -132695 -6354 -132651
rect -6310 -132695 -6254 -132651
rect -6210 -132695 -6154 -132651
rect -6110 -132695 -6054 -132651
rect -6010 -132695 -5954 -132651
rect -5910 -132695 -5854 -132651
rect -5810 -132695 -2893 -132651
rect -16409 -132751 -2893 -132695
rect -16409 -132795 -13354 -132751
rect -13310 -132795 -13254 -132751
rect -13210 -132795 -13154 -132751
rect -13110 -132795 -13054 -132751
rect -13010 -132795 -12954 -132751
rect -12910 -132795 -12854 -132751
rect -12810 -132795 -12754 -132751
rect -12710 -132795 -12654 -132751
rect -12610 -132795 -12554 -132751
rect -12510 -132795 -12454 -132751
rect -12410 -132795 -12354 -132751
rect -12310 -132795 -12254 -132751
rect -12210 -132795 -12154 -132751
rect -12110 -132795 -12054 -132751
rect -12010 -132795 -11954 -132751
rect -11910 -132795 -11854 -132751
rect -11810 -132795 -11354 -132751
rect -11310 -132795 -11254 -132751
rect -11210 -132795 -11154 -132751
rect -11110 -132795 -11054 -132751
rect -11010 -132795 -10954 -132751
rect -10910 -132795 -10854 -132751
rect -10810 -132795 -10754 -132751
rect -10710 -132795 -10654 -132751
rect -10610 -132795 -10554 -132751
rect -10510 -132795 -10454 -132751
rect -10410 -132795 -10354 -132751
rect -10310 -132795 -10254 -132751
rect -10210 -132795 -10154 -132751
rect -10110 -132795 -10054 -132751
rect -10010 -132795 -9954 -132751
rect -9910 -132795 -9854 -132751
rect -9810 -132795 -9354 -132751
rect -9310 -132795 -9254 -132751
rect -9210 -132795 -9154 -132751
rect -9110 -132795 -9054 -132751
rect -9010 -132795 -8954 -132751
rect -8910 -132795 -8854 -132751
rect -8810 -132795 -8754 -132751
rect -8710 -132795 -8654 -132751
rect -8610 -132795 -8554 -132751
rect -8510 -132795 -8454 -132751
rect -8410 -132795 -8354 -132751
rect -8310 -132795 -8254 -132751
rect -8210 -132795 -8154 -132751
rect -8110 -132795 -8054 -132751
rect -8010 -132795 -7954 -132751
rect -7910 -132795 -7854 -132751
rect -7810 -132795 -7354 -132751
rect -7310 -132795 -7254 -132751
rect -7210 -132795 -7154 -132751
rect -7110 -132795 -7054 -132751
rect -7010 -132795 -6954 -132751
rect -6910 -132795 -6854 -132751
rect -6810 -132795 -6754 -132751
rect -6710 -132795 -6654 -132751
rect -6610 -132795 -6554 -132751
rect -6510 -132795 -6454 -132751
rect -6410 -132795 -6354 -132751
rect -6310 -132795 -6254 -132751
rect -6210 -132795 -6154 -132751
rect -6110 -132795 -6054 -132751
rect -6010 -132795 -5954 -132751
rect -5910 -132795 -5854 -132751
rect -5810 -132795 -2893 -132751
rect -16409 -133867 -2893 -132795
rect 34207 -131385 47953 -11182
rect 178461 -11978 181332 9144
rect 173132 -13446 181332 -11978
rect 188605 6863 192404 6987
rect 188605 6200 190005 6863
rect 191144 6200 192404 6863
rect 142660 -17445 154949 -15886
rect 142660 -17489 144904 -17445
rect 144948 -17489 145004 -17445
rect 145048 -17489 145104 -17445
rect 145148 -17489 145204 -17445
rect 145248 -17489 145304 -17445
rect 145348 -17489 145404 -17445
rect 145448 -17489 145504 -17445
rect 145548 -17489 145604 -17445
rect 145648 -17489 145704 -17445
rect 145748 -17489 145804 -17445
rect 145848 -17489 145904 -17445
rect 145948 -17489 146004 -17445
rect 146048 -17489 146104 -17445
rect 146148 -17489 146204 -17445
rect 146248 -17489 146304 -17445
rect 146348 -17489 146404 -17445
rect 146448 -17489 146904 -17445
rect 146948 -17489 147004 -17445
rect 147048 -17489 147104 -17445
rect 147148 -17489 147204 -17445
rect 147248 -17489 147304 -17445
rect 147348 -17489 147404 -17445
rect 147448 -17489 147504 -17445
rect 147548 -17489 147604 -17445
rect 147648 -17489 147704 -17445
rect 147748 -17489 147804 -17445
rect 147848 -17489 147904 -17445
rect 147948 -17489 148004 -17445
rect 148048 -17489 148104 -17445
rect 148148 -17489 148204 -17445
rect 148248 -17489 148304 -17445
rect 148348 -17489 148404 -17445
rect 148448 -17489 148904 -17445
rect 148948 -17489 149004 -17445
rect 149048 -17489 149104 -17445
rect 149148 -17489 149204 -17445
rect 149248 -17489 149304 -17445
rect 149348 -17489 149404 -17445
rect 149448 -17489 149504 -17445
rect 149548 -17489 149604 -17445
rect 149648 -17489 149704 -17445
rect 149748 -17489 149804 -17445
rect 149848 -17489 149904 -17445
rect 149948 -17489 150004 -17445
rect 150048 -17489 150104 -17445
rect 150148 -17489 150204 -17445
rect 150248 -17489 150304 -17445
rect 150348 -17489 150404 -17445
rect 150448 -17489 150904 -17445
rect 150948 -17489 151004 -17445
rect 151048 -17489 151104 -17445
rect 151148 -17489 151204 -17445
rect 151248 -17489 151304 -17445
rect 151348 -17489 151404 -17445
rect 151448 -17489 151504 -17445
rect 151548 -17489 151604 -17445
rect 151648 -17489 151704 -17445
rect 151748 -17489 151804 -17445
rect 151848 -17489 151904 -17445
rect 151948 -17489 152004 -17445
rect 152048 -17489 152104 -17445
rect 152148 -17489 152204 -17445
rect 152248 -17489 152304 -17445
rect 152348 -17489 152404 -17445
rect 152448 -17489 154949 -17445
rect 142660 -17545 154949 -17489
rect 142660 -17589 144904 -17545
rect 144948 -17589 145004 -17545
rect 145048 -17589 145104 -17545
rect 145148 -17589 145204 -17545
rect 145248 -17589 145304 -17545
rect 145348 -17589 145404 -17545
rect 145448 -17589 145504 -17545
rect 145548 -17589 145604 -17545
rect 145648 -17589 145704 -17545
rect 145748 -17589 145804 -17545
rect 145848 -17589 145904 -17545
rect 145948 -17589 146004 -17545
rect 146048 -17589 146104 -17545
rect 146148 -17589 146204 -17545
rect 146248 -17589 146304 -17545
rect 146348 -17589 146404 -17545
rect 146448 -17589 146904 -17545
rect 146948 -17589 147004 -17545
rect 147048 -17589 147104 -17545
rect 147148 -17589 147204 -17545
rect 147248 -17589 147304 -17545
rect 147348 -17589 147404 -17545
rect 147448 -17589 147504 -17545
rect 147548 -17589 147604 -17545
rect 147648 -17589 147704 -17545
rect 147748 -17589 147804 -17545
rect 147848 -17589 147904 -17545
rect 147948 -17589 148004 -17545
rect 148048 -17589 148104 -17545
rect 148148 -17589 148204 -17545
rect 148248 -17589 148304 -17545
rect 148348 -17589 148404 -17545
rect 148448 -17589 148904 -17545
rect 148948 -17589 149004 -17545
rect 149048 -17589 149104 -17545
rect 149148 -17589 149204 -17545
rect 149248 -17589 149304 -17545
rect 149348 -17589 149404 -17545
rect 149448 -17589 149504 -17545
rect 149548 -17589 149604 -17545
rect 149648 -17589 149704 -17545
rect 149748 -17589 149804 -17545
rect 149848 -17589 149904 -17545
rect 149948 -17589 150004 -17545
rect 150048 -17589 150104 -17545
rect 150148 -17589 150204 -17545
rect 150248 -17589 150304 -17545
rect 150348 -17589 150404 -17545
rect 150448 -17589 150904 -17545
rect 150948 -17589 151004 -17545
rect 151048 -17589 151104 -17545
rect 151148 -17589 151204 -17545
rect 151248 -17589 151304 -17545
rect 151348 -17589 151404 -17545
rect 151448 -17589 151504 -17545
rect 151548 -17589 151604 -17545
rect 151648 -17589 151704 -17545
rect 151748 -17589 151804 -17545
rect 151848 -17589 151904 -17545
rect 151948 -17589 152004 -17545
rect 152048 -17589 152104 -17545
rect 152148 -17589 152204 -17545
rect 152248 -17589 152304 -17545
rect 152348 -17589 152404 -17545
rect 152448 -17589 154949 -17545
rect 142660 -17645 154949 -17589
rect 142660 -17689 144904 -17645
rect 144948 -17689 145004 -17645
rect 145048 -17689 145104 -17645
rect 145148 -17689 145204 -17645
rect 145248 -17689 145304 -17645
rect 145348 -17689 145404 -17645
rect 145448 -17689 145504 -17645
rect 145548 -17689 145604 -17645
rect 145648 -17689 145704 -17645
rect 145748 -17689 145804 -17645
rect 145848 -17689 145904 -17645
rect 145948 -17689 146004 -17645
rect 146048 -17689 146104 -17645
rect 146148 -17689 146204 -17645
rect 146248 -17689 146304 -17645
rect 146348 -17689 146404 -17645
rect 146448 -17689 146904 -17645
rect 146948 -17689 147004 -17645
rect 147048 -17689 147104 -17645
rect 147148 -17689 147204 -17645
rect 147248 -17689 147304 -17645
rect 147348 -17689 147404 -17645
rect 147448 -17689 147504 -17645
rect 147548 -17689 147604 -17645
rect 147648 -17689 147704 -17645
rect 147748 -17689 147804 -17645
rect 147848 -17689 147904 -17645
rect 147948 -17689 148004 -17645
rect 148048 -17689 148104 -17645
rect 148148 -17689 148204 -17645
rect 148248 -17689 148304 -17645
rect 148348 -17689 148404 -17645
rect 148448 -17689 148904 -17645
rect 148948 -17689 149004 -17645
rect 149048 -17689 149104 -17645
rect 149148 -17689 149204 -17645
rect 149248 -17689 149304 -17645
rect 149348 -17689 149404 -17645
rect 149448 -17689 149504 -17645
rect 149548 -17689 149604 -17645
rect 149648 -17689 149704 -17645
rect 149748 -17689 149804 -17645
rect 149848 -17689 149904 -17645
rect 149948 -17689 150004 -17645
rect 150048 -17689 150104 -17645
rect 150148 -17689 150204 -17645
rect 150248 -17689 150304 -17645
rect 150348 -17689 150404 -17645
rect 150448 -17689 150904 -17645
rect 150948 -17689 151004 -17645
rect 151048 -17689 151104 -17645
rect 151148 -17689 151204 -17645
rect 151248 -17689 151304 -17645
rect 151348 -17689 151404 -17645
rect 151448 -17689 151504 -17645
rect 151548 -17689 151604 -17645
rect 151648 -17689 151704 -17645
rect 151748 -17689 151804 -17645
rect 151848 -17689 151904 -17645
rect 151948 -17689 152004 -17645
rect 152048 -17689 152104 -17645
rect 152148 -17689 152204 -17645
rect 152248 -17689 152304 -17645
rect 152348 -17689 152404 -17645
rect 152448 -17689 154949 -17645
rect 142660 -17745 154949 -17689
rect 142660 -17789 144904 -17745
rect 144948 -17789 145004 -17745
rect 145048 -17789 145104 -17745
rect 145148 -17789 145204 -17745
rect 145248 -17789 145304 -17745
rect 145348 -17789 145404 -17745
rect 145448 -17789 145504 -17745
rect 145548 -17789 145604 -17745
rect 145648 -17789 145704 -17745
rect 145748 -17789 145804 -17745
rect 145848 -17789 145904 -17745
rect 145948 -17789 146004 -17745
rect 146048 -17789 146104 -17745
rect 146148 -17789 146204 -17745
rect 146248 -17789 146304 -17745
rect 146348 -17789 146404 -17745
rect 146448 -17789 146904 -17745
rect 146948 -17789 147004 -17745
rect 147048 -17789 147104 -17745
rect 147148 -17789 147204 -17745
rect 147248 -17789 147304 -17745
rect 147348 -17789 147404 -17745
rect 147448 -17789 147504 -17745
rect 147548 -17789 147604 -17745
rect 147648 -17789 147704 -17745
rect 147748 -17789 147804 -17745
rect 147848 -17789 147904 -17745
rect 147948 -17789 148004 -17745
rect 148048 -17789 148104 -17745
rect 148148 -17789 148204 -17745
rect 148248 -17789 148304 -17745
rect 148348 -17789 148404 -17745
rect 148448 -17789 148904 -17745
rect 148948 -17789 149004 -17745
rect 149048 -17789 149104 -17745
rect 149148 -17789 149204 -17745
rect 149248 -17789 149304 -17745
rect 149348 -17789 149404 -17745
rect 149448 -17789 149504 -17745
rect 149548 -17789 149604 -17745
rect 149648 -17789 149704 -17745
rect 149748 -17789 149804 -17745
rect 149848 -17789 149904 -17745
rect 149948 -17789 150004 -17745
rect 150048 -17789 150104 -17745
rect 150148 -17789 150204 -17745
rect 150248 -17789 150304 -17745
rect 150348 -17789 150404 -17745
rect 150448 -17789 150904 -17745
rect 150948 -17789 151004 -17745
rect 151048 -17789 151104 -17745
rect 151148 -17789 151204 -17745
rect 151248 -17789 151304 -17745
rect 151348 -17789 151404 -17745
rect 151448 -17789 151504 -17745
rect 151548 -17789 151604 -17745
rect 151648 -17789 151704 -17745
rect 151748 -17789 151804 -17745
rect 151848 -17789 151904 -17745
rect 151948 -17789 152004 -17745
rect 152048 -17789 152104 -17745
rect 152148 -17789 152204 -17745
rect 152248 -17789 152304 -17745
rect 152348 -17789 152404 -17745
rect 152448 -17789 154949 -17745
rect 142660 -17845 154949 -17789
rect 142660 -17889 144904 -17845
rect 144948 -17889 145004 -17845
rect 145048 -17889 145104 -17845
rect 145148 -17889 145204 -17845
rect 145248 -17889 145304 -17845
rect 145348 -17889 145404 -17845
rect 145448 -17889 145504 -17845
rect 145548 -17889 145604 -17845
rect 145648 -17889 145704 -17845
rect 145748 -17889 145804 -17845
rect 145848 -17889 145904 -17845
rect 145948 -17889 146004 -17845
rect 146048 -17889 146104 -17845
rect 146148 -17889 146204 -17845
rect 146248 -17889 146304 -17845
rect 146348 -17889 146404 -17845
rect 146448 -17889 146904 -17845
rect 146948 -17889 147004 -17845
rect 147048 -17889 147104 -17845
rect 147148 -17889 147204 -17845
rect 147248 -17889 147304 -17845
rect 147348 -17889 147404 -17845
rect 147448 -17889 147504 -17845
rect 147548 -17889 147604 -17845
rect 147648 -17889 147704 -17845
rect 147748 -17889 147804 -17845
rect 147848 -17889 147904 -17845
rect 147948 -17889 148004 -17845
rect 148048 -17889 148104 -17845
rect 148148 -17889 148204 -17845
rect 148248 -17889 148304 -17845
rect 148348 -17889 148404 -17845
rect 148448 -17889 148904 -17845
rect 148948 -17889 149004 -17845
rect 149048 -17889 149104 -17845
rect 149148 -17889 149204 -17845
rect 149248 -17889 149304 -17845
rect 149348 -17889 149404 -17845
rect 149448 -17889 149504 -17845
rect 149548 -17889 149604 -17845
rect 149648 -17889 149704 -17845
rect 149748 -17889 149804 -17845
rect 149848 -17889 149904 -17845
rect 149948 -17889 150004 -17845
rect 150048 -17889 150104 -17845
rect 150148 -17889 150204 -17845
rect 150248 -17889 150304 -17845
rect 150348 -17889 150404 -17845
rect 150448 -17889 150904 -17845
rect 150948 -17889 151004 -17845
rect 151048 -17889 151104 -17845
rect 151148 -17889 151204 -17845
rect 151248 -17889 151304 -17845
rect 151348 -17889 151404 -17845
rect 151448 -17889 151504 -17845
rect 151548 -17889 151604 -17845
rect 151648 -17889 151704 -17845
rect 151748 -17889 151804 -17845
rect 151848 -17889 151904 -17845
rect 151948 -17889 152004 -17845
rect 152048 -17889 152104 -17845
rect 152148 -17889 152204 -17845
rect 152248 -17889 152304 -17845
rect 152348 -17889 152404 -17845
rect 152448 -17889 154949 -17845
rect 142660 -17945 154949 -17889
rect 142660 -17989 144904 -17945
rect 144948 -17989 145004 -17945
rect 145048 -17989 145104 -17945
rect 145148 -17989 145204 -17945
rect 145248 -17989 145304 -17945
rect 145348 -17989 145404 -17945
rect 145448 -17989 145504 -17945
rect 145548 -17989 145604 -17945
rect 145648 -17989 145704 -17945
rect 145748 -17989 145804 -17945
rect 145848 -17989 145904 -17945
rect 145948 -17989 146004 -17945
rect 146048 -17989 146104 -17945
rect 146148 -17989 146204 -17945
rect 146248 -17989 146304 -17945
rect 146348 -17989 146404 -17945
rect 146448 -17989 146904 -17945
rect 146948 -17989 147004 -17945
rect 147048 -17989 147104 -17945
rect 147148 -17989 147204 -17945
rect 147248 -17989 147304 -17945
rect 147348 -17989 147404 -17945
rect 147448 -17989 147504 -17945
rect 147548 -17989 147604 -17945
rect 147648 -17989 147704 -17945
rect 147748 -17989 147804 -17945
rect 147848 -17989 147904 -17945
rect 147948 -17989 148004 -17945
rect 148048 -17989 148104 -17945
rect 148148 -17989 148204 -17945
rect 148248 -17989 148304 -17945
rect 148348 -17989 148404 -17945
rect 148448 -17989 148904 -17945
rect 148948 -17989 149004 -17945
rect 149048 -17989 149104 -17945
rect 149148 -17989 149204 -17945
rect 149248 -17989 149304 -17945
rect 149348 -17989 149404 -17945
rect 149448 -17989 149504 -17945
rect 149548 -17989 149604 -17945
rect 149648 -17989 149704 -17945
rect 149748 -17989 149804 -17945
rect 149848 -17989 149904 -17945
rect 149948 -17989 150004 -17945
rect 150048 -17989 150104 -17945
rect 150148 -17989 150204 -17945
rect 150248 -17989 150304 -17945
rect 150348 -17989 150404 -17945
rect 150448 -17989 150904 -17945
rect 150948 -17989 151004 -17945
rect 151048 -17989 151104 -17945
rect 151148 -17989 151204 -17945
rect 151248 -17989 151304 -17945
rect 151348 -17989 151404 -17945
rect 151448 -17989 151504 -17945
rect 151548 -17989 151604 -17945
rect 151648 -17989 151704 -17945
rect 151748 -17989 151804 -17945
rect 151848 -17989 151904 -17945
rect 151948 -17989 152004 -17945
rect 152048 -17989 152104 -17945
rect 152148 -17989 152204 -17945
rect 152248 -17989 152304 -17945
rect 152348 -17989 152404 -17945
rect 152448 -17989 154949 -17945
rect 142660 -18045 154949 -17989
rect 142660 -18089 144904 -18045
rect 144948 -18089 145004 -18045
rect 145048 -18089 145104 -18045
rect 145148 -18089 145204 -18045
rect 145248 -18089 145304 -18045
rect 145348 -18089 145404 -18045
rect 145448 -18089 145504 -18045
rect 145548 -18089 145604 -18045
rect 145648 -18089 145704 -18045
rect 145748 -18089 145804 -18045
rect 145848 -18089 145904 -18045
rect 145948 -18089 146004 -18045
rect 146048 -18089 146104 -18045
rect 146148 -18089 146204 -18045
rect 146248 -18089 146304 -18045
rect 146348 -18089 146404 -18045
rect 146448 -18089 146904 -18045
rect 146948 -18089 147004 -18045
rect 147048 -18089 147104 -18045
rect 147148 -18089 147204 -18045
rect 147248 -18089 147304 -18045
rect 147348 -18089 147404 -18045
rect 147448 -18089 147504 -18045
rect 147548 -18089 147604 -18045
rect 147648 -18089 147704 -18045
rect 147748 -18089 147804 -18045
rect 147848 -18089 147904 -18045
rect 147948 -18089 148004 -18045
rect 148048 -18089 148104 -18045
rect 148148 -18089 148204 -18045
rect 148248 -18089 148304 -18045
rect 148348 -18089 148404 -18045
rect 148448 -18089 148904 -18045
rect 148948 -18089 149004 -18045
rect 149048 -18089 149104 -18045
rect 149148 -18089 149204 -18045
rect 149248 -18089 149304 -18045
rect 149348 -18089 149404 -18045
rect 149448 -18089 149504 -18045
rect 149548 -18089 149604 -18045
rect 149648 -18089 149704 -18045
rect 149748 -18089 149804 -18045
rect 149848 -18089 149904 -18045
rect 149948 -18089 150004 -18045
rect 150048 -18089 150104 -18045
rect 150148 -18089 150204 -18045
rect 150248 -18089 150304 -18045
rect 150348 -18089 150404 -18045
rect 150448 -18089 150904 -18045
rect 150948 -18089 151004 -18045
rect 151048 -18089 151104 -18045
rect 151148 -18089 151204 -18045
rect 151248 -18089 151304 -18045
rect 151348 -18089 151404 -18045
rect 151448 -18089 151504 -18045
rect 151548 -18089 151604 -18045
rect 151648 -18089 151704 -18045
rect 151748 -18089 151804 -18045
rect 151848 -18089 151904 -18045
rect 151948 -18089 152004 -18045
rect 152048 -18089 152104 -18045
rect 152148 -18089 152204 -18045
rect 152248 -18089 152304 -18045
rect 152348 -18089 152404 -18045
rect 152448 -18089 154949 -18045
rect 142660 -18145 154949 -18089
rect 142660 -18189 144904 -18145
rect 144948 -18189 145004 -18145
rect 145048 -18189 145104 -18145
rect 145148 -18189 145204 -18145
rect 145248 -18189 145304 -18145
rect 145348 -18189 145404 -18145
rect 145448 -18189 145504 -18145
rect 145548 -18189 145604 -18145
rect 145648 -18189 145704 -18145
rect 145748 -18189 145804 -18145
rect 145848 -18189 145904 -18145
rect 145948 -18189 146004 -18145
rect 146048 -18189 146104 -18145
rect 146148 -18189 146204 -18145
rect 146248 -18189 146304 -18145
rect 146348 -18189 146404 -18145
rect 146448 -18189 146904 -18145
rect 146948 -18189 147004 -18145
rect 147048 -18189 147104 -18145
rect 147148 -18189 147204 -18145
rect 147248 -18189 147304 -18145
rect 147348 -18189 147404 -18145
rect 147448 -18189 147504 -18145
rect 147548 -18189 147604 -18145
rect 147648 -18189 147704 -18145
rect 147748 -18189 147804 -18145
rect 147848 -18189 147904 -18145
rect 147948 -18189 148004 -18145
rect 148048 -18189 148104 -18145
rect 148148 -18189 148204 -18145
rect 148248 -18189 148304 -18145
rect 148348 -18189 148404 -18145
rect 148448 -18189 148904 -18145
rect 148948 -18189 149004 -18145
rect 149048 -18189 149104 -18145
rect 149148 -18189 149204 -18145
rect 149248 -18189 149304 -18145
rect 149348 -18189 149404 -18145
rect 149448 -18189 149504 -18145
rect 149548 -18189 149604 -18145
rect 149648 -18189 149704 -18145
rect 149748 -18189 149804 -18145
rect 149848 -18189 149904 -18145
rect 149948 -18189 150004 -18145
rect 150048 -18189 150104 -18145
rect 150148 -18189 150204 -18145
rect 150248 -18189 150304 -18145
rect 150348 -18189 150404 -18145
rect 150448 -18189 150904 -18145
rect 150948 -18189 151004 -18145
rect 151048 -18189 151104 -18145
rect 151148 -18189 151204 -18145
rect 151248 -18189 151304 -18145
rect 151348 -18189 151404 -18145
rect 151448 -18189 151504 -18145
rect 151548 -18189 151604 -18145
rect 151648 -18189 151704 -18145
rect 151748 -18189 151804 -18145
rect 151848 -18189 151904 -18145
rect 151948 -18189 152004 -18145
rect 152048 -18189 152104 -18145
rect 152148 -18189 152204 -18145
rect 152248 -18189 152304 -18145
rect 152348 -18189 152404 -18145
rect 152448 -18189 154949 -18145
rect 142660 -18245 154949 -18189
rect 142660 -18289 144904 -18245
rect 144948 -18289 145004 -18245
rect 145048 -18289 145104 -18245
rect 145148 -18289 145204 -18245
rect 145248 -18289 145304 -18245
rect 145348 -18289 145404 -18245
rect 145448 -18289 145504 -18245
rect 145548 -18289 145604 -18245
rect 145648 -18289 145704 -18245
rect 145748 -18289 145804 -18245
rect 145848 -18289 145904 -18245
rect 145948 -18289 146004 -18245
rect 146048 -18289 146104 -18245
rect 146148 -18289 146204 -18245
rect 146248 -18289 146304 -18245
rect 146348 -18289 146404 -18245
rect 146448 -18289 146904 -18245
rect 146948 -18289 147004 -18245
rect 147048 -18289 147104 -18245
rect 147148 -18289 147204 -18245
rect 147248 -18289 147304 -18245
rect 147348 -18289 147404 -18245
rect 147448 -18289 147504 -18245
rect 147548 -18289 147604 -18245
rect 147648 -18289 147704 -18245
rect 147748 -18289 147804 -18245
rect 147848 -18289 147904 -18245
rect 147948 -18289 148004 -18245
rect 148048 -18289 148104 -18245
rect 148148 -18289 148204 -18245
rect 148248 -18289 148304 -18245
rect 148348 -18289 148404 -18245
rect 148448 -18289 148904 -18245
rect 148948 -18289 149004 -18245
rect 149048 -18289 149104 -18245
rect 149148 -18289 149204 -18245
rect 149248 -18289 149304 -18245
rect 149348 -18289 149404 -18245
rect 149448 -18289 149504 -18245
rect 149548 -18289 149604 -18245
rect 149648 -18289 149704 -18245
rect 149748 -18289 149804 -18245
rect 149848 -18289 149904 -18245
rect 149948 -18289 150004 -18245
rect 150048 -18289 150104 -18245
rect 150148 -18289 150204 -18245
rect 150248 -18289 150304 -18245
rect 150348 -18289 150404 -18245
rect 150448 -18289 150904 -18245
rect 150948 -18289 151004 -18245
rect 151048 -18289 151104 -18245
rect 151148 -18289 151204 -18245
rect 151248 -18289 151304 -18245
rect 151348 -18289 151404 -18245
rect 151448 -18289 151504 -18245
rect 151548 -18289 151604 -18245
rect 151648 -18289 151704 -18245
rect 151748 -18289 151804 -18245
rect 151848 -18289 151904 -18245
rect 151948 -18289 152004 -18245
rect 152048 -18289 152104 -18245
rect 152148 -18289 152204 -18245
rect 152248 -18289 152304 -18245
rect 152348 -18289 152404 -18245
rect 152448 -18289 154949 -18245
rect 142660 -18345 154949 -18289
rect 142660 -18389 144904 -18345
rect 144948 -18389 145004 -18345
rect 145048 -18389 145104 -18345
rect 145148 -18389 145204 -18345
rect 145248 -18389 145304 -18345
rect 145348 -18389 145404 -18345
rect 145448 -18389 145504 -18345
rect 145548 -18389 145604 -18345
rect 145648 -18389 145704 -18345
rect 145748 -18389 145804 -18345
rect 145848 -18389 145904 -18345
rect 145948 -18389 146004 -18345
rect 146048 -18389 146104 -18345
rect 146148 -18389 146204 -18345
rect 146248 -18389 146304 -18345
rect 146348 -18389 146404 -18345
rect 146448 -18389 146904 -18345
rect 146948 -18389 147004 -18345
rect 147048 -18389 147104 -18345
rect 147148 -18389 147204 -18345
rect 147248 -18389 147304 -18345
rect 147348 -18389 147404 -18345
rect 147448 -18389 147504 -18345
rect 147548 -18389 147604 -18345
rect 147648 -18389 147704 -18345
rect 147748 -18389 147804 -18345
rect 147848 -18389 147904 -18345
rect 147948 -18389 148004 -18345
rect 148048 -18389 148104 -18345
rect 148148 -18389 148204 -18345
rect 148248 -18389 148304 -18345
rect 148348 -18389 148404 -18345
rect 148448 -18389 148904 -18345
rect 148948 -18389 149004 -18345
rect 149048 -18389 149104 -18345
rect 149148 -18389 149204 -18345
rect 149248 -18389 149304 -18345
rect 149348 -18389 149404 -18345
rect 149448 -18389 149504 -18345
rect 149548 -18389 149604 -18345
rect 149648 -18389 149704 -18345
rect 149748 -18389 149804 -18345
rect 149848 -18389 149904 -18345
rect 149948 -18389 150004 -18345
rect 150048 -18389 150104 -18345
rect 150148 -18389 150204 -18345
rect 150248 -18389 150304 -18345
rect 150348 -18389 150404 -18345
rect 150448 -18389 150904 -18345
rect 150948 -18389 151004 -18345
rect 151048 -18389 151104 -18345
rect 151148 -18389 151204 -18345
rect 151248 -18389 151304 -18345
rect 151348 -18389 151404 -18345
rect 151448 -18389 151504 -18345
rect 151548 -18389 151604 -18345
rect 151648 -18389 151704 -18345
rect 151748 -18389 151804 -18345
rect 151848 -18389 151904 -18345
rect 151948 -18389 152004 -18345
rect 152048 -18389 152104 -18345
rect 152148 -18389 152204 -18345
rect 152248 -18389 152304 -18345
rect 152348 -18389 152404 -18345
rect 152448 -18389 154949 -18345
rect 142660 -18445 154949 -18389
rect 142660 -18489 144904 -18445
rect 144948 -18489 145004 -18445
rect 145048 -18489 145104 -18445
rect 145148 -18489 145204 -18445
rect 145248 -18489 145304 -18445
rect 145348 -18489 145404 -18445
rect 145448 -18489 145504 -18445
rect 145548 -18489 145604 -18445
rect 145648 -18489 145704 -18445
rect 145748 -18489 145804 -18445
rect 145848 -18489 145904 -18445
rect 145948 -18489 146004 -18445
rect 146048 -18489 146104 -18445
rect 146148 -18489 146204 -18445
rect 146248 -18489 146304 -18445
rect 146348 -18489 146404 -18445
rect 146448 -18489 146904 -18445
rect 146948 -18489 147004 -18445
rect 147048 -18489 147104 -18445
rect 147148 -18489 147204 -18445
rect 147248 -18489 147304 -18445
rect 147348 -18489 147404 -18445
rect 147448 -18489 147504 -18445
rect 147548 -18489 147604 -18445
rect 147648 -18489 147704 -18445
rect 147748 -18489 147804 -18445
rect 147848 -18489 147904 -18445
rect 147948 -18489 148004 -18445
rect 148048 -18489 148104 -18445
rect 148148 -18489 148204 -18445
rect 148248 -18489 148304 -18445
rect 148348 -18489 148404 -18445
rect 148448 -18489 148904 -18445
rect 148948 -18489 149004 -18445
rect 149048 -18489 149104 -18445
rect 149148 -18489 149204 -18445
rect 149248 -18489 149304 -18445
rect 149348 -18489 149404 -18445
rect 149448 -18489 149504 -18445
rect 149548 -18489 149604 -18445
rect 149648 -18489 149704 -18445
rect 149748 -18489 149804 -18445
rect 149848 -18489 149904 -18445
rect 149948 -18489 150004 -18445
rect 150048 -18489 150104 -18445
rect 150148 -18489 150204 -18445
rect 150248 -18489 150304 -18445
rect 150348 -18489 150404 -18445
rect 150448 -18489 150904 -18445
rect 150948 -18489 151004 -18445
rect 151048 -18489 151104 -18445
rect 151148 -18489 151204 -18445
rect 151248 -18489 151304 -18445
rect 151348 -18489 151404 -18445
rect 151448 -18489 151504 -18445
rect 151548 -18489 151604 -18445
rect 151648 -18489 151704 -18445
rect 151748 -18489 151804 -18445
rect 151848 -18489 151904 -18445
rect 151948 -18489 152004 -18445
rect 152048 -18489 152104 -18445
rect 152148 -18489 152204 -18445
rect 152248 -18489 152304 -18445
rect 152348 -18489 152404 -18445
rect 152448 -18489 154949 -18445
rect 142660 -18545 154949 -18489
rect 142660 -18589 144904 -18545
rect 144948 -18589 145004 -18545
rect 145048 -18589 145104 -18545
rect 145148 -18589 145204 -18545
rect 145248 -18589 145304 -18545
rect 145348 -18589 145404 -18545
rect 145448 -18589 145504 -18545
rect 145548 -18589 145604 -18545
rect 145648 -18589 145704 -18545
rect 145748 -18589 145804 -18545
rect 145848 -18589 145904 -18545
rect 145948 -18589 146004 -18545
rect 146048 -18589 146104 -18545
rect 146148 -18589 146204 -18545
rect 146248 -18589 146304 -18545
rect 146348 -18589 146404 -18545
rect 146448 -18589 146904 -18545
rect 146948 -18589 147004 -18545
rect 147048 -18589 147104 -18545
rect 147148 -18589 147204 -18545
rect 147248 -18589 147304 -18545
rect 147348 -18589 147404 -18545
rect 147448 -18589 147504 -18545
rect 147548 -18589 147604 -18545
rect 147648 -18589 147704 -18545
rect 147748 -18589 147804 -18545
rect 147848 -18589 147904 -18545
rect 147948 -18589 148004 -18545
rect 148048 -18589 148104 -18545
rect 148148 -18589 148204 -18545
rect 148248 -18589 148304 -18545
rect 148348 -18589 148404 -18545
rect 148448 -18589 148904 -18545
rect 148948 -18589 149004 -18545
rect 149048 -18589 149104 -18545
rect 149148 -18589 149204 -18545
rect 149248 -18589 149304 -18545
rect 149348 -18589 149404 -18545
rect 149448 -18589 149504 -18545
rect 149548 -18589 149604 -18545
rect 149648 -18589 149704 -18545
rect 149748 -18589 149804 -18545
rect 149848 -18589 149904 -18545
rect 149948 -18589 150004 -18545
rect 150048 -18589 150104 -18545
rect 150148 -18589 150204 -18545
rect 150248 -18589 150304 -18545
rect 150348 -18589 150404 -18545
rect 150448 -18589 150904 -18545
rect 150948 -18589 151004 -18545
rect 151048 -18589 151104 -18545
rect 151148 -18589 151204 -18545
rect 151248 -18589 151304 -18545
rect 151348 -18589 151404 -18545
rect 151448 -18589 151504 -18545
rect 151548 -18589 151604 -18545
rect 151648 -18589 151704 -18545
rect 151748 -18589 151804 -18545
rect 151848 -18589 151904 -18545
rect 151948 -18589 152004 -18545
rect 152048 -18589 152104 -18545
rect 152148 -18589 152204 -18545
rect 152248 -18589 152304 -18545
rect 152348 -18589 152404 -18545
rect 152448 -18589 154949 -18545
rect 142660 -18645 154949 -18589
rect 173132 -17214 174740 -13446
rect 173132 -17830 173611 -17214
rect 174124 -17830 174740 -17214
rect 173132 -18617 174740 -17830
rect 142660 -18689 144904 -18645
rect 144948 -18689 145004 -18645
rect 145048 -18689 145104 -18645
rect 145148 -18689 145204 -18645
rect 145248 -18689 145304 -18645
rect 145348 -18689 145404 -18645
rect 145448 -18689 145504 -18645
rect 145548 -18689 145604 -18645
rect 145648 -18689 145704 -18645
rect 145748 -18689 145804 -18645
rect 145848 -18689 145904 -18645
rect 145948 -18689 146004 -18645
rect 146048 -18689 146104 -18645
rect 146148 -18689 146204 -18645
rect 146248 -18689 146304 -18645
rect 146348 -18689 146404 -18645
rect 146448 -18689 146904 -18645
rect 146948 -18689 147004 -18645
rect 147048 -18689 147104 -18645
rect 147148 -18689 147204 -18645
rect 147248 -18689 147304 -18645
rect 147348 -18689 147404 -18645
rect 147448 -18689 147504 -18645
rect 147548 -18689 147604 -18645
rect 147648 -18689 147704 -18645
rect 147748 -18689 147804 -18645
rect 147848 -18689 147904 -18645
rect 147948 -18689 148004 -18645
rect 148048 -18689 148104 -18645
rect 148148 -18689 148204 -18645
rect 148248 -18689 148304 -18645
rect 148348 -18689 148404 -18645
rect 148448 -18689 148904 -18645
rect 148948 -18689 149004 -18645
rect 149048 -18689 149104 -18645
rect 149148 -18689 149204 -18645
rect 149248 -18689 149304 -18645
rect 149348 -18689 149404 -18645
rect 149448 -18689 149504 -18645
rect 149548 -18689 149604 -18645
rect 149648 -18689 149704 -18645
rect 149748 -18689 149804 -18645
rect 149848 -18689 149904 -18645
rect 149948 -18689 150004 -18645
rect 150048 -18689 150104 -18645
rect 150148 -18689 150204 -18645
rect 150248 -18689 150304 -18645
rect 150348 -18689 150404 -18645
rect 150448 -18689 150904 -18645
rect 150948 -18689 151004 -18645
rect 151048 -18689 151104 -18645
rect 151148 -18689 151204 -18645
rect 151248 -18689 151304 -18645
rect 151348 -18689 151404 -18645
rect 151448 -18689 151504 -18645
rect 151548 -18689 151604 -18645
rect 151648 -18689 151704 -18645
rect 151748 -18689 151804 -18645
rect 151848 -18689 151904 -18645
rect 151948 -18689 152004 -18645
rect 152048 -18689 152104 -18645
rect 152148 -18689 152204 -18645
rect 152248 -18689 152304 -18645
rect 152348 -18689 152404 -18645
rect 152448 -18689 154949 -18645
rect 142660 -18745 154949 -18689
rect 142660 -18789 144904 -18745
rect 144948 -18789 145004 -18745
rect 145048 -18789 145104 -18745
rect 145148 -18789 145204 -18745
rect 145248 -18789 145304 -18745
rect 145348 -18789 145404 -18745
rect 145448 -18789 145504 -18745
rect 145548 -18789 145604 -18745
rect 145648 -18789 145704 -18745
rect 145748 -18789 145804 -18745
rect 145848 -18789 145904 -18745
rect 145948 -18789 146004 -18745
rect 146048 -18789 146104 -18745
rect 146148 -18789 146204 -18745
rect 146248 -18789 146304 -18745
rect 146348 -18789 146404 -18745
rect 146448 -18789 146904 -18745
rect 146948 -18789 147004 -18745
rect 147048 -18789 147104 -18745
rect 147148 -18789 147204 -18745
rect 147248 -18789 147304 -18745
rect 147348 -18789 147404 -18745
rect 147448 -18789 147504 -18745
rect 147548 -18789 147604 -18745
rect 147648 -18789 147704 -18745
rect 147748 -18789 147804 -18745
rect 147848 -18789 147904 -18745
rect 147948 -18789 148004 -18745
rect 148048 -18789 148104 -18745
rect 148148 -18789 148204 -18745
rect 148248 -18789 148304 -18745
rect 148348 -18789 148404 -18745
rect 148448 -18789 148904 -18745
rect 148948 -18789 149004 -18745
rect 149048 -18789 149104 -18745
rect 149148 -18789 149204 -18745
rect 149248 -18789 149304 -18745
rect 149348 -18789 149404 -18745
rect 149448 -18789 149504 -18745
rect 149548 -18789 149604 -18745
rect 149648 -18789 149704 -18745
rect 149748 -18789 149804 -18745
rect 149848 -18789 149904 -18745
rect 149948 -18789 150004 -18745
rect 150048 -18789 150104 -18745
rect 150148 -18789 150204 -18745
rect 150248 -18789 150304 -18745
rect 150348 -18789 150404 -18745
rect 150448 -18789 150904 -18745
rect 150948 -18789 151004 -18745
rect 151048 -18789 151104 -18745
rect 151148 -18789 151204 -18745
rect 151248 -18789 151304 -18745
rect 151348 -18789 151404 -18745
rect 151448 -18789 151504 -18745
rect 151548 -18789 151604 -18745
rect 151648 -18789 151704 -18745
rect 151748 -18789 151804 -18745
rect 151848 -18789 151904 -18745
rect 151948 -18789 152004 -18745
rect 152048 -18789 152104 -18745
rect 152148 -18789 152204 -18745
rect 152248 -18789 152304 -18745
rect 152348 -18789 152404 -18745
rect 152448 -18789 154949 -18745
rect 142660 -18845 154949 -18789
rect 142660 -18889 144904 -18845
rect 144948 -18889 145004 -18845
rect 145048 -18889 145104 -18845
rect 145148 -18889 145204 -18845
rect 145248 -18889 145304 -18845
rect 145348 -18889 145404 -18845
rect 145448 -18889 145504 -18845
rect 145548 -18889 145604 -18845
rect 145648 -18889 145704 -18845
rect 145748 -18889 145804 -18845
rect 145848 -18889 145904 -18845
rect 145948 -18889 146004 -18845
rect 146048 -18889 146104 -18845
rect 146148 -18889 146204 -18845
rect 146248 -18889 146304 -18845
rect 146348 -18889 146404 -18845
rect 146448 -18889 146904 -18845
rect 146948 -18889 147004 -18845
rect 147048 -18889 147104 -18845
rect 147148 -18889 147204 -18845
rect 147248 -18889 147304 -18845
rect 147348 -18889 147404 -18845
rect 147448 -18889 147504 -18845
rect 147548 -18889 147604 -18845
rect 147648 -18889 147704 -18845
rect 147748 -18889 147804 -18845
rect 147848 -18889 147904 -18845
rect 147948 -18889 148004 -18845
rect 148048 -18889 148104 -18845
rect 148148 -18889 148204 -18845
rect 148248 -18889 148304 -18845
rect 148348 -18889 148404 -18845
rect 148448 -18889 148904 -18845
rect 148948 -18889 149004 -18845
rect 149048 -18889 149104 -18845
rect 149148 -18889 149204 -18845
rect 149248 -18889 149304 -18845
rect 149348 -18889 149404 -18845
rect 149448 -18889 149504 -18845
rect 149548 -18889 149604 -18845
rect 149648 -18889 149704 -18845
rect 149748 -18889 149804 -18845
rect 149848 -18889 149904 -18845
rect 149948 -18889 150004 -18845
rect 150048 -18889 150104 -18845
rect 150148 -18889 150204 -18845
rect 150248 -18889 150304 -18845
rect 150348 -18889 150404 -18845
rect 150448 -18889 150904 -18845
rect 150948 -18889 151004 -18845
rect 151048 -18889 151104 -18845
rect 151148 -18889 151204 -18845
rect 151248 -18889 151304 -18845
rect 151348 -18889 151404 -18845
rect 151448 -18889 151504 -18845
rect 151548 -18889 151604 -18845
rect 151648 -18889 151704 -18845
rect 151748 -18889 151804 -18845
rect 151848 -18889 151904 -18845
rect 151948 -18889 152004 -18845
rect 152048 -18889 152104 -18845
rect 152148 -18889 152204 -18845
rect 152248 -18889 152304 -18845
rect 152348 -18889 152404 -18845
rect 152448 -18889 154949 -18845
rect 142660 -18945 154949 -18889
rect 142660 -18989 144904 -18945
rect 144948 -18989 145004 -18945
rect 145048 -18989 145104 -18945
rect 145148 -18989 145204 -18945
rect 145248 -18989 145304 -18945
rect 145348 -18989 145404 -18945
rect 145448 -18989 145504 -18945
rect 145548 -18989 145604 -18945
rect 145648 -18989 145704 -18945
rect 145748 -18989 145804 -18945
rect 145848 -18989 145904 -18945
rect 145948 -18989 146004 -18945
rect 146048 -18989 146104 -18945
rect 146148 -18989 146204 -18945
rect 146248 -18989 146304 -18945
rect 146348 -18989 146404 -18945
rect 146448 -18989 146904 -18945
rect 146948 -18989 147004 -18945
rect 147048 -18989 147104 -18945
rect 147148 -18989 147204 -18945
rect 147248 -18989 147304 -18945
rect 147348 -18989 147404 -18945
rect 147448 -18989 147504 -18945
rect 147548 -18989 147604 -18945
rect 147648 -18989 147704 -18945
rect 147748 -18989 147804 -18945
rect 147848 -18989 147904 -18945
rect 147948 -18989 148004 -18945
rect 148048 -18989 148104 -18945
rect 148148 -18989 148204 -18945
rect 148248 -18989 148304 -18945
rect 148348 -18989 148404 -18945
rect 148448 -18989 148904 -18945
rect 148948 -18989 149004 -18945
rect 149048 -18989 149104 -18945
rect 149148 -18989 149204 -18945
rect 149248 -18989 149304 -18945
rect 149348 -18989 149404 -18945
rect 149448 -18989 149504 -18945
rect 149548 -18989 149604 -18945
rect 149648 -18989 149704 -18945
rect 149748 -18989 149804 -18945
rect 149848 -18989 149904 -18945
rect 149948 -18989 150004 -18945
rect 150048 -18989 150104 -18945
rect 150148 -18989 150204 -18945
rect 150248 -18989 150304 -18945
rect 150348 -18989 150404 -18945
rect 150448 -18989 150904 -18945
rect 150948 -18989 151004 -18945
rect 151048 -18989 151104 -18945
rect 151148 -18989 151204 -18945
rect 151248 -18989 151304 -18945
rect 151348 -18989 151404 -18945
rect 151448 -18989 151504 -18945
rect 151548 -18989 151604 -18945
rect 151648 -18989 151704 -18945
rect 151748 -18989 151804 -18945
rect 151848 -18989 151904 -18945
rect 151948 -18989 152004 -18945
rect 152048 -18989 152104 -18945
rect 152148 -18989 152204 -18945
rect 152248 -18989 152304 -18945
rect 152348 -18989 152404 -18945
rect 152448 -18989 154949 -18945
rect 79796 -24026 89254 -23015
rect 79796 -24070 80849 -24026
rect 80893 -24070 80949 -24026
rect 80993 -24070 81049 -24026
rect 81093 -24070 81149 -24026
rect 81193 -24070 81249 -24026
rect 81293 -24070 81349 -24026
rect 81393 -24070 81449 -24026
rect 81493 -24070 81549 -24026
rect 81593 -24070 81649 -24026
rect 81693 -24070 81749 -24026
rect 81793 -24070 81849 -24026
rect 81893 -24070 81949 -24026
rect 81993 -24070 82049 -24026
rect 82093 -24070 82149 -24026
rect 82193 -24070 82249 -24026
rect 82293 -24070 82349 -24026
rect 82393 -24070 82849 -24026
rect 82893 -24070 82949 -24026
rect 82993 -24070 83049 -24026
rect 83093 -24070 83149 -24026
rect 83193 -24070 83249 -24026
rect 83293 -24070 83349 -24026
rect 83393 -24070 83449 -24026
rect 83493 -24070 83549 -24026
rect 83593 -24070 83649 -24026
rect 83693 -24070 83749 -24026
rect 83793 -24070 83849 -24026
rect 83893 -24070 83949 -24026
rect 83993 -24070 84049 -24026
rect 84093 -24070 84149 -24026
rect 84193 -24070 84249 -24026
rect 84293 -24070 84349 -24026
rect 84393 -24070 84849 -24026
rect 84893 -24070 84949 -24026
rect 84993 -24070 85049 -24026
rect 85093 -24070 85149 -24026
rect 85193 -24070 85249 -24026
rect 85293 -24070 85349 -24026
rect 85393 -24070 85449 -24026
rect 85493 -24070 85549 -24026
rect 85593 -24070 85649 -24026
rect 85693 -24070 85749 -24026
rect 85793 -24070 85849 -24026
rect 85893 -24070 85949 -24026
rect 85993 -24070 86049 -24026
rect 86093 -24070 86149 -24026
rect 86193 -24070 86249 -24026
rect 86293 -24070 86349 -24026
rect 86393 -24070 86849 -24026
rect 86893 -24070 86949 -24026
rect 86993 -24070 87049 -24026
rect 87093 -24070 87149 -24026
rect 87193 -24070 87249 -24026
rect 87293 -24070 87349 -24026
rect 87393 -24070 87449 -24026
rect 87493 -24070 87549 -24026
rect 87593 -24070 87649 -24026
rect 87693 -24070 87749 -24026
rect 87793 -24070 87849 -24026
rect 87893 -24070 87949 -24026
rect 87993 -24070 88049 -24026
rect 88093 -24070 88149 -24026
rect 88193 -24070 88249 -24026
rect 88293 -24070 88349 -24026
rect 88393 -24070 89254 -24026
rect 79796 -24126 89254 -24070
rect 79796 -24170 80849 -24126
rect 80893 -24170 80949 -24126
rect 80993 -24170 81049 -24126
rect 81093 -24170 81149 -24126
rect 81193 -24170 81249 -24126
rect 81293 -24170 81349 -24126
rect 81393 -24170 81449 -24126
rect 81493 -24170 81549 -24126
rect 81593 -24170 81649 -24126
rect 81693 -24170 81749 -24126
rect 81793 -24170 81849 -24126
rect 81893 -24170 81949 -24126
rect 81993 -24170 82049 -24126
rect 82093 -24170 82149 -24126
rect 82193 -24170 82249 -24126
rect 82293 -24170 82349 -24126
rect 82393 -24170 82849 -24126
rect 82893 -24170 82949 -24126
rect 82993 -24170 83049 -24126
rect 83093 -24170 83149 -24126
rect 83193 -24170 83249 -24126
rect 83293 -24170 83349 -24126
rect 83393 -24170 83449 -24126
rect 83493 -24170 83549 -24126
rect 83593 -24170 83649 -24126
rect 83693 -24170 83749 -24126
rect 83793 -24170 83849 -24126
rect 83893 -24170 83949 -24126
rect 83993 -24170 84049 -24126
rect 84093 -24170 84149 -24126
rect 84193 -24170 84249 -24126
rect 84293 -24170 84349 -24126
rect 84393 -24170 84849 -24126
rect 84893 -24170 84949 -24126
rect 84993 -24170 85049 -24126
rect 85093 -24170 85149 -24126
rect 85193 -24170 85249 -24126
rect 85293 -24170 85349 -24126
rect 85393 -24170 85449 -24126
rect 85493 -24170 85549 -24126
rect 85593 -24170 85649 -24126
rect 85693 -24170 85749 -24126
rect 85793 -24170 85849 -24126
rect 85893 -24170 85949 -24126
rect 85993 -24170 86049 -24126
rect 86093 -24170 86149 -24126
rect 86193 -24170 86249 -24126
rect 86293 -24170 86349 -24126
rect 86393 -24170 86849 -24126
rect 86893 -24170 86949 -24126
rect 86993 -24170 87049 -24126
rect 87093 -24170 87149 -24126
rect 87193 -24170 87249 -24126
rect 87293 -24170 87349 -24126
rect 87393 -24170 87449 -24126
rect 87493 -24170 87549 -24126
rect 87593 -24170 87649 -24126
rect 87693 -24170 87749 -24126
rect 87793 -24170 87849 -24126
rect 87893 -24170 87949 -24126
rect 87993 -24170 88049 -24126
rect 88093 -24170 88149 -24126
rect 88193 -24170 88249 -24126
rect 88293 -24170 88349 -24126
rect 88393 -24170 89254 -24126
rect 79796 -24226 89254 -24170
rect 79796 -24270 80849 -24226
rect 80893 -24270 80949 -24226
rect 80993 -24270 81049 -24226
rect 81093 -24270 81149 -24226
rect 81193 -24270 81249 -24226
rect 81293 -24270 81349 -24226
rect 81393 -24270 81449 -24226
rect 81493 -24270 81549 -24226
rect 81593 -24270 81649 -24226
rect 81693 -24270 81749 -24226
rect 81793 -24270 81849 -24226
rect 81893 -24270 81949 -24226
rect 81993 -24270 82049 -24226
rect 82093 -24270 82149 -24226
rect 82193 -24270 82249 -24226
rect 82293 -24270 82349 -24226
rect 82393 -24270 82849 -24226
rect 82893 -24270 82949 -24226
rect 82993 -24270 83049 -24226
rect 83093 -24270 83149 -24226
rect 83193 -24270 83249 -24226
rect 83293 -24270 83349 -24226
rect 83393 -24270 83449 -24226
rect 83493 -24270 83549 -24226
rect 83593 -24270 83649 -24226
rect 83693 -24270 83749 -24226
rect 83793 -24270 83849 -24226
rect 83893 -24270 83949 -24226
rect 83993 -24270 84049 -24226
rect 84093 -24270 84149 -24226
rect 84193 -24270 84249 -24226
rect 84293 -24270 84349 -24226
rect 84393 -24270 84849 -24226
rect 84893 -24270 84949 -24226
rect 84993 -24270 85049 -24226
rect 85093 -24270 85149 -24226
rect 85193 -24270 85249 -24226
rect 85293 -24270 85349 -24226
rect 85393 -24270 85449 -24226
rect 85493 -24270 85549 -24226
rect 85593 -24270 85649 -24226
rect 85693 -24270 85749 -24226
rect 85793 -24270 85849 -24226
rect 85893 -24270 85949 -24226
rect 85993 -24270 86049 -24226
rect 86093 -24270 86149 -24226
rect 86193 -24270 86249 -24226
rect 86293 -24270 86349 -24226
rect 86393 -24270 86849 -24226
rect 86893 -24270 86949 -24226
rect 86993 -24270 87049 -24226
rect 87093 -24270 87149 -24226
rect 87193 -24270 87249 -24226
rect 87293 -24270 87349 -24226
rect 87393 -24270 87449 -24226
rect 87493 -24270 87549 -24226
rect 87593 -24270 87649 -24226
rect 87693 -24270 87749 -24226
rect 87793 -24270 87849 -24226
rect 87893 -24270 87949 -24226
rect 87993 -24270 88049 -24226
rect 88093 -24270 88149 -24226
rect 88193 -24270 88249 -24226
rect 88293 -24270 88349 -24226
rect 88393 -24270 89254 -24226
rect 79796 -24326 89254 -24270
rect 79796 -24370 80849 -24326
rect 80893 -24370 80949 -24326
rect 80993 -24370 81049 -24326
rect 81093 -24370 81149 -24326
rect 81193 -24370 81249 -24326
rect 81293 -24370 81349 -24326
rect 81393 -24370 81449 -24326
rect 81493 -24370 81549 -24326
rect 81593 -24370 81649 -24326
rect 81693 -24370 81749 -24326
rect 81793 -24370 81849 -24326
rect 81893 -24370 81949 -24326
rect 81993 -24370 82049 -24326
rect 82093 -24370 82149 -24326
rect 82193 -24370 82249 -24326
rect 82293 -24370 82349 -24326
rect 82393 -24370 82849 -24326
rect 82893 -24370 82949 -24326
rect 82993 -24370 83049 -24326
rect 83093 -24370 83149 -24326
rect 83193 -24370 83249 -24326
rect 83293 -24370 83349 -24326
rect 83393 -24370 83449 -24326
rect 83493 -24370 83549 -24326
rect 83593 -24370 83649 -24326
rect 83693 -24370 83749 -24326
rect 83793 -24370 83849 -24326
rect 83893 -24370 83949 -24326
rect 83993 -24370 84049 -24326
rect 84093 -24370 84149 -24326
rect 84193 -24370 84249 -24326
rect 84293 -24370 84349 -24326
rect 84393 -24370 84849 -24326
rect 84893 -24370 84949 -24326
rect 84993 -24370 85049 -24326
rect 85093 -24370 85149 -24326
rect 85193 -24370 85249 -24326
rect 85293 -24370 85349 -24326
rect 85393 -24370 85449 -24326
rect 85493 -24370 85549 -24326
rect 85593 -24370 85649 -24326
rect 85693 -24370 85749 -24326
rect 85793 -24370 85849 -24326
rect 85893 -24370 85949 -24326
rect 85993 -24370 86049 -24326
rect 86093 -24370 86149 -24326
rect 86193 -24370 86249 -24326
rect 86293 -24370 86349 -24326
rect 86393 -24370 86849 -24326
rect 86893 -24370 86949 -24326
rect 86993 -24370 87049 -24326
rect 87093 -24370 87149 -24326
rect 87193 -24370 87249 -24326
rect 87293 -24370 87349 -24326
rect 87393 -24370 87449 -24326
rect 87493 -24370 87549 -24326
rect 87593 -24370 87649 -24326
rect 87693 -24370 87749 -24326
rect 87793 -24370 87849 -24326
rect 87893 -24370 87949 -24326
rect 87993 -24370 88049 -24326
rect 88093 -24370 88149 -24326
rect 88193 -24370 88249 -24326
rect 88293 -24370 88349 -24326
rect 88393 -24370 89254 -24326
rect 79796 -24426 89254 -24370
rect 79796 -24470 80849 -24426
rect 80893 -24470 80949 -24426
rect 80993 -24470 81049 -24426
rect 81093 -24470 81149 -24426
rect 81193 -24470 81249 -24426
rect 81293 -24470 81349 -24426
rect 81393 -24470 81449 -24426
rect 81493 -24470 81549 -24426
rect 81593 -24470 81649 -24426
rect 81693 -24470 81749 -24426
rect 81793 -24470 81849 -24426
rect 81893 -24470 81949 -24426
rect 81993 -24470 82049 -24426
rect 82093 -24470 82149 -24426
rect 82193 -24470 82249 -24426
rect 82293 -24470 82349 -24426
rect 82393 -24470 82849 -24426
rect 82893 -24470 82949 -24426
rect 82993 -24470 83049 -24426
rect 83093 -24470 83149 -24426
rect 83193 -24470 83249 -24426
rect 83293 -24470 83349 -24426
rect 83393 -24470 83449 -24426
rect 83493 -24470 83549 -24426
rect 83593 -24470 83649 -24426
rect 83693 -24470 83749 -24426
rect 83793 -24470 83849 -24426
rect 83893 -24470 83949 -24426
rect 83993 -24470 84049 -24426
rect 84093 -24470 84149 -24426
rect 84193 -24470 84249 -24426
rect 84293 -24470 84349 -24426
rect 84393 -24470 84849 -24426
rect 84893 -24470 84949 -24426
rect 84993 -24470 85049 -24426
rect 85093 -24470 85149 -24426
rect 85193 -24470 85249 -24426
rect 85293 -24470 85349 -24426
rect 85393 -24470 85449 -24426
rect 85493 -24470 85549 -24426
rect 85593 -24470 85649 -24426
rect 85693 -24470 85749 -24426
rect 85793 -24470 85849 -24426
rect 85893 -24470 85949 -24426
rect 85993 -24470 86049 -24426
rect 86093 -24470 86149 -24426
rect 86193 -24470 86249 -24426
rect 86293 -24470 86349 -24426
rect 86393 -24470 86849 -24426
rect 86893 -24470 86949 -24426
rect 86993 -24470 87049 -24426
rect 87093 -24470 87149 -24426
rect 87193 -24470 87249 -24426
rect 87293 -24470 87349 -24426
rect 87393 -24470 87449 -24426
rect 87493 -24470 87549 -24426
rect 87593 -24470 87649 -24426
rect 87693 -24470 87749 -24426
rect 87793 -24470 87849 -24426
rect 87893 -24470 87949 -24426
rect 87993 -24470 88049 -24426
rect 88093 -24470 88149 -24426
rect 88193 -24470 88249 -24426
rect 88293 -24470 88349 -24426
rect 88393 -24470 89254 -24426
rect 79796 -24526 89254 -24470
rect 79796 -24570 80849 -24526
rect 80893 -24570 80949 -24526
rect 80993 -24570 81049 -24526
rect 81093 -24570 81149 -24526
rect 81193 -24570 81249 -24526
rect 81293 -24570 81349 -24526
rect 81393 -24570 81449 -24526
rect 81493 -24570 81549 -24526
rect 81593 -24570 81649 -24526
rect 81693 -24570 81749 -24526
rect 81793 -24570 81849 -24526
rect 81893 -24570 81949 -24526
rect 81993 -24570 82049 -24526
rect 82093 -24570 82149 -24526
rect 82193 -24570 82249 -24526
rect 82293 -24570 82349 -24526
rect 82393 -24570 82849 -24526
rect 82893 -24570 82949 -24526
rect 82993 -24570 83049 -24526
rect 83093 -24570 83149 -24526
rect 83193 -24570 83249 -24526
rect 83293 -24570 83349 -24526
rect 83393 -24570 83449 -24526
rect 83493 -24570 83549 -24526
rect 83593 -24570 83649 -24526
rect 83693 -24570 83749 -24526
rect 83793 -24570 83849 -24526
rect 83893 -24570 83949 -24526
rect 83993 -24570 84049 -24526
rect 84093 -24570 84149 -24526
rect 84193 -24570 84249 -24526
rect 84293 -24570 84349 -24526
rect 84393 -24570 84849 -24526
rect 84893 -24570 84949 -24526
rect 84993 -24570 85049 -24526
rect 85093 -24570 85149 -24526
rect 85193 -24570 85249 -24526
rect 85293 -24570 85349 -24526
rect 85393 -24570 85449 -24526
rect 85493 -24570 85549 -24526
rect 85593 -24570 85649 -24526
rect 85693 -24570 85749 -24526
rect 85793 -24570 85849 -24526
rect 85893 -24570 85949 -24526
rect 85993 -24570 86049 -24526
rect 86093 -24570 86149 -24526
rect 86193 -24570 86249 -24526
rect 86293 -24570 86349 -24526
rect 86393 -24570 86849 -24526
rect 86893 -24570 86949 -24526
rect 86993 -24570 87049 -24526
rect 87093 -24570 87149 -24526
rect 87193 -24570 87249 -24526
rect 87293 -24570 87349 -24526
rect 87393 -24570 87449 -24526
rect 87493 -24570 87549 -24526
rect 87593 -24570 87649 -24526
rect 87693 -24570 87749 -24526
rect 87793 -24570 87849 -24526
rect 87893 -24570 87949 -24526
rect 87993 -24570 88049 -24526
rect 88093 -24570 88149 -24526
rect 88193 -24570 88249 -24526
rect 88293 -24570 88349 -24526
rect 88393 -24570 89254 -24526
rect 79796 -24626 89254 -24570
rect 79796 -24670 80849 -24626
rect 80893 -24670 80949 -24626
rect 80993 -24670 81049 -24626
rect 81093 -24670 81149 -24626
rect 81193 -24670 81249 -24626
rect 81293 -24670 81349 -24626
rect 81393 -24670 81449 -24626
rect 81493 -24670 81549 -24626
rect 81593 -24670 81649 -24626
rect 81693 -24670 81749 -24626
rect 81793 -24670 81849 -24626
rect 81893 -24670 81949 -24626
rect 81993 -24670 82049 -24626
rect 82093 -24670 82149 -24626
rect 82193 -24670 82249 -24626
rect 82293 -24670 82349 -24626
rect 82393 -24670 82849 -24626
rect 82893 -24670 82949 -24626
rect 82993 -24670 83049 -24626
rect 83093 -24670 83149 -24626
rect 83193 -24670 83249 -24626
rect 83293 -24670 83349 -24626
rect 83393 -24670 83449 -24626
rect 83493 -24670 83549 -24626
rect 83593 -24670 83649 -24626
rect 83693 -24670 83749 -24626
rect 83793 -24670 83849 -24626
rect 83893 -24670 83949 -24626
rect 83993 -24670 84049 -24626
rect 84093 -24670 84149 -24626
rect 84193 -24670 84249 -24626
rect 84293 -24670 84349 -24626
rect 84393 -24670 84849 -24626
rect 84893 -24670 84949 -24626
rect 84993 -24670 85049 -24626
rect 85093 -24670 85149 -24626
rect 85193 -24670 85249 -24626
rect 85293 -24670 85349 -24626
rect 85393 -24670 85449 -24626
rect 85493 -24670 85549 -24626
rect 85593 -24670 85649 -24626
rect 85693 -24670 85749 -24626
rect 85793 -24670 85849 -24626
rect 85893 -24670 85949 -24626
rect 85993 -24670 86049 -24626
rect 86093 -24670 86149 -24626
rect 86193 -24670 86249 -24626
rect 86293 -24670 86349 -24626
rect 86393 -24670 86849 -24626
rect 86893 -24670 86949 -24626
rect 86993 -24670 87049 -24626
rect 87093 -24670 87149 -24626
rect 87193 -24670 87249 -24626
rect 87293 -24670 87349 -24626
rect 87393 -24670 87449 -24626
rect 87493 -24670 87549 -24626
rect 87593 -24670 87649 -24626
rect 87693 -24670 87749 -24626
rect 87793 -24670 87849 -24626
rect 87893 -24670 87949 -24626
rect 87993 -24670 88049 -24626
rect 88093 -24670 88149 -24626
rect 88193 -24670 88249 -24626
rect 88293 -24670 88349 -24626
rect 88393 -24670 89254 -24626
rect 79796 -24726 89254 -24670
rect 79796 -24770 80849 -24726
rect 80893 -24770 80949 -24726
rect 80993 -24770 81049 -24726
rect 81093 -24770 81149 -24726
rect 81193 -24770 81249 -24726
rect 81293 -24770 81349 -24726
rect 81393 -24770 81449 -24726
rect 81493 -24770 81549 -24726
rect 81593 -24770 81649 -24726
rect 81693 -24770 81749 -24726
rect 81793 -24770 81849 -24726
rect 81893 -24770 81949 -24726
rect 81993 -24770 82049 -24726
rect 82093 -24770 82149 -24726
rect 82193 -24770 82249 -24726
rect 82293 -24770 82349 -24726
rect 82393 -24770 82849 -24726
rect 82893 -24770 82949 -24726
rect 82993 -24770 83049 -24726
rect 83093 -24770 83149 -24726
rect 83193 -24770 83249 -24726
rect 83293 -24770 83349 -24726
rect 83393 -24770 83449 -24726
rect 83493 -24770 83549 -24726
rect 83593 -24770 83649 -24726
rect 83693 -24770 83749 -24726
rect 83793 -24770 83849 -24726
rect 83893 -24770 83949 -24726
rect 83993 -24770 84049 -24726
rect 84093 -24770 84149 -24726
rect 84193 -24770 84249 -24726
rect 84293 -24770 84349 -24726
rect 84393 -24770 84849 -24726
rect 84893 -24770 84949 -24726
rect 84993 -24770 85049 -24726
rect 85093 -24770 85149 -24726
rect 85193 -24770 85249 -24726
rect 85293 -24770 85349 -24726
rect 85393 -24770 85449 -24726
rect 85493 -24770 85549 -24726
rect 85593 -24770 85649 -24726
rect 85693 -24770 85749 -24726
rect 85793 -24770 85849 -24726
rect 85893 -24770 85949 -24726
rect 85993 -24770 86049 -24726
rect 86093 -24770 86149 -24726
rect 86193 -24770 86249 -24726
rect 86293 -24770 86349 -24726
rect 86393 -24770 86849 -24726
rect 86893 -24770 86949 -24726
rect 86993 -24770 87049 -24726
rect 87093 -24770 87149 -24726
rect 87193 -24770 87249 -24726
rect 87293 -24770 87349 -24726
rect 87393 -24770 87449 -24726
rect 87493 -24770 87549 -24726
rect 87593 -24770 87649 -24726
rect 87693 -24770 87749 -24726
rect 87793 -24770 87849 -24726
rect 87893 -24770 87949 -24726
rect 87993 -24770 88049 -24726
rect 88093 -24770 88149 -24726
rect 88193 -24770 88249 -24726
rect 88293 -24770 88349 -24726
rect 88393 -24770 89254 -24726
rect 79796 -24826 89254 -24770
rect 79796 -24870 80849 -24826
rect 80893 -24870 80949 -24826
rect 80993 -24870 81049 -24826
rect 81093 -24870 81149 -24826
rect 81193 -24870 81249 -24826
rect 81293 -24870 81349 -24826
rect 81393 -24870 81449 -24826
rect 81493 -24870 81549 -24826
rect 81593 -24870 81649 -24826
rect 81693 -24870 81749 -24826
rect 81793 -24870 81849 -24826
rect 81893 -24870 81949 -24826
rect 81993 -24870 82049 -24826
rect 82093 -24870 82149 -24826
rect 82193 -24870 82249 -24826
rect 82293 -24870 82349 -24826
rect 82393 -24870 82849 -24826
rect 82893 -24870 82949 -24826
rect 82993 -24870 83049 -24826
rect 83093 -24870 83149 -24826
rect 83193 -24870 83249 -24826
rect 83293 -24870 83349 -24826
rect 83393 -24870 83449 -24826
rect 83493 -24870 83549 -24826
rect 83593 -24870 83649 -24826
rect 83693 -24870 83749 -24826
rect 83793 -24870 83849 -24826
rect 83893 -24870 83949 -24826
rect 83993 -24870 84049 -24826
rect 84093 -24870 84149 -24826
rect 84193 -24870 84249 -24826
rect 84293 -24870 84349 -24826
rect 84393 -24870 84849 -24826
rect 84893 -24870 84949 -24826
rect 84993 -24870 85049 -24826
rect 85093 -24870 85149 -24826
rect 85193 -24870 85249 -24826
rect 85293 -24870 85349 -24826
rect 85393 -24870 85449 -24826
rect 85493 -24870 85549 -24826
rect 85593 -24870 85649 -24826
rect 85693 -24870 85749 -24826
rect 85793 -24870 85849 -24826
rect 85893 -24870 85949 -24826
rect 85993 -24870 86049 -24826
rect 86093 -24870 86149 -24826
rect 86193 -24870 86249 -24826
rect 86293 -24870 86349 -24826
rect 86393 -24870 86849 -24826
rect 86893 -24870 86949 -24826
rect 86993 -24870 87049 -24826
rect 87093 -24870 87149 -24826
rect 87193 -24870 87249 -24826
rect 87293 -24870 87349 -24826
rect 87393 -24870 87449 -24826
rect 87493 -24870 87549 -24826
rect 87593 -24870 87649 -24826
rect 87693 -24870 87749 -24826
rect 87793 -24870 87849 -24826
rect 87893 -24870 87949 -24826
rect 87993 -24870 88049 -24826
rect 88093 -24870 88149 -24826
rect 88193 -24870 88249 -24826
rect 88293 -24870 88349 -24826
rect 88393 -24870 89254 -24826
rect 79796 -24926 89254 -24870
rect 79796 -24970 80849 -24926
rect 80893 -24970 80949 -24926
rect 80993 -24970 81049 -24926
rect 81093 -24970 81149 -24926
rect 81193 -24970 81249 -24926
rect 81293 -24970 81349 -24926
rect 81393 -24970 81449 -24926
rect 81493 -24970 81549 -24926
rect 81593 -24970 81649 -24926
rect 81693 -24970 81749 -24926
rect 81793 -24970 81849 -24926
rect 81893 -24970 81949 -24926
rect 81993 -24970 82049 -24926
rect 82093 -24970 82149 -24926
rect 82193 -24970 82249 -24926
rect 82293 -24970 82349 -24926
rect 82393 -24970 82849 -24926
rect 82893 -24970 82949 -24926
rect 82993 -24970 83049 -24926
rect 83093 -24970 83149 -24926
rect 83193 -24970 83249 -24926
rect 83293 -24970 83349 -24926
rect 83393 -24970 83449 -24926
rect 83493 -24970 83549 -24926
rect 83593 -24970 83649 -24926
rect 83693 -24970 83749 -24926
rect 83793 -24970 83849 -24926
rect 83893 -24970 83949 -24926
rect 83993 -24970 84049 -24926
rect 84093 -24970 84149 -24926
rect 84193 -24970 84249 -24926
rect 84293 -24970 84349 -24926
rect 84393 -24970 84849 -24926
rect 84893 -24970 84949 -24926
rect 84993 -24970 85049 -24926
rect 85093 -24970 85149 -24926
rect 85193 -24970 85249 -24926
rect 85293 -24970 85349 -24926
rect 85393 -24970 85449 -24926
rect 85493 -24970 85549 -24926
rect 85593 -24970 85649 -24926
rect 85693 -24970 85749 -24926
rect 85793 -24970 85849 -24926
rect 85893 -24970 85949 -24926
rect 85993 -24970 86049 -24926
rect 86093 -24970 86149 -24926
rect 86193 -24970 86249 -24926
rect 86293 -24970 86349 -24926
rect 86393 -24970 86849 -24926
rect 86893 -24970 86949 -24926
rect 86993 -24970 87049 -24926
rect 87093 -24970 87149 -24926
rect 87193 -24970 87249 -24926
rect 87293 -24970 87349 -24926
rect 87393 -24970 87449 -24926
rect 87493 -24970 87549 -24926
rect 87593 -24970 87649 -24926
rect 87693 -24970 87749 -24926
rect 87793 -24970 87849 -24926
rect 87893 -24970 87949 -24926
rect 87993 -24970 88049 -24926
rect 88093 -24970 88149 -24926
rect 88193 -24970 88249 -24926
rect 88293 -24970 88349 -24926
rect 88393 -24970 89254 -24926
rect 79796 -25026 89254 -24970
rect 79796 -25070 80849 -25026
rect 80893 -25070 80949 -25026
rect 80993 -25070 81049 -25026
rect 81093 -25070 81149 -25026
rect 81193 -25070 81249 -25026
rect 81293 -25070 81349 -25026
rect 81393 -25070 81449 -25026
rect 81493 -25070 81549 -25026
rect 81593 -25070 81649 -25026
rect 81693 -25070 81749 -25026
rect 81793 -25070 81849 -25026
rect 81893 -25070 81949 -25026
rect 81993 -25070 82049 -25026
rect 82093 -25070 82149 -25026
rect 82193 -25070 82249 -25026
rect 82293 -25070 82349 -25026
rect 82393 -25070 82849 -25026
rect 82893 -25070 82949 -25026
rect 82993 -25070 83049 -25026
rect 83093 -25070 83149 -25026
rect 83193 -25070 83249 -25026
rect 83293 -25070 83349 -25026
rect 83393 -25070 83449 -25026
rect 83493 -25070 83549 -25026
rect 83593 -25070 83649 -25026
rect 83693 -25070 83749 -25026
rect 83793 -25070 83849 -25026
rect 83893 -25070 83949 -25026
rect 83993 -25070 84049 -25026
rect 84093 -25070 84149 -25026
rect 84193 -25070 84249 -25026
rect 84293 -25070 84349 -25026
rect 84393 -25070 84849 -25026
rect 84893 -25070 84949 -25026
rect 84993 -25070 85049 -25026
rect 85093 -25070 85149 -25026
rect 85193 -25070 85249 -25026
rect 85293 -25070 85349 -25026
rect 85393 -25070 85449 -25026
rect 85493 -25070 85549 -25026
rect 85593 -25070 85649 -25026
rect 85693 -25070 85749 -25026
rect 85793 -25070 85849 -25026
rect 85893 -25070 85949 -25026
rect 85993 -25070 86049 -25026
rect 86093 -25070 86149 -25026
rect 86193 -25070 86249 -25026
rect 86293 -25070 86349 -25026
rect 86393 -25070 86849 -25026
rect 86893 -25070 86949 -25026
rect 86993 -25070 87049 -25026
rect 87093 -25070 87149 -25026
rect 87193 -25070 87249 -25026
rect 87293 -25070 87349 -25026
rect 87393 -25070 87449 -25026
rect 87493 -25070 87549 -25026
rect 87593 -25070 87649 -25026
rect 87693 -25070 87749 -25026
rect 87793 -25070 87849 -25026
rect 87893 -25070 87949 -25026
rect 87993 -25070 88049 -25026
rect 88093 -25070 88149 -25026
rect 88193 -25070 88249 -25026
rect 88293 -25070 88349 -25026
rect 88393 -25070 89254 -25026
rect 79796 -25126 89254 -25070
rect 79796 -25170 80849 -25126
rect 80893 -25170 80949 -25126
rect 80993 -25170 81049 -25126
rect 81093 -25170 81149 -25126
rect 81193 -25170 81249 -25126
rect 81293 -25170 81349 -25126
rect 81393 -25170 81449 -25126
rect 81493 -25170 81549 -25126
rect 81593 -25170 81649 -25126
rect 81693 -25170 81749 -25126
rect 81793 -25170 81849 -25126
rect 81893 -25170 81949 -25126
rect 81993 -25170 82049 -25126
rect 82093 -25170 82149 -25126
rect 82193 -25170 82249 -25126
rect 82293 -25170 82349 -25126
rect 82393 -25170 82849 -25126
rect 82893 -25170 82949 -25126
rect 82993 -25170 83049 -25126
rect 83093 -25170 83149 -25126
rect 83193 -25170 83249 -25126
rect 83293 -25170 83349 -25126
rect 83393 -25170 83449 -25126
rect 83493 -25170 83549 -25126
rect 83593 -25170 83649 -25126
rect 83693 -25170 83749 -25126
rect 83793 -25170 83849 -25126
rect 83893 -25170 83949 -25126
rect 83993 -25170 84049 -25126
rect 84093 -25170 84149 -25126
rect 84193 -25170 84249 -25126
rect 84293 -25170 84349 -25126
rect 84393 -25170 84849 -25126
rect 84893 -25170 84949 -25126
rect 84993 -25170 85049 -25126
rect 85093 -25170 85149 -25126
rect 85193 -25170 85249 -25126
rect 85293 -25170 85349 -25126
rect 85393 -25170 85449 -25126
rect 85493 -25170 85549 -25126
rect 85593 -25170 85649 -25126
rect 85693 -25170 85749 -25126
rect 85793 -25170 85849 -25126
rect 85893 -25170 85949 -25126
rect 85993 -25170 86049 -25126
rect 86093 -25170 86149 -25126
rect 86193 -25170 86249 -25126
rect 86293 -25170 86349 -25126
rect 86393 -25170 86849 -25126
rect 86893 -25170 86949 -25126
rect 86993 -25170 87049 -25126
rect 87093 -25170 87149 -25126
rect 87193 -25170 87249 -25126
rect 87293 -25170 87349 -25126
rect 87393 -25170 87449 -25126
rect 87493 -25170 87549 -25126
rect 87593 -25170 87649 -25126
rect 87693 -25170 87749 -25126
rect 87793 -25170 87849 -25126
rect 87893 -25170 87949 -25126
rect 87993 -25170 88049 -25126
rect 88093 -25170 88149 -25126
rect 88193 -25170 88249 -25126
rect 88293 -25170 88349 -25126
rect 88393 -25170 89254 -25126
rect 79796 -25226 89254 -25170
rect 79796 -25270 80849 -25226
rect 80893 -25270 80949 -25226
rect 80993 -25270 81049 -25226
rect 81093 -25270 81149 -25226
rect 81193 -25270 81249 -25226
rect 81293 -25270 81349 -25226
rect 81393 -25270 81449 -25226
rect 81493 -25270 81549 -25226
rect 81593 -25270 81649 -25226
rect 81693 -25270 81749 -25226
rect 81793 -25270 81849 -25226
rect 81893 -25270 81949 -25226
rect 81993 -25270 82049 -25226
rect 82093 -25270 82149 -25226
rect 82193 -25270 82249 -25226
rect 82293 -25270 82349 -25226
rect 82393 -25270 82849 -25226
rect 82893 -25270 82949 -25226
rect 82993 -25270 83049 -25226
rect 83093 -25270 83149 -25226
rect 83193 -25270 83249 -25226
rect 83293 -25270 83349 -25226
rect 83393 -25270 83449 -25226
rect 83493 -25270 83549 -25226
rect 83593 -25270 83649 -25226
rect 83693 -25270 83749 -25226
rect 83793 -25270 83849 -25226
rect 83893 -25270 83949 -25226
rect 83993 -25270 84049 -25226
rect 84093 -25270 84149 -25226
rect 84193 -25270 84249 -25226
rect 84293 -25270 84349 -25226
rect 84393 -25270 84849 -25226
rect 84893 -25270 84949 -25226
rect 84993 -25270 85049 -25226
rect 85093 -25270 85149 -25226
rect 85193 -25270 85249 -25226
rect 85293 -25270 85349 -25226
rect 85393 -25270 85449 -25226
rect 85493 -25270 85549 -25226
rect 85593 -25270 85649 -25226
rect 85693 -25270 85749 -25226
rect 85793 -25270 85849 -25226
rect 85893 -25270 85949 -25226
rect 85993 -25270 86049 -25226
rect 86093 -25270 86149 -25226
rect 86193 -25270 86249 -25226
rect 86293 -25270 86349 -25226
rect 86393 -25270 86849 -25226
rect 86893 -25270 86949 -25226
rect 86993 -25270 87049 -25226
rect 87093 -25270 87149 -25226
rect 87193 -25270 87249 -25226
rect 87293 -25270 87349 -25226
rect 87393 -25270 87449 -25226
rect 87493 -25270 87549 -25226
rect 87593 -25270 87649 -25226
rect 87693 -25270 87749 -25226
rect 87793 -25270 87849 -25226
rect 87893 -25270 87949 -25226
rect 87993 -25270 88049 -25226
rect 88093 -25270 88149 -25226
rect 88193 -25270 88249 -25226
rect 88293 -25270 88349 -25226
rect 88393 -25270 89254 -25226
rect 79796 -25326 89254 -25270
rect 79796 -25370 80849 -25326
rect 80893 -25370 80949 -25326
rect 80993 -25370 81049 -25326
rect 81093 -25370 81149 -25326
rect 81193 -25370 81249 -25326
rect 81293 -25370 81349 -25326
rect 81393 -25370 81449 -25326
rect 81493 -25370 81549 -25326
rect 81593 -25370 81649 -25326
rect 81693 -25370 81749 -25326
rect 81793 -25370 81849 -25326
rect 81893 -25370 81949 -25326
rect 81993 -25370 82049 -25326
rect 82093 -25370 82149 -25326
rect 82193 -25370 82249 -25326
rect 82293 -25370 82349 -25326
rect 82393 -25370 82849 -25326
rect 82893 -25370 82949 -25326
rect 82993 -25370 83049 -25326
rect 83093 -25370 83149 -25326
rect 83193 -25370 83249 -25326
rect 83293 -25370 83349 -25326
rect 83393 -25370 83449 -25326
rect 83493 -25370 83549 -25326
rect 83593 -25370 83649 -25326
rect 83693 -25370 83749 -25326
rect 83793 -25370 83849 -25326
rect 83893 -25370 83949 -25326
rect 83993 -25370 84049 -25326
rect 84093 -25370 84149 -25326
rect 84193 -25370 84249 -25326
rect 84293 -25370 84349 -25326
rect 84393 -25370 84849 -25326
rect 84893 -25370 84949 -25326
rect 84993 -25370 85049 -25326
rect 85093 -25370 85149 -25326
rect 85193 -25370 85249 -25326
rect 85293 -25370 85349 -25326
rect 85393 -25370 85449 -25326
rect 85493 -25370 85549 -25326
rect 85593 -25370 85649 -25326
rect 85693 -25370 85749 -25326
rect 85793 -25370 85849 -25326
rect 85893 -25370 85949 -25326
rect 85993 -25370 86049 -25326
rect 86093 -25370 86149 -25326
rect 86193 -25370 86249 -25326
rect 86293 -25370 86349 -25326
rect 86393 -25370 86849 -25326
rect 86893 -25370 86949 -25326
rect 86993 -25370 87049 -25326
rect 87093 -25370 87149 -25326
rect 87193 -25370 87249 -25326
rect 87293 -25370 87349 -25326
rect 87393 -25370 87449 -25326
rect 87493 -25370 87549 -25326
rect 87593 -25370 87649 -25326
rect 87693 -25370 87749 -25326
rect 87793 -25370 87849 -25326
rect 87893 -25370 87949 -25326
rect 87993 -25370 88049 -25326
rect 88093 -25370 88149 -25326
rect 88193 -25370 88249 -25326
rect 88293 -25370 88349 -25326
rect 88393 -25370 89254 -25326
rect 79796 -25426 89254 -25370
rect 79796 -25470 80849 -25426
rect 80893 -25470 80949 -25426
rect 80993 -25470 81049 -25426
rect 81093 -25470 81149 -25426
rect 81193 -25470 81249 -25426
rect 81293 -25470 81349 -25426
rect 81393 -25470 81449 -25426
rect 81493 -25470 81549 -25426
rect 81593 -25470 81649 -25426
rect 81693 -25470 81749 -25426
rect 81793 -25470 81849 -25426
rect 81893 -25470 81949 -25426
rect 81993 -25470 82049 -25426
rect 82093 -25470 82149 -25426
rect 82193 -25470 82249 -25426
rect 82293 -25470 82349 -25426
rect 82393 -25470 82849 -25426
rect 82893 -25470 82949 -25426
rect 82993 -25470 83049 -25426
rect 83093 -25470 83149 -25426
rect 83193 -25470 83249 -25426
rect 83293 -25470 83349 -25426
rect 83393 -25470 83449 -25426
rect 83493 -25470 83549 -25426
rect 83593 -25470 83649 -25426
rect 83693 -25470 83749 -25426
rect 83793 -25470 83849 -25426
rect 83893 -25470 83949 -25426
rect 83993 -25470 84049 -25426
rect 84093 -25470 84149 -25426
rect 84193 -25470 84249 -25426
rect 84293 -25470 84349 -25426
rect 84393 -25470 84849 -25426
rect 84893 -25470 84949 -25426
rect 84993 -25470 85049 -25426
rect 85093 -25470 85149 -25426
rect 85193 -25470 85249 -25426
rect 85293 -25470 85349 -25426
rect 85393 -25470 85449 -25426
rect 85493 -25470 85549 -25426
rect 85593 -25470 85649 -25426
rect 85693 -25470 85749 -25426
rect 85793 -25470 85849 -25426
rect 85893 -25470 85949 -25426
rect 85993 -25470 86049 -25426
rect 86093 -25470 86149 -25426
rect 86193 -25470 86249 -25426
rect 86293 -25470 86349 -25426
rect 86393 -25470 86849 -25426
rect 86893 -25470 86949 -25426
rect 86993 -25470 87049 -25426
rect 87093 -25470 87149 -25426
rect 87193 -25470 87249 -25426
rect 87293 -25470 87349 -25426
rect 87393 -25470 87449 -25426
rect 87493 -25470 87549 -25426
rect 87593 -25470 87649 -25426
rect 87693 -25470 87749 -25426
rect 87793 -25470 87849 -25426
rect 87893 -25470 87949 -25426
rect 87993 -25470 88049 -25426
rect 88093 -25470 88149 -25426
rect 88193 -25470 88249 -25426
rect 88293 -25470 88349 -25426
rect 88393 -25470 89254 -25426
rect 79796 -25526 89254 -25470
rect 79796 -25570 80849 -25526
rect 80893 -25570 80949 -25526
rect 80993 -25570 81049 -25526
rect 81093 -25570 81149 -25526
rect 81193 -25570 81249 -25526
rect 81293 -25570 81349 -25526
rect 81393 -25570 81449 -25526
rect 81493 -25570 81549 -25526
rect 81593 -25570 81649 -25526
rect 81693 -25570 81749 -25526
rect 81793 -25570 81849 -25526
rect 81893 -25570 81949 -25526
rect 81993 -25570 82049 -25526
rect 82093 -25570 82149 -25526
rect 82193 -25570 82249 -25526
rect 82293 -25570 82349 -25526
rect 82393 -25570 82849 -25526
rect 82893 -25570 82949 -25526
rect 82993 -25570 83049 -25526
rect 83093 -25570 83149 -25526
rect 83193 -25570 83249 -25526
rect 83293 -25570 83349 -25526
rect 83393 -25570 83449 -25526
rect 83493 -25570 83549 -25526
rect 83593 -25570 83649 -25526
rect 83693 -25570 83749 -25526
rect 83793 -25570 83849 -25526
rect 83893 -25570 83949 -25526
rect 83993 -25570 84049 -25526
rect 84093 -25570 84149 -25526
rect 84193 -25570 84249 -25526
rect 84293 -25570 84349 -25526
rect 84393 -25570 84849 -25526
rect 84893 -25570 84949 -25526
rect 84993 -25570 85049 -25526
rect 85093 -25570 85149 -25526
rect 85193 -25570 85249 -25526
rect 85293 -25570 85349 -25526
rect 85393 -25570 85449 -25526
rect 85493 -25570 85549 -25526
rect 85593 -25570 85649 -25526
rect 85693 -25570 85749 -25526
rect 85793 -25570 85849 -25526
rect 85893 -25570 85949 -25526
rect 85993 -25570 86049 -25526
rect 86093 -25570 86149 -25526
rect 86193 -25570 86249 -25526
rect 86293 -25570 86349 -25526
rect 86393 -25570 86849 -25526
rect 86893 -25570 86949 -25526
rect 86993 -25570 87049 -25526
rect 87093 -25570 87149 -25526
rect 87193 -25570 87249 -25526
rect 87293 -25570 87349 -25526
rect 87393 -25570 87449 -25526
rect 87493 -25570 87549 -25526
rect 87593 -25570 87649 -25526
rect 87693 -25570 87749 -25526
rect 87793 -25570 87849 -25526
rect 87893 -25570 87949 -25526
rect 87993 -25570 88049 -25526
rect 88093 -25570 88149 -25526
rect 88193 -25570 88249 -25526
rect 88293 -25570 88349 -25526
rect 88393 -25570 89254 -25526
rect 79796 -80455 89254 -25570
rect 108496 -24195 117196 -23015
rect 108496 -24239 109104 -24195
rect 109148 -24239 109204 -24195
rect 109248 -24239 109304 -24195
rect 109348 -24239 109404 -24195
rect 109448 -24239 109504 -24195
rect 109548 -24239 109604 -24195
rect 109648 -24239 109704 -24195
rect 109748 -24239 109804 -24195
rect 109848 -24239 109904 -24195
rect 109948 -24239 110004 -24195
rect 110048 -24239 110104 -24195
rect 110148 -24239 110204 -24195
rect 110248 -24239 110304 -24195
rect 110348 -24239 110404 -24195
rect 110448 -24239 110504 -24195
rect 110548 -24239 110604 -24195
rect 110648 -24239 111104 -24195
rect 111148 -24239 111204 -24195
rect 111248 -24239 111304 -24195
rect 111348 -24239 111404 -24195
rect 111448 -24239 111504 -24195
rect 111548 -24239 111604 -24195
rect 111648 -24239 111704 -24195
rect 111748 -24239 111804 -24195
rect 111848 -24239 111904 -24195
rect 111948 -24239 112004 -24195
rect 112048 -24239 112104 -24195
rect 112148 -24239 112204 -24195
rect 112248 -24239 112304 -24195
rect 112348 -24239 112404 -24195
rect 112448 -24239 112504 -24195
rect 112548 -24239 112604 -24195
rect 112648 -24239 113104 -24195
rect 113148 -24239 113204 -24195
rect 113248 -24239 113304 -24195
rect 113348 -24239 113404 -24195
rect 113448 -24239 113504 -24195
rect 113548 -24239 113604 -24195
rect 113648 -24239 113704 -24195
rect 113748 -24239 113804 -24195
rect 113848 -24239 113904 -24195
rect 113948 -24239 114004 -24195
rect 114048 -24239 114104 -24195
rect 114148 -24239 114204 -24195
rect 114248 -24239 114304 -24195
rect 114348 -24239 114404 -24195
rect 114448 -24239 114504 -24195
rect 114548 -24239 114604 -24195
rect 114648 -24239 115104 -24195
rect 115148 -24239 115204 -24195
rect 115248 -24239 115304 -24195
rect 115348 -24239 115404 -24195
rect 115448 -24239 115504 -24195
rect 115548 -24239 115604 -24195
rect 115648 -24239 115704 -24195
rect 115748 -24239 115804 -24195
rect 115848 -24239 115904 -24195
rect 115948 -24239 116004 -24195
rect 116048 -24239 116104 -24195
rect 116148 -24239 116204 -24195
rect 116248 -24239 116304 -24195
rect 116348 -24239 116404 -24195
rect 116448 -24239 116504 -24195
rect 116548 -24239 116604 -24195
rect 116648 -24239 117196 -24195
rect 108496 -24295 117196 -24239
rect 108496 -24339 109104 -24295
rect 109148 -24339 109204 -24295
rect 109248 -24339 109304 -24295
rect 109348 -24339 109404 -24295
rect 109448 -24339 109504 -24295
rect 109548 -24339 109604 -24295
rect 109648 -24339 109704 -24295
rect 109748 -24339 109804 -24295
rect 109848 -24339 109904 -24295
rect 109948 -24339 110004 -24295
rect 110048 -24339 110104 -24295
rect 110148 -24339 110204 -24295
rect 110248 -24339 110304 -24295
rect 110348 -24339 110404 -24295
rect 110448 -24339 110504 -24295
rect 110548 -24339 110604 -24295
rect 110648 -24339 111104 -24295
rect 111148 -24339 111204 -24295
rect 111248 -24339 111304 -24295
rect 111348 -24339 111404 -24295
rect 111448 -24339 111504 -24295
rect 111548 -24339 111604 -24295
rect 111648 -24339 111704 -24295
rect 111748 -24339 111804 -24295
rect 111848 -24339 111904 -24295
rect 111948 -24339 112004 -24295
rect 112048 -24339 112104 -24295
rect 112148 -24339 112204 -24295
rect 112248 -24339 112304 -24295
rect 112348 -24339 112404 -24295
rect 112448 -24339 112504 -24295
rect 112548 -24339 112604 -24295
rect 112648 -24339 113104 -24295
rect 113148 -24339 113204 -24295
rect 113248 -24339 113304 -24295
rect 113348 -24339 113404 -24295
rect 113448 -24339 113504 -24295
rect 113548 -24339 113604 -24295
rect 113648 -24339 113704 -24295
rect 113748 -24339 113804 -24295
rect 113848 -24339 113904 -24295
rect 113948 -24339 114004 -24295
rect 114048 -24339 114104 -24295
rect 114148 -24339 114204 -24295
rect 114248 -24339 114304 -24295
rect 114348 -24339 114404 -24295
rect 114448 -24339 114504 -24295
rect 114548 -24339 114604 -24295
rect 114648 -24339 115104 -24295
rect 115148 -24339 115204 -24295
rect 115248 -24339 115304 -24295
rect 115348 -24339 115404 -24295
rect 115448 -24339 115504 -24295
rect 115548 -24339 115604 -24295
rect 115648 -24339 115704 -24295
rect 115748 -24339 115804 -24295
rect 115848 -24339 115904 -24295
rect 115948 -24339 116004 -24295
rect 116048 -24339 116104 -24295
rect 116148 -24339 116204 -24295
rect 116248 -24339 116304 -24295
rect 116348 -24339 116404 -24295
rect 116448 -24339 116504 -24295
rect 116548 -24339 116604 -24295
rect 116648 -24339 117196 -24295
rect 108496 -24395 117196 -24339
rect 108496 -24439 109104 -24395
rect 109148 -24439 109204 -24395
rect 109248 -24439 109304 -24395
rect 109348 -24439 109404 -24395
rect 109448 -24439 109504 -24395
rect 109548 -24439 109604 -24395
rect 109648 -24439 109704 -24395
rect 109748 -24439 109804 -24395
rect 109848 -24439 109904 -24395
rect 109948 -24439 110004 -24395
rect 110048 -24439 110104 -24395
rect 110148 -24439 110204 -24395
rect 110248 -24439 110304 -24395
rect 110348 -24439 110404 -24395
rect 110448 -24439 110504 -24395
rect 110548 -24439 110604 -24395
rect 110648 -24439 111104 -24395
rect 111148 -24439 111204 -24395
rect 111248 -24439 111304 -24395
rect 111348 -24439 111404 -24395
rect 111448 -24439 111504 -24395
rect 111548 -24439 111604 -24395
rect 111648 -24439 111704 -24395
rect 111748 -24439 111804 -24395
rect 111848 -24439 111904 -24395
rect 111948 -24439 112004 -24395
rect 112048 -24439 112104 -24395
rect 112148 -24439 112204 -24395
rect 112248 -24439 112304 -24395
rect 112348 -24439 112404 -24395
rect 112448 -24439 112504 -24395
rect 112548 -24439 112604 -24395
rect 112648 -24439 113104 -24395
rect 113148 -24439 113204 -24395
rect 113248 -24439 113304 -24395
rect 113348 -24439 113404 -24395
rect 113448 -24439 113504 -24395
rect 113548 -24439 113604 -24395
rect 113648 -24439 113704 -24395
rect 113748 -24439 113804 -24395
rect 113848 -24439 113904 -24395
rect 113948 -24439 114004 -24395
rect 114048 -24439 114104 -24395
rect 114148 -24439 114204 -24395
rect 114248 -24439 114304 -24395
rect 114348 -24439 114404 -24395
rect 114448 -24439 114504 -24395
rect 114548 -24439 114604 -24395
rect 114648 -24439 115104 -24395
rect 115148 -24439 115204 -24395
rect 115248 -24439 115304 -24395
rect 115348 -24439 115404 -24395
rect 115448 -24439 115504 -24395
rect 115548 -24439 115604 -24395
rect 115648 -24439 115704 -24395
rect 115748 -24439 115804 -24395
rect 115848 -24439 115904 -24395
rect 115948 -24439 116004 -24395
rect 116048 -24439 116104 -24395
rect 116148 -24439 116204 -24395
rect 116248 -24439 116304 -24395
rect 116348 -24439 116404 -24395
rect 116448 -24439 116504 -24395
rect 116548 -24439 116604 -24395
rect 116648 -24439 117196 -24395
rect 108496 -24495 117196 -24439
rect 108496 -24539 109104 -24495
rect 109148 -24539 109204 -24495
rect 109248 -24539 109304 -24495
rect 109348 -24539 109404 -24495
rect 109448 -24539 109504 -24495
rect 109548 -24539 109604 -24495
rect 109648 -24539 109704 -24495
rect 109748 -24539 109804 -24495
rect 109848 -24539 109904 -24495
rect 109948 -24539 110004 -24495
rect 110048 -24539 110104 -24495
rect 110148 -24539 110204 -24495
rect 110248 -24539 110304 -24495
rect 110348 -24539 110404 -24495
rect 110448 -24539 110504 -24495
rect 110548 -24539 110604 -24495
rect 110648 -24539 111104 -24495
rect 111148 -24539 111204 -24495
rect 111248 -24539 111304 -24495
rect 111348 -24539 111404 -24495
rect 111448 -24539 111504 -24495
rect 111548 -24539 111604 -24495
rect 111648 -24539 111704 -24495
rect 111748 -24539 111804 -24495
rect 111848 -24539 111904 -24495
rect 111948 -24539 112004 -24495
rect 112048 -24539 112104 -24495
rect 112148 -24539 112204 -24495
rect 112248 -24539 112304 -24495
rect 112348 -24539 112404 -24495
rect 112448 -24539 112504 -24495
rect 112548 -24539 112604 -24495
rect 112648 -24539 113104 -24495
rect 113148 -24539 113204 -24495
rect 113248 -24539 113304 -24495
rect 113348 -24539 113404 -24495
rect 113448 -24539 113504 -24495
rect 113548 -24539 113604 -24495
rect 113648 -24539 113704 -24495
rect 113748 -24539 113804 -24495
rect 113848 -24539 113904 -24495
rect 113948 -24539 114004 -24495
rect 114048 -24539 114104 -24495
rect 114148 -24539 114204 -24495
rect 114248 -24539 114304 -24495
rect 114348 -24539 114404 -24495
rect 114448 -24539 114504 -24495
rect 114548 -24539 114604 -24495
rect 114648 -24539 115104 -24495
rect 115148 -24539 115204 -24495
rect 115248 -24539 115304 -24495
rect 115348 -24539 115404 -24495
rect 115448 -24539 115504 -24495
rect 115548 -24539 115604 -24495
rect 115648 -24539 115704 -24495
rect 115748 -24539 115804 -24495
rect 115848 -24539 115904 -24495
rect 115948 -24539 116004 -24495
rect 116048 -24539 116104 -24495
rect 116148 -24539 116204 -24495
rect 116248 -24539 116304 -24495
rect 116348 -24539 116404 -24495
rect 116448 -24539 116504 -24495
rect 116548 -24539 116604 -24495
rect 116648 -24539 117196 -24495
rect 108496 -24595 117196 -24539
rect 108496 -24639 109104 -24595
rect 109148 -24639 109204 -24595
rect 109248 -24639 109304 -24595
rect 109348 -24639 109404 -24595
rect 109448 -24639 109504 -24595
rect 109548 -24639 109604 -24595
rect 109648 -24639 109704 -24595
rect 109748 -24639 109804 -24595
rect 109848 -24639 109904 -24595
rect 109948 -24639 110004 -24595
rect 110048 -24639 110104 -24595
rect 110148 -24639 110204 -24595
rect 110248 -24639 110304 -24595
rect 110348 -24639 110404 -24595
rect 110448 -24639 110504 -24595
rect 110548 -24639 110604 -24595
rect 110648 -24639 111104 -24595
rect 111148 -24639 111204 -24595
rect 111248 -24639 111304 -24595
rect 111348 -24639 111404 -24595
rect 111448 -24639 111504 -24595
rect 111548 -24639 111604 -24595
rect 111648 -24639 111704 -24595
rect 111748 -24639 111804 -24595
rect 111848 -24639 111904 -24595
rect 111948 -24639 112004 -24595
rect 112048 -24639 112104 -24595
rect 112148 -24639 112204 -24595
rect 112248 -24639 112304 -24595
rect 112348 -24639 112404 -24595
rect 112448 -24639 112504 -24595
rect 112548 -24639 112604 -24595
rect 112648 -24639 113104 -24595
rect 113148 -24639 113204 -24595
rect 113248 -24639 113304 -24595
rect 113348 -24639 113404 -24595
rect 113448 -24639 113504 -24595
rect 113548 -24639 113604 -24595
rect 113648 -24639 113704 -24595
rect 113748 -24639 113804 -24595
rect 113848 -24639 113904 -24595
rect 113948 -24639 114004 -24595
rect 114048 -24639 114104 -24595
rect 114148 -24639 114204 -24595
rect 114248 -24639 114304 -24595
rect 114348 -24639 114404 -24595
rect 114448 -24639 114504 -24595
rect 114548 -24639 114604 -24595
rect 114648 -24639 115104 -24595
rect 115148 -24639 115204 -24595
rect 115248 -24639 115304 -24595
rect 115348 -24639 115404 -24595
rect 115448 -24639 115504 -24595
rect 115548 -24639 115604 -24595
rect 115648 -24639 115704 -24595
rect 115748 -24639 115804 -24595
rect 115848 -24639 115904 -24595
rect 115948 -24639 116004 -24595
rect 116048 -24639 116104 -24595
rect 116148 -24639 116204 -24595
rect 116248 -24639 116304 -24595
rect 116348 -24639 116404 -24595
rect 116448 -24639 116504 -24595
rect 116548 -24639 116604 -24595
rect 116648 -24639 117196 -24595
rect 108496 -24695 117196 -24639
rect 108496 -24739 109104 -24695
rect 109148 -24739 109204 -24695
rect 109248 -24739 109304 -24695
rect 109348 -24739 109404 -24695
rect 109448 -24739 109504 -24695
rect 109548 -24739 109604 -24695
rect 109648 -24739 109704 -24695
rect 109748 -24739 109804 -24695
rect 109848 -24739 109904 -24695
rect 109948 -24739 110004 -24695
rect 110048 -24739 110104 -24695
rect 110148 -24739 110204 -24695
rect 110248 -24739 110304 -24695
rect 110348 -24739 110404 -24695
rect 110448 -24739 110504 -24695
rect 110548 -24739 110604 -24695
rect 110648 -24739 111104 -24695
rect 111148 -24739 111204 -24695
rect 111248 -24739 111304 -24695
rect 111348 -24739 111404 -24695
rect 111448 -24739 111504 -24695
rect 111548 -24739 111604 -24695
rect 111648 -24739 111704 -24695
rect 111748 -24739 111804 -24695
rect 111848 -24739 111904 -24695
rect 111948 -24739 112004 -24695
rect 112048 -24739 112104 -24695
rect 112148 -24739 112204 -24695
rect 112248 -24739 112304 -24695
rect 112348 -24739 112404 -24695
rect 112448 -24739 112504 -24695
rect 112548 -24739 112604 -24695
rect 112648 -24739 113104 -24695
rect 113148 -24739 113204 -24695
rect 113248 -24739 113304 -24695
rect 113348 -24739 113404 -24695
rect 113448 -24739 113504 -24695
rect 113548 -24739 113604 -24695
rect 113648 -24739 113704 -24695
rect 113748 -24739 113804 -24695
rect 113848 -24739 113904 -24695
rect 113948 -24739 114004 -24695
rect 114048 -24739 114104 -24695
rect 114148 -24739 114204 -24695
rect 114248 -24739 114304 -24695
rect 114348 -24739 114404 -24695
rect 114448 -24739 114504 -24695
rect 114548 -24739 114604 -24695
rect 114648 -24739 115104 -24695
rect 115148 -24739 115204 -24695
rect 115248 -24739 115304 -24695
rect 115348 -24739 115404 -24695
rect 115448 -24739 115504 -24695
rect 115548 -24739 115604 -24695
rect 115648 -24739 115704 -24695
rect 115748 -24739 115804 -24695
rect 115848 -24739 115904 -24695
rect 115948 -24739 116004 -24695
rect 116048 -24739 116104 -24695
rect 116148 -24739 116204 -24695
rect 116248 -24739 116304 -24695
rect 116348 -24739 116404 -24695
rect 116448 -24739 116504 -24695
rect 116548 -24739 116604 -24695
rect 116648 -24739 117196 -24695
rect 108496 -24795 117196 -24739
rect 108496 -24839 109104 -24795
rect 109148 -24839 109204 -24795
rect 109248 -24839 109304 -24795
rect 109348 -24839 109404 -24795
rect 109448 -24839 109504 -24795
rect 109548 -24839 109604 -24795
rect 109648 -24839 109704 -24795
rect 109748 -24839 109804 -24795
rect 109848 -24839 109904 -24795
rect 109948 -24839 110004 -24795
rect 110048 -24839 110104 -24795
rect 110148 -24839 110204 -24795
rect 110248 -24839 110304 -24795
rect 110348 -24839 110404 -24795
rect 110448 -24839 110504 -24795
rect 110548 -24839 110604 -24795
rect 110648 -24839 111104 -24795
rect 111148 -24839 111204 -24795
rect 111248 -24839 111304 -24795
rect 111348 -24839 111404 -24795
rect 111448 -24839 111504 -24795
rect 111548 -24839 111604 -24795
rect 111648 -24839 111704 -24795
rect 111748 -24839 111804 -24795
rect 111848 -24839 111904 -24795
rect 111948 -24839 112004 -24795
rect 112048 -24839 112104 -24795
rect 112148 -24839 112204 -24795
rect 112248 -24839 112304 -24795
rect 112348 -24839 112404 -24795
rect 112448 -24839 112504 -24795
rect 112548 -24839 112604 -24795
rect 112648 -24839 113104 -24795
rect 113148 -24839 113204 -24795
rect 113248 -24839 113304 -24795
rect 113348 -24839 113404 -24795
rect 113448 -24839 113504 -24795
rect 113548 -24839 113604 -24795
rect 113648 -24839 113704 -24795
rect 113748 -24839 113804 -24795
rect 113848 -24839 113904 -24795
rect 113948 -24839 114004 -24795
rect 114048 -24839 114104 -24795
rect 114148 -24839 114204 -24795
rect 114248 -24839 114304 -24795
rect 114348 -24839 114404 -24795
rect 114448 -24839 114504 -24795
rect 114548 -24839 114604 -24795
rect 114648 -24839 115104 -24795
rect 115148 -24839 115204 -24795
rect 115248 -24839 115304 -24795
rect 115348 -24839 115404 -24795
rect 115448 -24839 115504 -24795
rect 115548 -24839 115604 -24795
rect 115648 -24839 115704 -24795
rect 115748 -24839 115804 -24795
rect 115848 -24839 115904 -24795
rect 115948 -24839 116004 -24795
rect 116048 -24839 116104 -24795
rect 116148 -24839 116204 -24795
rect 116248 -24839 116304 -24795
rect 116348 -24839 116404 -24795
rect 116448 -24839 116504 -24795
rect 116548 -24839 116604 -24795
rect 116648 -24839 117196 -24795
rect 108496 -24895 117196 -24839
rect 108496 -24939 109104 -24895
rect 109148 -24939 109204 -24895
rect 109248 -24939 109304 -24895
rect 109348 -24939 109404 -24895
rect 109448 -24939 109504 -24895
rect 109548 -24939 109604 -24895
rect 109648 -24939 109704 -24895
rect 109748 -24939 109804 -24895
rect 109848 -24939 109904 -24895
rect 109948 -24939 110004 -24895
rect 110048 -24939 110104 -24895
rect 110148 -24939 110204 -24895
rect 110248 -24939 110304 -24895
rect 110348 -24939 110404 -24895
rect 110448 -24939 110504 -24895
rect 110548 -24939 110604 -24895
rect 110648 -24939 111104 -24895
rect 111148 -24939 111204 -24895
rect 111248 -24939 111304 -24895
rect 111348 -24939 111404 -24895
rect 111448 -24939 111504 -24895
rect 111548 -24939 111604 -24895
rect 111648 -24939 111704 -24895
rect 111748 -24939 111804 -24895
rect 111848 -24939 111904 -24895
rect 111948 -24939 112004 -24895
rect 112048 -24939 112104 -24895
rect 112148 -24939 112204 -24895
rect 112248 -24939 112304 -24895
rect 112348 -24939 112404 -24895
rect 112448 -24939 112504 -24895
rect 112548 -24939 112604 -24895
rect 112648 -24939 113104 -24895
rect 113148 -24939 113204 -24895
rect 113248 -24939 113304 -24895
rect 113348 -24939 113404 -24895
rect 113448 -24939 113504 -24895
rect 113548 -24939 113604 -24895
rect 113648 -24939 113704 -24895
rect 113748 -24939 113804 -24895
rect 113848 -24939 113904 -24895
rect 113948 -24939 114004 -24895
rect 114048 -24939 114104 -24895
rect 114148 -24939 114204 -24895
rect 114248 -24939 114304 -24895
rect 114348 -24939 114404 -24895
rect 114448 -24939 114504 -24895
rect 114548 -24939 114604 -24895
rect 114648 -24939 115104 -24895
rect 115148 -24939 115204 -24895
rect 115248 -24939 115304 -24895
rect 115348 -24939 115404 -24895
rect 115448 -24939 115504 -24895
rect 115548 -24939 115604 -24895
rect 115648 -24939 115704 -24895
rect 115748 -24939 115804 -24895
rect 115848 -24939 115904 -24895
rect 115948 -24939 116004 -24895
rect 116048 -24939 116104 -24895
rect 116148 -24939 116204 -24895
rect 116248 -24939 116304 -24895
rect 116348 -24939 116404 -24895
rect 116448 -24939 116504 -24895
rect 116548 -24939 116604 -24895
rect 116648 -24939 117196 -24895
rect 108496 -24995 117196 -24939
rect 108496 -25039 109104 -24995
rect 109148 -25039 109204 -24995
rect 109248 -25039 109304 -24995
rect 109348 -25039 109404 -24995
rect 109448 -25039 109504 -24995
rect 109548 -25039 109604 -24995
rect 109648 -25039 109704 -24995
rect 109748 -25039 109804 -24995
rect 109848 -25039 109904 -24995
rect 109948 -25039 110004 -24995
rect 110048 -25039 110104 -24995
rect 110148 -25039 110204 -24995
rect 110248 -25039 110304 -24995
rect 110348 -25039 110404 -24995
rect 110448 -25039 110504 -24995
rect 110548 -25039 110604 -24995
rect 110648 -25039 111104 -24995
rect 111148 -25039 111204 -24995
rect 111248 -25039 111304 -24995
rect 111348 -25039 111404 -24995
rect 111448 -25039 111504 -24995
rect 111548 -25039 111604 -24995
rect 111648 -25039 111704 -24995
rect 111748 -25039 111804 -24995
rect 111848 -25039 111904 -24995
rect 111948 -25039 112004 -24995
rect 112048 -25039 112104 -24995
rect 112148 -25039 112204 -24995
rect 112248 -25039 112304 -24995
rect 112348 -25039 112404 -24995
rect 112448 -25039 112504 -24995
rect 112548 -25039 112604 -24995
rect 112648 -25039 113104 -24995
rect 113148 -25039 113204 -24995
rect 113248 -25039 113304 -24995
rect 113348 -25039 113404 -24995
rect 113448 -25039 113504 -24995
rect 113548 -25039 113604 -24995
rect 113648 -25039 113704 -24995
rect 113748 -25039 113804 -24995
rect 113848 -25039 113904 -24995
rect 113948 -25039 114004 -24995
rect 114048 -25039 114104 -24995
rect 114148 -25039 114204 -24995
rect 114248 -25039 114304 -24995
rect 114348 -25039 114404 -24995
rect 114448 -25039 114504 -24995
rect 114548 -25039 114604 -24995
rect 114648 -25039 115104 -24995
rect 115148 -25039 115204 -24995
rect 115248 -25039 115304 -24995
rect 115348 -25039 115404 -24995
rect 115448 -25039 115504 -24995
rect 115548 -25039 115604 -24995
rect 115648 -25039 115704 -24995
rect 115748 -25039 115804 -24995
rect 115848 -25039 115904 -24995
rect 115948 -25039 116004 -24995
rect 116048 -25039 116104 -24995
rect 116148 -25039 116204 -24995
rect 116248 -25039 116304 -24995
rect 116348 -25039 116404 -24995
rect 116448 -25039 116504 -24995
rect 116548 -25039 116604 -24995
rect 116648 -25039 117196 -24995
rect 108496 -25095 117196 -25039
rect 108496 -25139 109104 -25095
rect 109148 -25139 109204 -25095
rect 109248 -25139 109304 -25095
rect 109348 -25139 109404 -25095
rect 109448 -25139 109504 -25095
rect 109548 -25139 109604 -25095
rect 109648 -25139 109704 -25095
rect 109748 -25139 109804 -25095
rect 109848 -25139 109904 -25095
rect 109948 -25139 110004 -25095
rect 110048 -25139 110104 -25095
rect 110148 -25139 110204 -25095
rect 110248 -25139 110304 -25095
rect 110348 -25139 110404 -25095
rect 110448 -25139 110504 -25095
rect 110548 -25139 110604 -25095
rect 110648 -25139 111104 -25095
rect 111148 -25139 111204 -25095
rect 111248 -25139 111304 -25095
rect 111348 -25139 111404 -25095
rect 111448 -25139 111504 -25095
rect 111548 -25139 111604 -25095
rect 111648 -25139 111704 -25095
rect 111748 -25139 111804 -25095
rect 111848 -25139 111904 -25095
rect 111948 -25139 112004 -25095
rect 112048 -25139 112104 -25095
rect 112148 -25139 112204 -25095
rect 112248 -25139 112304 -25095
rect 112348 -25139 112404 -25095
rect 112448 -25139 112504 -25095
rect 112548 -25139 112604 -25095
rect 112648 -25139 113104 -25095
rect 113148 -25139 113204 -25095
rect 113248 -25139 113304 -25095
rect 113348 -25139 113404 -25095
rect 113448 -25139 113504 -25095
rect 113548 -25139 113604 -25095
rect 113648 -25139 113704 -25095
rect 113748 -25139 113804 -25095
rect 113848 -25139 113904 -25095
rect 113948 -25139 114004 -25095
rect 114048 -25139 114104 -25095
rect 114148 -25139 114204 -25095
rect 114248 -25139 114304 -25095
rect 114348 -25139 114404 -25095
rect 114448 -25139 114504 -25095
rect 114548 -25139 114604 -25095
rect 114648 -25139 115104 -25095
rect 115148 -25139 115204 -25095
rect 115248 -25139 115304 -25095
rect 115348 -25139 115404 -25095
rect 115448 -25139 115504 -25095
rect 115548 -25139 115604 -25095
rect 115648 -25139 115704 -25095
rect 115748 -25139 115804 -25095
rect 115848 -25139 115904 -25095
rect 115948 -25139 116004 -25095
rect 116048 -25139 116104 -25095
rect 116148 -25139 116204 -25095
rect 116248 -25139 116304 -25095
rect 116348 -25139 116404 -25095
rect 116448 -25139 116504 -25095
rect 116548 -25139 116604 -25095
rect 116648 -25139 117196 -25095
rect 108496 -25195 117196 -25139
rect 108496 -25239 109104 -25195
rect 109148 -25239 109204 -25195
rect 109248 -25239 109304 -25195
rect 109348 -25239 109404 -25195
rect 109448 -25239 109504 -25195
rect 109548 -25239 109604 -25195
rect 109648 -25239 109704 -25195
rect 109748 -25239 109804 -25195
rect 109848 -25239 109904 -25195
rect 109948 -25239 110004 -25195
rect 110048 -25239 110104 -25195
rect 110148 -25239 110204 -25195
rect 110248 -25239 110304 -25195
rect 110348 -25239 110404 -25195
rect 110448 -25239 110504 -25195
rect 110548 -25239 110604 -25195
rect 110648 -25239 111104 -25195
rect 111148 -25239 111204 -25195
rect 111248 -25239 111304 -25195
rect 111348 -25239 111404 -25195
rect 111448 -25239 111504 -25195
rect 111548 -25239 111604 -25195
rect 111648 -25239 111704 -25195
rect 111748 -25239 111804 -25195
rect 111848 -25239 111904 -25195
rect 111948 -25239 112004 -25195
rect 112048 -25239 112104 -25195
rect 112148 -25239 112204 -25195
rect 112248 -25239 112304 -25195
rect 112348 -25239 112404 -25195
rect 112448 -25239 112504 -25195
rect 112548 -25239 112604 -25195
rect 112648 -25239 113104 -25195
rect 113148 -25239 113204 -25195
rect 113248 -25239 113304 -25195
rect 113348 -25239 113404 -25195
rect 113448 -25239 113504 -25195
rect 113548 -25239 113604 -25195
rect 113648 -25239 113704 -25195
rect 113748 -25239 113804 -25195
rect 113848 -25239 113904 -25195
rect 113948 -25239 114004 -25195
rect 114048 -25239 114104 -25195
rect 114148 -25239 114204 -25195
rect 114248 -25239 114304 -25195
rect 114348 -25239 114404 -25195
rect 114448 -25239 114504 -25195
rect 114548 -25239 114604 -25195
rect 114648 -25239 115104 -25195
rect 115148 -25239 115204 -25195
rect 115248 -25239 115304 -25195
rect 115348 -25239 115404 -25195
rect 115448 -25239 115504 -25195
rect 115548 -25239 115604 -25195
rect 115648 -25239 115704 -25195
rect 115748 -25239 115804 -25195
rect 115848 -25239 115904 -25195
rect 115948 -25239 116004 -25195
rect 116048 -25239 116104 -25195
rect 116148 -25239 116204 -25195
rect 116248 -25239 116304 -25195
rect 116348 -25239 116404 -25195
rect 116448 -25239 116504 -25195
rect 116548 -25239 116604 -25195
rect 116648 -25239 117196 -25195
rect 108496 -25295 117196 -25239
rect 108496 -25339 109104 -25295
rect 109148 -25339 109204 -25295
rect 109248 -25339 109304 -25295
rect 109348 -25339 109404 -25295
rect 109448 -25339 109504 -25295
rect 109548 -25339 109604 -25295
rect 109648 -25339 109704 -25295
rect 109748 -25339 109804 -25295
rect 109848 -25339 109904 -25295
rect 109948 -25339 110004 -25295
rect 110048 -25339 110104 -25295
rect 110148 -25339 110204 -25295
rect 110248 -25339 110304 -25295
rect 110348 -25339 110404 -25295
rect 110448 -25339 110504 -25295
rect 110548 -25339 110604 -25295
rect 110648 -25339 111104 -25295
rect 111148 -25339 111204 -25295
rect 111248 -25339 111304 -25295
rect 111348 -25339 111404 -25295
rect 111448 -25339 111504 -25295
rect 111548 -25339 111604 -25295
rect 111648 -25339 111704 -25295
rect 111748 -25339 111804 -25295
rect 111848 -25339 111904 -25295
rect 111948 -25339 112004 -25295
rect 112048 -25339 112104 -25295
rect 112148 -25339 112204 -25295
rect 112248 -25339 112304 -25295
rect 112348 -25339 112404 -25295
rect 112448 -25339 112504 -25295
rect 112548 -25339 112604 -25295
rect 112648 -25339 113104 -25295
rect 113148 -25339 113204 -25295
rect 113248 -25339 113304 -25295
rect 113348 -25339 113404 -25295
rect 113448 -25339 113504 -25295
rect 113548 -25339 113604 -25295
rect 113648 -25339 113704 -25295
rect 113748 -25339 113804 -25295
rect 113848 -25339 113904 -25295
rect 113948 -25339 114004 -25295
rect 114048 -25339 114104 -25295
rect 114148 -25339 114204 -25295
rect 114248 -25339 114304 -25295
rect 114348 -25339 114404 -25295
rect 114448 -25339 114504 -25295
rect 114548 -25339 114604 -25295
rect 114648 -25339 115104 -25295
rect 115148 -25339 115204 -25295
rect 115248 -25339 115304 -25295
rect 115348 -25339 115404 -25295
rect 115448 -25339 115504 -25295
rect 115548 -25339 115604 -25295
rect 115648 -25339 115704 -25295
rect 115748 -25339 115804 -25295
rect 115848 -25339 115904 -25295
rect 115948 -25339 116004 -25295
rect 116048 -25339 116104 -25295
rect 116148 -25339 116204 -25295
rect 116248 -25339 116304 -25295
rect 116348 -25339 116404 -25295
rect 116448 -25339 116504 -25295
rect 116548 -25339 116604 -25295
rect 116648 -25339 117196 -25295
rect 108496 -25395 117196 -25339
rect 108496 -25439 109104 -25395
rect 109148 -25439 109204 -25395
rect 109248 -25439 109304 -25395
rect 109348 -25439 109404 -25395
rect 109448 -25439 109504 -25395
rect 109548 -25439 109604 -25395
rect 109648 -25439 109704 -25395
rect 109748 -25439 109804 -25395
rect 109848 -25439 109904 -25395
rect 109948 -25439 110004 -25395
rect 110048 -25439 110104 -25395
rect 110148 -25439 110204 -25395
rect 110248 -25439 110304 -25395
rect 110348 -25439 110404 -25395
rect 110448 -25439 110504 -25395
rect 110548 -25439 110604 -25395
rect 110648 -25439 111104 -25395
rect 111148 -25439 111204 -25395
rect 111248 -25439 111304 -25395
rect 111348 -25439 111404 -25395
rect 111448 -25439 111504 -25395
rect 111548 -25439 111604 -25395
rect 111648 -25439 111704 -25395
rect 111748 -25439 111804 -25395
rect 111848 -25439 111904 -25395
rect 111948 -25439 112004 -25395
rect 112048 -25439 112104 -25395
rect 112148 -25439 112204 -25395
rect 112248 -25439 112304 -25395
rect 112348 -25439 112404 -25395
rect 112448 -25439 112504 -25395
rect 112548 -25439 112604 -25395
rect 112648 -25439 113104 -25395
rect 113148 -25439 113204 -25395
rect 113248 -25439 113304 -25395
rect 113348 -25439 113404 -25395
rect 113448 -25439 113504 -25395
rect 113548 -25439 113604 -25395
rect 113648 -25439 113704 -25395
rect 113748 -25439 113804 -25395
rect 113848 -25439 113904 -25395
rect 113948 -25439 114004 -25395
rect 114048 -25439 114104 -25395
rect 114148 -25439 114204 -25395
rect 114248 -25439 114304 -25395
rect 114348 -25439 114404 -25395
rect 114448 -25439 114504 -25395
rect 114548 -25439 114604 -25395
rect 114648 -25439 115104 -25395
rect 115148 -25439 115204 -25395
rect 115248 -25439 115304 -25395
rect 115348 -25439 115404 -25395
rect 115448 -25439 115504 -25395
rect 115548 -25439 115604 -25395
rect 115648 -25439 115704 -25395
rect 115748 -25439 115804 -25395
rect 115848 -25439 115904 -25395
rect 115948 -25439 116004 -25395
rect 116048 -25439 116104 -25395
rect 116148 -25439 116204 -25395
rect 116248 -25439 116304 -25395
rect 116348 -25439 116404 -25395
rect 116448 -25439 116504 -25395
rect 116548 -25439 116604 -25395
rect 116648 -25439 117196 -25395
rect 108496 -25495 117196 -25439
rect 108496 -25539 109104 -25495
rect 109148 -25539 109204 -25495
rect 109248 -25539 109304 -25495
rect 109348 -25539 109404 -25495
rect 109448 -25539 109504 -25495
rect 109548 -25539 109604 -25495
rect 109648 -25539 109704 -25495
rect 109748 -25539 109804 -25495
rect 109848 -25539 109904 -25495
rect 109948 -25539 110004 -25495
rect 110048 -25539 110104 -25495
rect 110148 -25539 110204 -25495
rect 110248 -25539 110304 -25495
rect 110348 -25539 110404 -25495
rect 110448 -25539 110504 -25495
rect 110548 -25539 110604 -25495
rect 110648 -25539 111104 -25495
rect 111148 -25539 111204 -25495
rect 111248 -25539 111304 -25495
rect 111348 -25539 111404 -25495
rect 111448 -25539 111504 -25495
rect 111548 -25539 111604 -25495
rect 111648 -25539 111704 -25495
rect 111748 -25539 111804 -25495
rect 111848 -25539 111904 -25495
rect 111948 -25539 112004 -25495
rect 112048 -25539 112104 -25495
rect 112148 -25539 112204 -25495
rect 112248 -25539 112304 -25495
rect 112348 -25539 112404 -25495
rect 112448 -25539 112504 -25495
rect 112548 -25539 112604 -25495
rect 112648 -25539 113104 -25495
rect 113148 -25539 113204 -25495
rect 113248 -25539 113304 -25495
rect 113348 -25539 113404 -25495
rect 113448 -25539 113504 -25495
rect 113548 -25539 113604 -25495
rect 113648 -25539 113704 -25495
rect 113748 -25539 113804 -25495
rect 113848 -25539 113904 -25495
rect 113948 -25539 114004 -25495
rect 114048 -25539 114104 -25495
rect 114148 -25539 114204 -25495
rect 114248 -25539 114304 -25495
rect 114348 -25539 114404 -25495
rect 114448 -25539 114504 -25495
rect 114548 -25539 114604 -25495
rect 114648 -25539 115104 -25495
rect 115148 -25539 115204 -25495
rect 115248 -25539 115304 -25495
rect 115348 -25539 115404 -25495
rect 115448 -25539 115504 -25495
rect 115548 -25539 115604 -25495
rect 115648 -25539 115704 -25495
rect 115748 -25539 115804 -25495
rect 115848 -25539 115904 -25495
rect 115948 -25539 116004 -25495
rect 116048 -25539 116104 -25495
rect 116148 -25539 116204 -25495
rect 116248 -25539 116304 -25495
rect 116348 -25539 116404 -25495
rect 116448 -25539 116504 -25495
rect 116548 -25539 116604 -25495
rect 116648 -25539 117196 -25495
rect 108496 -25595 117196 -25539
rect 108496 -25639 109104 -25595
rect 109148 -25639 109204 -25595
rect 109248 -25639 109304 -25595
rect 109348 -25639 109404 -25595
rect 109448 -25639 109504 -25595
rect 109548 -25639 109604 -25595
rect 109648 -25639 109704 -25595
rect 109748 -25639 109804 -25595
rect 109848 -25639 109904 -25595
rect 109948 -25639 110004 -25595
rect 110048 -25639 110104 -25595
rect 110148 -25639 110204 -25595
rect 110248 -25639 110304 -25595
rect 110348 -25639 110404 -25595
rect 110448 -25639 110504 -25595
rect 110548 -25639 110604 -25595
rect 110648 -25639 111104 -25595
rect 111148 -25639 111204 -25595
rect 111248 -25639 111304 -25595
rect 111348 -25639 111404 -25595
rect 111448 -25639 111504 -25595
rect 111548 -25639 111604 -25595
rect 111648 -25639 111704 -25595
rect 111748 -25639 111804 -25595
rect 111848 -25639 111904 -25595
rect 111948 -25639 112004 -25595
rect 112048 -25639 112104 -25595
rect 112148 -25639 112204 -25595
rect 112248 -25639 112304 -25595
rect 112348 -25639 112404 -25595
rect 112448 -25639 112504 -25595
rect 112548 -25639 112604 -25595
rect 112648 -25639 113104 -25595
rect 113148 -25639 113204 -25595
rect 113248 -25639 113304 -25595
rect 113348 -25639 113404 -25595
rect 113448 -25639 113504 -25595
rect 113548 -25639 113604 -25595
rect 113648 -25639 113704 -25595
rect 113748 -25639 113804 -25595
rect 113848 -25639 113904 -25595
rect 113948 -25639 114004 -25595
rect 114048 -25639 114104 -25595
rect 114148 -25639 114204 -25595
rect 114248 -25639 114304 -25595
rect 114348 -25639 114404 -25595
rect 114448 -25639 114504 -25595
rect 114548 -25639 114604 -25595
rect 114648 -25639 115104 -25595
rect 115148 -25639 115204 -25595
rect 115248 -25639 115304 -25595
rect 115348 -25639 115404 -25595
rect 115448 -25639 115504 -25595
rect 115548 -25639 115604 -25595
rect 115648 -25639 115704 -25595
rect 115748 -25639 115804 -25595
rect 115848 -25639 115904 -25595
rect 115948 -25639 116004 -25595
rect 116048 -25639 116104 -25595
rect 116148 -25639 116204 -25595
rect 116248 -25639 116304 -25595
rect 116348 -25639 116404 -25595
rect 116448 -25639 116504 -25595
rect 116548 -25639 116604 -25595
rect 116648 -25639 117196 -25595
rect 108496 -25695 117196 -25639
rect 108496 -25739 109104 -25695
rect 109148 -25739 109204 -25695
rect 109248 -25739 109304 -25695
rect 109348 -25739 109404 -25695
rect 109448 -25739 109504 -25695
rect 109548 -25739 109604 -25695
rect 109648 -25739 109704 -25695
rect 109748 -25739 109804 -25695
rect 109848 -25739 109904 -25695
rect 109948 -25739 110004 -25695
rect 110048 -25739 110104 -25695
rect 110148 -25739 110204 -25695
rect 110248 -25739 110304 -25695
rect 110348 -25739 110404 -25695
rect 110448 -25739 110504 -25695
rect 110548 -25739 110604 -25695
rect 110648 -25739 111104 -25695
rect 111148 -25739 111204 -25695
rect 111248 -25739 111304 -25695
rect 111348 -25739 111404 -25695
rect 111448 -25739 111504 -25695
rect 111548 -25739 111604 -25695
rect 111648 -25739 111704 -25695
rect 111748 -25739 111804 -25695
rect 111848 -25739 111904 -25695
rect 111948 -25739 112004 -25695
rect 112048 -25739 112104 -25695
rect 112148 -25739 112204 -25695
rect 112248 -25739 112304 -25695
rect 112348 -25739 112404 -25695
rect 112448 -25739 112504 -25695
rect 112548 -25739 112604 -25695
rect 112648 -25739 113104 -25695
rect 113148 -25739 113204 -25695
rect 113248 -25739 113304 -25695
rect 113348 -25739 113404 -25695
rect 113448 -25739 113504 -25695
rect 113548 -25739 113604 -25695
rect 113648 -25739 113704 -25695
rect 113748 -25739 113804 -25695
rect 113848 -25739 113904 -25695
rect 113948 -25739 114004 -25695
rect 114048 -25739 114104 -25695
rect 114148 -25739 114204 -25695
rect 114248 -25739 114304 -25695
rect 114348 -25739 114404 -25695
rect 114448 -25739 114504 -25695
rect 114548 -25739 114604 -25695
rect 114648 -25739 115104 -25695
rect 115148 -25739 115204 -25695
rect 115248 -25739 115304 -25695
rect 115348 -25739 115404 -25695
rect 115448 -25739 115504 -25695
rect 115548 -25739 115604 -25695
rect 115648 -25739 115704 -25695
rect 115748 -25739 115804 -25695
rect 115848 -25739 115904 -25695
rect 115948 -25739 116004 -25695
rect 116048 -25739 116104 -25695
rect 116148 -25739 116204 -25695
rect 116248 -25739 116304 -25695
rect 116348 -25739 116404 -25695
rect 116448 -25739 116504 -25695
rect 116548 -25739 116604 -25695
rect 116648 -25739 117196 -25695
rect 108496 -51137 117196 -25739
rect 108496 -51181 109305 -51137
rect 109349 -51181 109405 -51137
rect 109449 -51181 109505 -51137
rect 109549 -51181 109605 -51137
rect 109649 -51181 109705 -51137
rect 109749 -51181 109805 -51137
rect 109849 -51181 109905 -51137
rect 109949 -51181 110005 -51137
rect 110049 -51181 110105 -51137
rect 110149 -51181 110205 -51137
rect 110249 -51181 110305 -51137
rect 110349 -51181 110405 -51137
rect 110449 -51181 110505 -51137
rect 110549 -51181 110605 -51137
rect 110649 -51181 110705 -51137
rect 110749 -51181 110805 -51137
rect 110849 -51181 111305 -51137
rect 111349 -51181 111405 -51137
rect 111449 -51181 111505 -51137
rect 111549 -51181 111605 -51137
rect 111649 -51181 111705 -51137
rect 111749 -51181 111805 -51137
rect 111849 -51181 111905 -51137
rect 111949 -51181 112005 -51137
rect 112049 -51181 112105 -51137
rect 112149 -51181 112205 -51137
rect 112249 -51181 112305 -51137
rect 112349 -51181 112405 -51137
rect 112449 -51181 112505 -51137
rect 112549 -51181 112605 -51137
rect 112649 -51181 112705 -51137
rect 112749 -51181 112805 -51137
rect 112849 -51181 113305 -51137
rect 113349 -51181 113405 -51137
rect 113449 -51181 113505 -51137
rect 113549 -51181 113605 -51137
rect 113649 -51181 113705 -51137
rect 113749 -51181 113805 -51137
rect 113849 -51181 113905 -51137
rect 113949 -51181 114005 -51137
rect 114049 -51181 114105 -51137
rect 114149 -51181 114205 -51137
rect 114249 -51181 114305 -51137
rect 114349 -51181 114405 -51137
rect 114449 -51181 114505 -51137
rect 114549 -51181 114605 -51137
rect 114649 -51181 114705 -51137
rect 114749 -51181 114805 -51137
rect 114849 -51181 115305 -51137
rect 115349 -51181 115405 -51137
rect 115449 -51181 115505 -51137
rect 115549 -51181 115605 -51137
rect 115649 -51181 115705 -51137
rect 115749 -51181 115805 -51137
rect 115849 -51181 115905 -51137
rect 115949 -51181 116005 -51137
rect 116049 -51181 116105 -51137
rect 116149 -51181 116205 -51137
rect 116249 -51181 116305 -51137
rect 116349 -51181 116405 -51137
rect 116449 -51181 116505 -51137
rect 116549 -51181 116605 -51137
rect 116649 -51181 116705 -51137
rect 116749 -51181 116805 -51137
rect 116849 -51181 117196 -51137
rect 108496 -51237 117196 -51181
rect 108496 -51281 109305 -51237
rect 109349 -51281 109405 -51237
rect 109449 -51281 109505 -51237
rect 109549 -51281 109605 -51237
rect 109649 -51281 109705 -51237
rect 109749 -51281 109805 -51237
rect 109849 -51281 109905 -51237
rect 109949 -51281 110005 -51237
rect 110049 -51281 110105 -51237
rect 110149 -51281 110205 -51237
rect 110249 -51281 110305 -51237
rect 110349 -51281 110405 -51237
rect 110449 -51281 110505 -51237
rect 110549 -51281 110605 -51237
rect 110649 -51281 110705 -51237
rect 110749 -51281 110805 -51237
rect 110849 -51281 111305 -51237
rect 111349 -51281 111405 -51237
rect 111449 -51281 111505 -51237
rect 111549 -51281 111605 -51237
rect 111649 -51281 111705 -51237
rect 111749 -51281 111805 -51237
rect 111849 -51281 111905 -51237
rect 111949 -51281 112005 -51237
rect 112049 -51281 112105 -51237
rect 112149 -51281 112205 -51237
rect 112249 -51281 112305 -51237
rect 112349 -51281 112405 -51237
rect 112449 -51281 112505 -51237
rect 112549 -51281 112605 -51237
rect 112649 -51281 112705 -51237
rect 112749 -51281 112805 -51237
rect 112849 -51281 113305 -51237
rect 113349 -51281 113405 -51237
rect 113449 -51281 113505 -51237
rect 113549 -51281 113605 -51237
rect 113649 -51281 113705 -51237
rect 113749 -51281 113805 -51237
rect 113849 -51281 113905 -51237
rect 113949 -51281 114005 -51237
rect 114049 -51281 114105 -51237
rect 114149 -51281 114205 -51237
rect 114249 -51281 114305 -51237
rect 114349 -51281 114405 -51237
rect 114449 -51281 114505 -51237
rect 114549 -51281 114605 -51237
rect 114649 -51281 114705 -51237
rect 114749 -51281 114805 -51237
rect 114849 -51281 115305 -51237
rect 115349 -51281 115405 -51237
rect 115449 -51281 115505 -51237
rect 115549 -51281 115605 -51237
rect 115649 -51281 115705 -51237
rect 115749 -51281 115805 -51237
rect 115849 -51281 115905 -51237
rect 115949 -51281 116005 -51237
rect 116049 -51281 116105 -51237
rect 116149 -51281 116205 -51237
rect 116249 -51281 116305 -51237
rect 116349 -51281 116405 -51237
rect 116449 -51281 116505 -51237
rect 116549 -51281 116605 -51237
rect 116649 -51281 116705 -51237
rect 116749 -51281 116805 -51237
rect 116849 -51281 117196 -51237
rect 108496 -51337 117196 -51281
rect 108496 -51381 109305 -51337
rect 109349 -51381 109405 -51337
rect 109449 -51381 109505 -51337
rect 109549 -51381 109605 -51337
rect 109649 -51381 109705 -51337
rect 109749 -51381 109805 -51337
rect 109849 -51381 109905 -51337
rect 109949 -51381 110005 -51337
rect 110049 -51381 110105 -51337
rect 110149 -51381 110205 -51337
rect 110249 -51381 110305 -51337
rect 110349 -51381 110405 -51337
rect 110449 -51381 110505 -51337
rect 110549 -51381 110605 -51337
rect 110649 -51381 110705 -51337
rect 110749 -51381 110805 -51337
rect 110849 -51381 111305 -51337
rect 111349 -51381 111405 -51337
rect 111449 -51381 111505 -51337
rect 111549 -51381 111605 -51337
rect 111649 -51381 111705 -51337
rect 111749 -51381 111805 -51337
rect 111849 -51381 111905 -51337
rect 111949 -51381 112005 -51337
rect 112049 -51381 112105 -51337
rect 112149 -51381 112205 -51337
rect 112249 -51381 112305 -51337
rect 112349 -51381 112405 -51337
rect 112449 -51381 112505 -51337
rect 112549 -51381 112605 -51337
rect 112649 -51381 112705 -51337
rect 112749 -51381 112805 -51337
rect 112849 -51381 113305 -51337
rect 113349 -51381 113405 -51337
rect 113449 -51381 113505 -51337
rect 113549 -51381 113605 -51337
rect 113649 -51381 113705 -51337
rect 113749 -51381 113805 -51337
rect 113849 -51381 113905 -51337
rect 113949 -51381 114005 -51337
rect 114049 -51381 114105 -51337
rect 114149 -51381 114205 -51337
rect 114249 -51381 114305 -51337
rect 114349 -51381 114405 -51337
rect 114449 -51381 114505 -51337
rect 114549 -51381 114605 -51337
rect 114649 -51381 114705 -51337
rect 114749 -51381 114805 -51337
rect 114849 -51381 115305 -51337
rect 115349 -51381 115405 -51337
rect 115449 -51381 115505 -51337
rect 115549 -51381 115605 -51337
rect 115649 -51381 115705 -51337
rect 115749 -51381 115805 -51337
rect 115849 -51381 115905 -51337
rect 115949 -51381 116005 -51337
rect 116049 -51381 116105 -51337
rect 116149 -51381 116205 -51337
rect 116249 -51381 116305 -51337
rect 116349 -51381 116405 -51337
rect 116449 -51381 116505 -51337
rect 116549 -51381 116605 -51337
rect 116649 -51381 116705 -51337
rect 116749 -51381 116805 -51337
rect 116849 -51381 117196 -51337
rect 108496 -51437 117196 -51381
rect 108496 -51481 109305 -51437
rect 109349 -51481 109405 -51437
rect 109449 -51481 109505 -51437
rect 109549 -51481 109605 -51437
rect 109649 -51481 109705 -51437
rect 109749 -51481 109805 -51437
rect 109849 -51481 109905 -51437
rect 109949 -51481 110005 -51437
rect 110049 -51481 110105 -51437
rect 110149 -51481 110205 -51437
rect 110249 -51481 110305 -51437
rect 110349 -51481 110405 -51437
rect 110449 -51481 110505 -51437
rect 110549 -51481 110605 -51437
rect 110649 -51481 110705 -51437
rect 110749 -51481 110805 -51437
rect 110849 -51481 111305 -51437
rect 111349 -51481 111405 -51437
rect 111449 -51481 111505 -51437
rect 111549 -51481 111605 -51437
rect 111649 -51481 111705 -51437
rect 111749 -51481 111805 -51437
rect 111849 -51481 111905 -51437
rect 111949 -51481 112005 -51437
rect 112049 -51481 112105 -51437
rect 112149 -51481 112205 -51437
rect 112249 -51481 112305 -51437
rect 112349 -51481 112405 -51437
rect 112449 -51481 112505 -51437
rect 112549 -51481 112605 -51437
rect 112649 -51481 112705 -51437
rect 112749 -51481 112805 -51437
rect 112849 -51481 113305 -51437
rect 113349 -51481 113405 -51437
rect 113449 -51481 113505 -51437
rect 113549 -51481 113605 -51437
rect 113649 -51481 113705 -51437
rect 113749 -51481 113805 -51437
rect 113849 -51481 113905 -51437
rect 113949 -51481 114005 -51437
rect 114049 -51481 114105 -51437
rect 114149 -51481 114205 -51437
rect 114249 -51481 114305 -51437
rect 114349 -51481 114405 -51437
rect 114449 -51481 114505 -51437
rect 114549 -51481 114605 -51437
rect 114649 -51481 114705 -51437
rect 114749 -51481 114805 -51437
rect 114849 -51481 115305 -51437
rect 115349 -51481 115405 -51437
rect 115449 -51481 115505 -51437
rect 115549 -51481 115605 -51437
rect 115649 -51481 115705 -51437
rect 115749 -51481 115805 -51437
rect 115849 -51481 115905 -51437
rect 115949 -51481 116005 -51437
rect 116049 -51481 116105 -51437
rect 116149 -51481 116205 -51437
rect 116249 -51481 116305 -51437
rect 116349 -51481 116405 -51437
rect 116449 -51481 116505 -51437
rect 116549 -51481 116605 -51437
rect 116649 -51481 116705 -51437
rect 116749 -51481 116805 -51437
rect 116849 -51481 117196 -51437
rect 108496 -51537 117196 -51481
rect 108496 -51581 109305 -51537
rect 109349 -51581 109405 -51537
rect 109449 -51581 109505 -51537
rect 109549 -51581 109605 -51537
rect 109649 -51581 109705 -51537
rect 109749 -51581 109805 -51537
rect 109849 -51581 109905 -51537
rect 109949 -51581 110005 -51537
rect 110049 -51581 110105 -51537
rect 110149 -51581 110205 -51537
rect 110249 -51581 110305 -51537
rect 110349 -51581 110405 -51537
rect 110449 -51581 110505 -51537
rect 110549 -51581 110605 -51537
rect 110649 -51581 110705 -51537
rect 110749 -51581 110805 -51537
rect 110849 -51581 111305 -51537
rect 111349 -51581 111405 -51537
rect 111449 -51581 111505 -51537
rect 111549 -51581 111605 -51537
rect 111649 -51581 111705 -51537
rect 111749 -51581 111805 -51537
rect 111849 -51581 111905 -51537
rect 111949 -51581 112005 -51537
rect 112049 -51581 112105 -51537
rect 112149 -51581 112205 -51537
rect 112249 -51581 112305 -51537
rect 112349 -51581 112405 -51537
rect 112449 -51581 112505 -51537
rect 112549 -51581 112605 -51537
rect 112649 -51581 112705 -51537
rect 112749 -51581 112805 -51537
rect 112849 -51581 113305 -51537
rect 113349 -51581 113405 -51537
rect 113449 -51581 113505 -51537
rect 113549 -51581 113605 -51537
rect 113649 -51581 113705 -51537
rect 113749 -51581 113805 -51537
rect 113849 -51581 113905 -51537
rect 113949 -51581 114005 -51537
rect 114049 -51581 114105 -51537
rect 114149 -51581 114205 -51537
rect 114249 -51581 114305 -51537
rect 114349 -51581 114405 -51537
rect 114449 -51581 114505 -51537
rect 114549 -51581 114605 -51537
rect 114649 -51581 114705 -51537
rect 114749 -51581 114805 -51537
rect 114849 -51581 115305 -51537
rect 115349 -51581 115405 -51537
rect 115449 -51581 115505 -51537
rect 115549 -51581 115605 -51537
rect 115649 -51581 115705 -51537
rect 115749 -51581 115805 -51537
rect 115849 -51581 115905 -51537
rect 115949 -51581 116005 -51537
rect 116049 -51581 116105 -51537
rect 116149 -51581 116205 -51537
rect 116249 -51581 116305 -51537
rect 116349 -51581 116405 -51537
rect 116449 -51581 116505 -51537
rect 116549 -51581 116605 -51537
rect 116649 -51581 116705 -51537
rect 116749 -51581 116805 -51537
rect 116849 -51581 117196 -51537
rect 108496 -51637 117196 -51581
rect 108496 -51681 109305 -51637
rect 109349 -51681 109405 -51637
rect 109449 -51681 109505 -51637
rect 109549 -51681 109605 -51637
rect 109649 -51681 109705 -51637
rect 109749 -51681 109805 -51637
rect 109849 -51681 109905 -51637
rect 109949 -51681 110005 -51637
rect 110049 -51681 110105 -51637
rect 110149 -51681 110205 -51637
rect 110249 -51681 110305 -51637
rect 110349 -51681 110405 -51637
rect 110449 -51681 110505 -51637
rect 110549 -51681 110605 -51637
rect 110649 -51681 110705 -51637
rect 110749 -51681 110805 -51637
rect 110849 -51681 111305 -51637
rect 111349 -51681 111405 -51637
rect 111449 -51681 111505 -51637
rect 111549 -51681 111605 -51637
rect 111649 -51681 111705 -51637
rect 111749 -51681 111805 -51637
rect 111849 -51681 111905 -51637
rect 111949 -51681 112005 -51637
rect 112049 -51681 112105 -51637
rect 112149 -51681 112205 -51637
rect 112249 -51681 112305 -51637
rect 112349 -51681 112405 -51637
rect 112449 -51681 112505 -51637
rect 112549 -51681 112605 -51637
rect 112649 -51681 112705 -51637
rect 112749 -51681 112805 -51637
rect 112849 -51681 113305 -51637
rect 113349 -51681 113405 -51637
rect 113449 -51681 113505 -51637
rect 113549 -51681 113605 -51637
rect 113649 -51681 113705 -51637
rect 113749 -51681 113805 -51637
rect 113849 -51681 113905 -51637
rect 113949 -51681 114005 -51637
rect 114049 -51681 114105 -51637
rect 114149 -51681 114205 -51637
rect 114249 -51681 114305 -51637
rect 114349 -51681 114405 -51637
rect 114449 -51681 114505 -51637
rect 114549 -51681 114605 -51637
rect 114649 -51681 114705 -51637
rect 114749 -51681 114805 -51637
rect 114849 -51681 115305 -51637
rect 115349 -51681 115405 -51637
rect 115449 -51681 115505 -51637
rect 115549 -51681 115605 -51637
rect 115649 -51681 115705 -51637
rect 115749 -51681 115805 -51637
rect 115849 -51681 115905 -51637
rect 115949 -51681 116005 -51637
rect 116049 -51681 116105 -51637
rect 116149 -51681 116205 -51637
rect 116249 -51681 116305 -51637
rect 116349 -51681 116405 -51637
rect 116449 -51681 116505 -51637
rect 116549 -51681 116605 -51637
rect 116649 -51681 116705 -51637
rect 116749 -51681 116805 -51637
rect 116849 -51681 117196 -51637
rect 108496 -51737 117196 -51681
rect 108496 -51781 109305 -51737
rect 109349 -51781 109405 -51737
rect 109449 -51781 109505 -51737
rect 109549 -51781 109605 -51737
rect 109649 -51781 109705 -51737
rect 109749 -51781 109805 -51737
rect 109849 -51781 109905 -51737
rect 109949 -51781 110005 -51737
rect 110049 -51781 110105 -51737
rect 110149 -51781 110205 -51737
rect 110249 -51781 110305 -51737
rect 110349 -51781 110405 -51737
rect 110449 -51781 110505 -51737
rect 110549 -51781 110605 -51737
rect 110649 -51781 110705 -51737
rect 110749 -51781 110805 -51737
rect 110849 -51781 111305 -51737
rect 111349 -51781 111405 -51737
rect 111449 -51781 111505 -51737
rect 111549 -51781 111605 -51737
rect 111649 -51781 111705 -51737
rect 111749 -51781 111805 -51737
rect 111849 -51781 111905 -51737
rect 111949 -51781 112005 -51737
rect 112049 -51781 112105 -51737
rect 112149 -51781 112205 -51737
rect 112249 -51781 112305 -51737
rect 112349 -51781 112405 -51737
rect 112449 -51781 112505 -51737
rect 112549 -51781 112605 -51737
rect 112649 -51781 112705 -51737
rect 112749 -51781 112805 -51737
rect 112849 -51781 113305 -51737
rect 113349 -51781 113405 -51737
rect 113449 -51781 113505 -51737
rect 113549 -51781 113605 -51737
rect 113649 -51781 113705 -51737
rect 113749 -51781 113805 -51737
rect 113849 -51781 113905 -51737
rect 113949 -51781 114005 -51737
rect 114049 -51781 114105 -51737
rect 114149 -51781 114205 -51737
rect 114249 -51781 114305 -51737
rect 114349 -51781 114405 -51737
rect 114449 -51781 114505 -51737
rect 114549 -51781 114605 -51737
rect 114649 -51781 114705 -51737
rect 114749 -51781 114805 -51737
rect 114849 -51781 115305 -51737
rect 115349 -51781 115405 -51737
rect 115449 -51781 115505 -51737
rect 115549 -51781 115605 -51737
rect 115649 -51781 115705 -51737
rect 115749 -51781 115805 -51737
rect 115849 -51781 115905 -51737
rect 115949 -51781 116005 -51737
rect 116049 -51781 116105 -51737
rect 116149 -51781 116205 -51737
rect 116249 -51781 116305 -51737
rect 116349 -51781 116405 -51737
rect 116449 -51781 116505 -51737
rect 116549 -51781 116605 -51737
rect 116649 -51781 116705 -51737
rect 116749 -51781 116805 -51737
rect 116849 -51781 117196 -51737
rect 108496 -51837 117196 -51781
rect 108496 -51881 109305 -51837
rect 109349 -51881 109405 -51837
rect 109449 -51881 109505 -51837
rect 109549 -51881 109605 -51837
rect 109649 -51881 109705 -51837
rect 109749 -51881 109805 -51837
rect 109849 -51881 109905 -51837
rect 109949 -51881 110005 -51837
rect 110049 -51881 110105 -51837
rect 110149 -51881 110205 -51837
rect 110249 -51881 110305 -51837
rect 110349 -51881 110405 -51837
rect 110449 -51881 110505 -51837
rect 110549 -51881 110605 -51837
rect 110649 -51881 110705 -51837
rect 110749 -51881 110805 -51837
rect 110849 -51881 111305 -51837
rect 111349 -51881 111405 -51837
rect 111449 -51881 111505 -51837
rect 111549 -51881 111605 -51837
rect 111649 -51881 111705 -51837
rect 111749 -51881 111805 -51837
rect 111849 -51881 111905 -51837
rect 111949 -51881 112005 -51837
rect 112049 -51881 112105 -51837
rect 112149 -51881 112205 -51837
rect 112249 -51881 112305 -51837
rect 112349 -51881 112405 -51837
rect 112449 -51881 112505 -51837
rect 112549 -51881 112605 -51837
rect 112649 -51881 112705 -51837
rect 112749 -51881 112805 -51837
rect 112849 -51881 113305 -51837
rect 113349 -51881 113405 -51837
rect 113449 -51881 113505 -51837
rect 113549 -51881 113605 -51837
rect 113649 -51881 113705 -51837
rect 113749 -51881 113805 -51837
rect 113849 -51881 113905 -51837
rect 113949 -51881 114005 -51837
rect 114049 -51881 114105 -51837
rect 114149 -51881 114205 -51837
rect 114249 -51881 114305 -51837
rect 114349 -51881 114405 -51837
rect 114449 -51881 114505 -51837
rect 114549 -51881 114605 -51837
rect 114649 -51881 114705 -51837
rect 114749 -51881 114805 -51837
rect 114849 -51881 115305 -51837
rect 115349 -51881 115405 -51837
rect 115449 -51881 115505 -51837
rect 115549 -51881 115605 -51837
rect 115649 -51881 115705 -51837
rect 115749 -51881 115805 -51837
rect 115849 -51881 115905 -51837
rect 115949 -51881 116005 -51837
rect 116049 -51881 116105 -51837
rect 116149 -51881 116205 -51837
rect 116249 -51881 116305 -51837
rect 116349 -51881 116405 -51837
rect 116449 -51881 116505 -51837
rect 116549 -51881 116605 -51837
rect 116649 -51881 116705 -51837
rect 116749 -51881 116805 -51837
rect 116849 -51881 117196 -51837
rect 108496 -51937 117196 -51881
rect 108496 -51981 109305 -51937
rect 109349 -51981 109405 -51937
rect 109449 -51981 109505 -51937
rect 109549 -51981 109605 -51937
rect 109649 -51981 109705 -51937
rect 109749 -51981 109805 -51937
rect 109849 -51981 109905 -51937
rect 109949 -51981 110005 -51937
rect 110049 -51981 110105 -51937
rect 110149 -51981 110205 -51937
rect 110249 -51981 110305 -51937
rect 110349 -51981 110405 -51937
rect 110449 -51981 110505 -51937
rect 110549 -51981 110605 -51937
rect 110649 -51981 110705 -51937
rect 110749 -51981 110805 -51937
rect 110849 -51981 111305 -51937
rect 111349 -51981 111405 -51937
rect 111449 -51981 111505 -51937
rect 111549 -51981 111605 -51937
rect 111649 -51981 111705 -51937
rect 111749 -51981 111805 -51937
rect 111849 -51981 111905 -51937
rect 111949 -51981 112005 -51937
rect 112049 -51981 112105 -51937
rect 112149 -51981 112205 -51937
rect 112249 -51981 112305 -51937
rect 112349 -51981 112405 -51937
rect 112449 -51981 112505 -51937
rect 112549 -51981 112605 -51937
rect 112649 -51981 112705 -51937
rect 112749 -51981 112805 -51937
rect 112849 -51981 113305 -51937
rect 113349 -51981 113405 -51937
rect 113449 -51981 113505 -51937
rect 113549 -51981 113605 -51937
rect 113649 -51981 113705 -51937
rect 113749 -51981 113805 -51937
rect 113849 -51981 113905 -51937
rect 113949 -51981 114005 -51937
rect 114049 -51981 114105 -51937
rect 114149 -51981 114205 -51937
rect 114249 -51981 114305 -51937
rect 114349 -51981 114405 -51937
rect 114449 -51981 114505 -51937
rect 114549 -51981 114605 -51937
rect 114649 -51981 114705 -51937
rect 114749 -51981 114805 -51937
rect 114849 -51981 115305 -51937
rect 115349 -51981 115405 -51937
rect 115449 -51981 115505 -51937
rect 115549 -51981 115605 -51937
rect 115649 -51981 115705 -51937
rect 115749 -51981 115805 -51937
rect 115849 -51981 115905 -51937
rect 115949 -51981 116005 -51937
rect 116049 -51981 116105 -51937
rect 116149 -51981 116205 -51937
rect 116249 -51981 116305 -51937
rect 116349 -51981 116405 -51937
rect 116449 -51981 116505 -51937
rect 116549 -51981 116605 -51937
rect 116649 -51981 116705 -51937
rect 116749 -51981 116805 -51937
rect 116849 -51981 117196 -51937
rect 108496 -52037 117196 -51981
rect 108496 -52081 109305 -52037
rect 109349 -52081 109405 -52037
rect 109449 -52081 109505 -52037
rect 109549 -52081 109605 -52037
rect 109649 -52081 109705 -52037
rect 109749 -52081 109805 -52037
rect 109849 -52081 109905 -52037
rect 109949 -52081 110005 -52037
rect 110049 -52081 110105 -52037
rect 110149 -52081 110205 -52037
rect 110249 -52081 110305 -52037
rect 110349 -52081 110405 -52037
rect 110449 -52081 110505 -52037
rect 110549 -52081 110605 -52037
rect 110649 -52081 110705 -52037
rect 110749 -52081 110805 -52037
rect 110849 -52081 111305 -52037
rect 111349 -52081 111405 -52037
rect 111449 -52081 111505 -52037
rect 111549 -52081 111605 -52037
rect 111649 -52081 111705 -52037
rect 111749 -52081 111805 -52037
rect 111849 -52081 111905 -52037
rect 111949 -52081 112005 -52037
rect 112049 -52081 112105 -52037
rect 112149 -52081 112205 -52037
rect 112249 -52081 112305 -52037
rect 112349 -52081 112405 -52037
rect 112449 -52081 112505 -52037
rect 112549 -52081 112605 -52037
rect 112649 -52081 112705 -52037
rect 112749 -52081 112805 -52037
rect 112849 -52081 113305 -52037
rect 113349 -52081 113405 -52037
rect 113449 -52081 113505 -52037
rect 113549 -52081 113605 -52037
rect 113649 -52081 113705 -52037
rect 113749 -52081 113805 -52037
rect 113849 -52081 113905 -52037
rect 113949 -52081 114005 -52037
rect 114049 -52081 114105 -52037
rect 114149 -52081 114205 -52037
rect 114249 -52081 114305 -52037
rect 114349 -52081 114405 -52037
rect 114449 -52081 114505 -52037
rect 114549 -52081 114605 -52037
rect 114649 -52081 114705 -52037
rect 114749 -52081 114805 -52037
rect 114849 -52081 115305 -52037
rect 115349 -52081 115405 -52037
rect 115449 -52081 115505 -52037
rect 115549 -52081 115605 -52037
rect 115649 -52081 115705 -52037
rect 115749 -52081 115805 -52037
rect 115849 -52081 115905 -52037
rect 115949 -52081 116005 -52037
rect 116049 -52081 116105 -52037
rect 116149 -52081 116205 -52037
rect 116249 -52081 116305 -52037
rect 116349 -52081 116405 -52037
rect 116449 -52081 116505 -52037
rect 116549 -52081 116605 -52037
rect 116649 -52081 116705 -52037
rect 116749 -52081 116805 -52037
rect 116849 -52081 117196 -52037
rect 108496 -52137 117196 -52081
rect 108496 -52181 109305 -52137
rect 109349 -52181 109405 -52137
rect 109449 -52181 109505 -52137
rect 109549 -52181 109605 -52137
rect 109649 -52181 109705 -52137
rect 109749 -52181 109805 -52137
rect 109849 -52181 109905 -52137
rect 109949 -52181 110005 -52137
rect 110049 -52181 110105 -52137
rect 110149 -52181 110205 -52137
rect 110249 -52181 110305 -52137
rect 110349 -52181 110405 -52137
rect 110449 -52181 110505 -52137
rect 110549 -52181 110605 -52137
rect 110649 -52181 110705 -52137
rect 110749 -52181 110805 -52137
rect 110849 -52181 111305 -52137
rect 111349 -52181 111405 -52137
rect 111449 -52181 111505 -52137
rect 111549 -52181 111605 -52137
rect 111649 -52181 111705 -52137
rect 111749 -52181 111805 -52137
rect 111849 -52181 111905 -52137
rect 111949 -52181 112005 -52137
rect 112049 -52181 112105 -52137
rect 112149 -52181 112205 -52137
rect 112249 -52181 112305 -52137
rect 112349 -52181 112405 -52137
rect 112449 -52181 112505 -52137
rect 112549 -52181 112605 -52137
rect 112649 -52181 112705 -52137
rect 112749 -52181 112805 -52137
rect 112849 -52181 113305 -52137
rect 113349 -52181 113405 -52137
rect 113449 -52181 113505 -52137
rect 113549 -52181 113605 -52137
rect 113649 -52181 113705 -52137
rect 113749 -52181 113805 -52137
rect 113849 -52181 113905 -52137
rect 113949 -52181 114005 -52137
rect 114049 -52181 114105 -52137
rect 114149 -52181 114205 -52137
rect 114249 -52181 114305 -52137
rect 114349 -52181 114405 -52137
rect 114449 -52181 114505 -52137
rect 114549 -52181 114605 -52137
rect 114649 -52181 114705 -52137
rect 114749 -52181 114805 -52137
rect 114849 -52181 115305 -52137
rect 115349 -52181 115405 -52137
rect 115449 -52181 115505 -52137
rect 115549 -52181 115605 -52137
rect 115649 -52181 115705 -52137
rect 115749 -52181 115805 -52137
rect 115849 -52181 115905 -52137
rect 115949 -52181 116005 -52137
rect 116049 -52181 116105 -52137
rect 116149 -52181 116205 -52137
rect 116249 -52181 116305 -52137
rect 116349 -52181 116405 -52137
rect 116449 -52181 116505 -52137
rect 116549 -52181 116605 -52137
rect 116649 -52181 116705 -52137
rect 116749 -52181 116805 -52137
rect 116849 -52181 117196 -52137
rect 108496 -52237 117196 -52181
rect 108496 -52281 109305 -52237
rect 109349 -52281 109405 -52237
rect 109449 -52281 109505 -52237
rect 109549 -52281 109605 -52237
rect 109649 -52281 109705 -52237
rect 109749 -52281 109805 -52237
rect 109849 -52281 109905 -52237
rect 109949 -52281 110005 -52237
rect 110049 -52281 110105 -52237
rect 110149 -52281 110205 -52237
rect 110249 -52281 110305 -52237
rect 110349 -52281 110405 -52237
rect 110449 -52281 110505 -52237
rect 110549 -52281 110605 -52237
rect 110649 -52281 110705 -52237
rect 110749 -52281 110805 -52237
rect 110849 -52281 111305 -52237
rect 111349 -52281 111405 -52237
rect 111449 -52281 111505 -52237
rect 111549 -52281 111605 -52237
rect 111649 -52281 111705 -52237
rect 111749 -52281 111805 -52237
rect 111849 -52281 111905 -52237
rect 111949 -52281 112005 -52237
rect 112049 -52281 112105 -52237
rect 112149 -52281 112205 -52237
rect 112249 -52281 112305 -52237
rect 112349 -52281 112405 -52237
rect 112449 -52281 112505 -52237
rect 112549 -52281 112605 -52237
rect 112649 -52281 112705 -52237
rect 112749 -52281 112805 -52237
rect 112849 -52281 113305 -52237
rect 113349 -52281 113405 -52237
rect 113449 -52281 113505 -52237
rect 113549 -52281 113605 -52237
rect 113649 -52281 113705 -52237
rect 113749 -52281 113805 -52237
rect 113849 -52281 113905 -52237
rect 113949 -52281 114005 -52237
rect 114049 -52281 114105 -52237
rect 114149 -52281 114205 -52237
rect 114249 -52281 114305 -52237
rect 114349 -52281 114405 -52237
rect 114449 -52281 114505 -52237
rect 114549 -52281 114605 -52237
rect 114649 -52281 114705 -52237
rect 114749 -52281 114805 -52237
rect 114849 -52281 115305 -52237
rect 115349 -52281 115405 -52237
rect 115449 -52281 115505 -52237
rect 115549 -52281 115605 -52237
rect 115649 -52281 115705 -52237
rect 115749 -52281 115805 -52237
rect 115849 -52281 115905 -52237
rect 115949 -52281 116005 -52237
rect 116049 -52281 116105 -52237
rect 116149 -52281 116205 -52237
rect 116249 -52281 116305 -52237
rect 116349 -52281 116405 -52237
rect 116449 -52281 116505 -52237
rect 116549 -52281 116605 -52237
rect 116649 -52281 116705 -52237
rect 116749 -52281 116805 -52237
rect 116849 -52281 117196 -52237
rect 108496 -52337 117196 -52281
rect 108496 -52381 109305 -52337
rect 109349 -52381 109405 -52337
rect 109449 -52381 109505 -52337
rect 109549 -52381 109605 -52337
rect 109649 -52381 109705 -52337
rect 109749 -52381 109805 -52337
rect 109849 -52381 109905 -52337
rect 109949 -52381 110005 -52337
rect 110049 -52381 110105 -52337
rect 110149 -52381 110205 -52337
rect 110249 -52381 110305 -52337
rect 110349 -52381 110405 -52337
rect 110449 -52381 110505 -52337
rect 110549 -52381 110605 -52337
rect 110649 -52381 110705 -52337
rect 110749 -52381 110805 -52337
rect 110849 -52381 111305 -52337
rect 111349 -52381 111405 -52337
rect 111449 -52381 111505 -52337
rect 111549 -52381 111605 -52337
rect 111649 -52381 111705 -52337
rect 111749 -52381 111805 -52337
rect 111849 -52381 111905 -52337
rect 111949 -52381 112005 -52337
rect 112049 -52381 112105 -52337
rect 112149 -52381 112205 -52337
rect 112249 -52381 112305 -52337
rect 112349 -52381 112405 -52337
rect 112449 -52381 112505 -52337
rect 112549 -52381 112605 -52337
rect 112649 -52381 112705 -52337
rect 112749 -52381 112805 -52337
rect 112849 -52381 113305 -52337
rect 113349 -52381 113405 -52337
rect 113449 -52381 113505 -52337
rect 113549 -52381 113605 -52337
rect 113649 -52381 113705 -52337
rect 113749 -52381 113805 -52337
rect 113849 -52381 113905 -52337
rect 113949 -52381 114005 -52337
rect 114049 -52381 114105 -52337
rect 114149 -52381 114205 -52337
rect 114249 -52381 114305 -52337
rect 114349 -52381 114405 -52337
rect 114449 -52381 114505 -52337
rect 114549 -52381 114605 -52337
rect 114649 -52381 114705 -52337
rect 114749 -52381 114805 -52337
rect 114849 -52381 115305 -52337
rect 115349 -52381 115405 -52337
rect 115449 -52381 115505 -52337
rect 115549 -52381 115605 -52337
rect 115649 -52381 115705 -52337
rect 115749 -52381 115805 -52337
rect 115849 -52381 115905 -52337
rect 115949 -52381 116005 -52337
rect 116049 -52381 116105 -52337
rect 116149 -52381 116205 -52337
rect 116249 -52381 116305 -52337
rect 116349 -52381 116405 -52337
rect 116449 -52381 116505 -52337
rect 116549 -52381 116605 -52337
rect 116649 -52381 116705 -52337
rect 116749 -52381 116805 -52337
rect 116849 -52381 117196 -52337
rect 108496 -52437 117196 -52381
rect 108496 -52481 109305 -52437
rect 109349 -52481 109405 -52437
rect 109449 -52481 109505 -52437
rect 109549 -52481 109605 -52437
rect 109649 -52481 109705 -52437
rect 109749 -52481 109805 -52437
rect 109849 -52481 109905 -52437
rect 109949 -52481 110005 -52437
rect 110049 -52481 110105 -52437
rect 110149 -52481 110205 -52437
rect 110249 -52481 110305 -52437
rect 110349 -52481 110405 -52437
rect 110449 -52481 110505 -52437
rect 110549 -52481 110605 -52437
rect 110649 -52481 110705 -52437
rect 110749 -52481 110805 -52437
rect 110849 -52481 111305 -52437
rect 111349 -52481 111405 -52437
rect 111449 -52481 111505 -52437
rect 111549 -52481 111605 -52437
rect 111649 -52481 111705 -52437
rect 111749 -52481 111805 -52437
rect 111849 -52481 111905 -52437
rect 111949 -52481 112005 -52437
rect 112049 -52481 112105 -52437
rect 112149 -52481 112205 -52437
rect 112249 -52481 112305 -52437
rect 112349 -52481 112405 -52437
rect 112449 -52481 112505 -52437
rect 112549 -52481 112605 -52437
rect 112649 -52481 112705 -52437
rect 112749 -52481 112805 -52437
rect 112849 -52481 113305 -52437
rect 113349 -52481 113405 -52437
rect 113449 -52481 113505 -52437
rect 113549 -52481 113605 -52437
rect 113649 -52481 113705 -52437
rect 113749 -52481 113805 -52437
rect 113849 -52481 113905 -52437
rect 113949 -52481 114005 -52437
rect 114049 -52481 114105 -52437
rect 114149 -52481 114205 -52437
rect 114249 -52481 114305 -52437
rect 114349 -52481 114405 -52437
rect 114449 -52481 114505 -52437
rect 114549 -52481 114605 -52437
rect 114649 -52481 114705 -52437
rect 114749 -52481 114805 -52437
rect 114849 -52481 115305 -52437
rect 115349 -52481 115405 -52437
rect 115449 -52481 115505 -52437
rect 115549 -52481 115605 -52437
rect 115649 -52481 115705 -52437
rect 115749 -52481 115805 -52437
rect 115849 -52481 115905 -52437
rect 115949 -52481 116005 -52437
rect 116049 -52481 116105 -52437
rect 116149 -52481 116205 -52437
rect 116249 -52481 116305 -52437
rect 116349 -52481 116405 -52437
rect 116449 -52481 116505 -52437
rect 116549 -52481 116605 -52437
rect 116649 -52481 116705 -52437
rect 116749 -52481 116805 -52437
rect 116849 -52481 117196 -52437
rect 108496 -52537 117196 -52481
rect 108496 -52581 109305 -52537
rect 109349 -52581 109405 -52537
rect 109449 -52581 109505 -52537
rect 109549 -52581 109605 -52537
rect 109649 -52581 109705 -52537
rect 109749 -52581 109805 -52537
rect 109849 -52581 109905 -52537
rect 109949 -52581 110005 -52537
rect 110049 -52581 110105 -52537
rect 110149 -52581 110205 -52537
rect 110249 -52581 110305 -52537
rect 110349 -52581 110405 -52537
rect 110449 -52581 110505 -52537
rect 110549 -52581 110605 -52537
rect 110649 -52581 110705 -52537
rect 110749 -52581 110805 -52537
rect 110849 -52581 111305 -52537
rect 111349 -52581 111405 -52537
rect 111449 -52581 111505 -52537
rect 111549 -52581 111605 -52537
rect 111649 -52581 111705 -52537
rect 111749 -52581 111805 -52537
rect 111849 -52581 111905 -52537
rect 111949 -52581 112005 -52537
rect 112049 -52581 112105 -52537
rect 112149 -52581 112205 -52537
rect 112249 -52581 112305 -52537
rect 112349 -52581 112405 -52537
rect 112449 -52581 112505 -52537
rect 112549 -52581 112605 -52537
rect 112649 -52581 112705 -52537
rect 112749 -52581 112805 -52537
rect 112849 -52581 113305 -52537
rect 113349 -52581 113405 -52537
rect 113449 -52581 113505 -52537
rect 113549 -52581 113605 -52537
rect 113649 -52581 113705 -52537
rect 113749 -52581 113805 -52537
rect 113849 -52581 113905 -52537
rect 113949 -52581 114005 -52537
rect 114049 -52581 114105 -52537
rect 114149 -52581 114205 -52537
rect 114249 -52581 114305 -52537
rect 114349 -52581 114405 -52537
rect 114449 -52581 114505 -52537
rect 114549 -52581 114605 -52537
rect 114649 -52581 114705 -52537
rect 114749 -52581 114805 -52537
rect 114849 -52581 115305 -52537
rect 115349 -52581 115405 -52537
rect 115449 -52581 115505 -52537
rect 115549 -52581 115605 -52537
rect 115649 -52581 115705 -52537
rect 115749 -52581 115805 -52537
rect 115849 -52581 115905 -52537
rect 115949 -52581 116005 -52537
rect 116049 -52581 116105 -52537
rect 116149 -52581 116205 -52537
rect 116249 -52581 116305 -52537
rect 116349 -52581 116405 -52537
rect 116449 -52581 116505 -52537
rect 116549 -52581 116605 -52537
rect 116649 -52581 116705 -52537
rect 116749 -52581 116805 -52537
rect 116849 -52581 117196 -52537
rect 108496 -52637 117196 -52581
rect 108496 -52681 109305 -52637
rect 109349 -52681 109405 -52637
rect 109449 -52681 109505 -52637
rect 109549 -52681 109605 -52637
rect 109649 -52681 109705 -52637
rect 109749 -52681 109805 -52637
rect 109849 -52681 109905 -52637
rect 109949 -52681 110005 -52637
rect 110049 -52681 110105 -52637
rect 110149 -52681 110205 -52637
rect 110249 -52681 110305 -52637
rect 110349 -52681 110405 -52637
rect 110449 -52681 110505 -52637
rect 110549 -52681 110605 -52637
rect 110649 -52681 110705 -52637
rect 110749 -52681 110805 -52637
rect 110849 -52681 111305 -52637
rect 111349 -52681 111405 -52637
rect 111449 -52681 111505 -52637
rect 111549 -52681 111605 -52637
rect 111649 -52681 111705 -52637
rect 111749 -52681 111805 -52637
rect 111849 -52681 111905 -52637
rect 111949 -52681 112005 -52637
rect 112049 -52681 112105 -52637
rect 112149 -52681 112205 -52637
rect 112249 -52681 112305 -52637
rect 112349 -52681 112405 -52637
rect 112449 -52681 112505 -52637
rect 112549 -52681 112605 -52637
rect 112649 -52681 112705 -52637
rect 112749 -52681 112805 -52637
rect 112849 -52681 113305 -52637
rect 113349 -52681 113405 -52637
rect 113449 -52681 113505 -52637
rect 113549 -52681 113605 -52637
rect 113649 -52681 113705 -52637
rect 113749 -52681 113805 -52637
rect 113849 -52681 113905 -52637
rect 113949 -52681 114005 -52637
rect 114049 -52681 114105 -52637
rect 114149 -52681 114205 -52637
rect 114249 -52681 114305 -52637
rect 114349 -52681 114405 -52637
rect 114449 -52681 114505 -52637
rect 114549 -52681 114605 -52637
rect 114649 -52681 114705 -52637
rect 114749 -52681 114805 -52637
rect 114849 -52681 115305 -52637
rect 115349 -52681 115405 -52637
rect 115449 -52681 115505 -52637
rect 115549 -52681 115605 -52637
rect 115649 -52681 115705 -52637
rect 115749 -52681 115805 -52637
rect 115849 -52681 115905 -52637
rect 115949 -52681 116005 -52637
rect 116049 -52681 116105 -52637
rect 116149 -52681 116205 -52637
rect 116249 -52681 116305 -52637
rect 116349 -52681 116405 -52637
rect 116449 -52681 116505 -52637
rect 116549 -52681 116605 -52637
rect 116649 -52681 116705 -52637
rect 116749 -52681 116805 -52637
rect 116849 -52681 117196 -52637
rect 108496 -54119 117196 -52681
rect 79796 -80499 80737 -80455
rect 80781 -80499 80837 -80455
rect 80881 -80499 80937 -80455
rect 80981 -80499 81037 -80455
rect 81081 -80499 81137 -80455
rect 81181 -80499 81237 -80455
rect 81281 -80499 81337 -80455
rect 81381 -80499 81437 -80455
rect 81481 -80499 81537 -80455
rect 81581 -80499 81637 -80455
rect 81681 -80499 81737 -80455
rect 81781 -80499 81837 -80455
rect 81881 -80499 81937 -80455
rect 81981 -80499 82037 -80455
rect 82081 -80499 82137 -80455
rect 82181 -80499 82237 -80455
rect 82281 -80499 82737 -80455
rect 82781 -80499 82837 -80455
rect 82881 -80499 82937 -80455
rect 82981 -80499 83037 -80455
rect 83081 -80499 83137 -80455
rect 83181 -80499 83237 -80455
rect 83281 -80499 83337 -80455
rect 83381 -80499 83437 -80455
rect 83481 -80499 83537 -80455
rect 83581 -80499 83637 -80455
rect 83681 -80499 83737 -80455
rect 83781 -80499 83837 -80455
rect 83881 -80499 83937 -80455
rect 83981 -80499 84037 -80455
rect 84081 -80499 84137 -80455
rect 84181 -80499 84237 -80455
rect 84281 -80499 84737 -80455
rect 84781 -80499 84837 -80455
rect 84881 -80499 84937 -80455
rect 84981 -80499 85037 -80455
rect 85081 -80499 85137 -80455
rect 85181 -80499 85237 -80455
rect 85281 -80499 85337 -80455
rect 85381 -80499 85437 -80455
rect 85481 -80499 85537 -80455
rect 85581 -80499 85637 -80455
rect 85681 -80499 85737 -80455
rect 85781 -80499 85837 -80455
rect 85881 -80499 85937 -80455
rect 85981 -80499 86037 -80455
rect 86081 -80499 86137 -80455
rect 86181 -80499 86237 -80455
rect 86281 -80499 86737 -80455
rect 86781 -80499 86837 -80455
rect 86881 -80499 86937 -80455
rect 86981 -80499 87037 -80455
rect 87081 -80499 87137 -80455
rect 87181 -80499 87237 -80455
rect 87281 -80499 87337 -80455
rect 87381 -80499 87437 -80455
rect 87481 -80499 87537 -80455
rect 87581 -80499 87637 -80455
rect 87681 -80499 87737 -80455
rect 87781 -80499 87837 -80455
rect 87881 -80499 87937 -80455
rect 87981 -80499 88037 -80455
rect 88081 -80499 88137 -80455
rect 88181 -80499 88237 -80455
rect 88281 -80499 89254 -80455
rect 79796 -80555 89254 -80499
rect 79796 -80599 80737 -80555
rect 80781 -80599 80837 -80555
rect 80881 -80599 80937 -80555
rect 80981 -80599 81037 -80555
rect 81081 -80599 81137 -80555
rect 81181 -80599 81237 -80555
rect 81281 -80599 81337 -80555
rect 81381 -80599 81437 -80555
rect 81481 -80599 81537 -80555
rect 81581 -80599 81637 -80555
rect 81681 -80599 81737 -80555
rect 81781 -80599 81837 -80555
rect 81881 -80599 81937 -80555
rect 81981 -80599 82037 -80555
rect 82081 -80599 82137 -80555
rect 82181 -80599 82237 -80555
rect 82281 -80599 82737 -80555
rect 82781 -80599 82837 -80555
rect 82881 -80599 82937 -80555
rect 82981 -80599 83037 -80555
rect 83081 -80599 83137 -80555
rect 83181 -80599 83237 -80555
rect 83281 -80599 83337 -80555
rect 83381 -80599 83437 -80555
rect 83481 -80599 83537 -80555
rect 83581 -80599 83637 -80555
rect 83681 -80599 83737 -80555
rect 83781 -80599 83837 -80555
rect 83881 -80599 83937 -80555
rect 83981 -80599 84037 -80555
rect 84081 -80599 84137 -80555
rect 84181 -80599 84237 -80555
rect 84281 -80599 84737 -80555
rect 84781 -80599 84837 -80555
rect 84881 -80599 84937 -80555
rect 84981 -80599 85037 -80555
rect 85081 -80599 85137 -80555
rect 85181 -80599 85237 -80555
rect 85281 -80599 85337 -80555
rect 85381 -80599 85437 -80555
rect 85481 -80599 85537 -80555
rect 85581 -80599 85637 -80555
rect 85681 -80599 85737 -80555
rect 85781 -80599 85837 -80555
rect 85881 -80599 85937 -80555
rect 85981 -80599 86037 -80555
rect 86081 -80599 86137 -80555
rect 86181 -80599 86237 -80555
rect 86281 -80599 86737 -80555
rect 86781 -80599 86837 -80555
rect 86881 -80599 86937 -80555
rect 86981 -80599 87037 -80555
rect 87081 -80599 87137 -80555
rect 87181 -80599 87237 -80555
rect 87281 -80599 87337 -80555
rect 87381 -80599 87437 -80555
rect 87481 -80599 87537 -80555
rect 87581 -80599 87637 -80555
rect 87681 -80599 87737 -80555
rect 87781 -80599 87837 -80555
rect 87881 -80599 87937 -80555
rect 87981 -80599 88037 -80555
rect 88081 -80599 88137 -80555
rect 88181 -80599 88237 -80555
rect 88281 -80599 89254 -80555
rect 79796 -80655 89254 -80599
rect 79796 -80699 80737 -80655
rect 80781 -80699 80837 -80655
rect 80881 -80699 80937 -80655
rect 80981 -80699 81037 -80655
rect 81081 -80699 81137 -80655
rect 81181 -80699 81237 -80655
rect 81281 -80699 81337 -80655
rect 81381 -80699 81437 -80655
rect 81481 -80699 81537 -80655
rect 81581 -80699 81637 -80655
rect 81681 -80699 81737 -80655
rect 81781 -80699 81837 -80655
rect 81881 -80699 81937 -80655
rect 81981 -80699 82037 -80655
rect 82081 -80699 82137 -80655
rect 82181 -80699 82237 -80655
rect 82281 -80699 82737 -80655
rect 82781 -80699 82837 -80655
rect 82881 -80699 82937 -80655
rect 82981 -80699 83037 -80655
rect 83081 -80699 83137 -80655
rect 83181 -80699 83237 -80655
rect 83281 -80699 83337 -80655
rect 83381 -80699 83437 -80655
rect 83481 -80699 83537 -80655
rect 83581 -80699 83637 -80655
rect 83681 -80699 83737 -80655
rect 83781 -80699 83837 -80655
rect 83881 -80699 83937 -80655
rect 83981 -80699 84037 -80655
rect 84081 -80699 84137 -80655
rect 84181 -80699 84237 -80655
rect 84281 -80699 84737 -80655
rect 84781 -80699 84837 -80655
rect 84881 -80699 84937 -80655
rect 84981 -80699 85037 -80655
rect 85081 -80699 85137 -80655
rect 85181 -80699 85237 -80655
rect 85281 -80699 85337 -80655
rect 85381 -80699 85437 -80655
rect 85481 -80699 85537 -80655
rect 85581 -80699 85637 -80655
rect 85681 -80699 85737 -80655
rect 85781 -80699 85837 -80655
rect 85881 -80699 85937 -80655
rect 85981 -80699 86037 -80655
rect 86081 -80699 86137 -80655
rect 86181 -80699 86237 -80655
rect 86281 -80699 86737 -80655
rect 86781 -80699 86837 -80655
rect 86881 -80699 86937 -80655
rect 86981 -80699 87037 -80655
rect 87081 -80699 87137 -80655
rect 87181 -80699 87237 -80655
rect 87281 -80699 87337 -80655
rect 87381 -80699 87437 -80655
rect 87481 -80699 87537 -80655
rect 87581 -80699 87637 -80655
rect 87681 -80699 87737 -80655
rect 87781 -80699 87837 -80655
rect 87881 -80699 87937 -80655
rect 87981 -80699 88037 -80655
rect 88081 -80699 88137 -80655
rect 88181 -80699 88237 -80655
rect 88281 -80699 89254 -80655
rect 79796 -80755 89254 -80699
rect 79796 -80799 80737 -80755
rect 80781 -80799 80837 -80755
rect 80881 -80799 80937 -80755
rect 80981 -80799 81037 -80755
rect 81081 -80799 81137 -80755
rect 81181 -80799 81237 -80755
rect 81281 -80799 81337 -80755
rect 81381 -80799 81437 -80755
rect 81481 -80799 81537 -80755
rect 81581 -80799 81637 -80755
rect 81681 -80799 81737 -80755
rect 81781 -80799 81837 -80755
rect 81881 -80799 81937 -80755
rect 81981 -80799 82037 -80755
rect 82081 -80799 82137 -80755
rect 82181 -80799 82237 -80755
rect 82281 -80799 82737 -80755
rect 82781 -80799 82837 -80755
rect 82881 -80799 82937 -80755
rect 82981 -80799 83037 -80755
rect 83081 -80799 83137 -80755
rect 83181 -80799 83237 -80755
rect 83281 -80799 83337 -80755
rect 83381 -80799 83437 -80755
rect 83481 -80799 83537 -80755
rect 83581 -80799 83637 -80755
rect 83681 -80799 83737 -80755
rect 83781 -80799 83837 -80755
rect 83881 -80799 83937 -80755
rect 83981 -80799 84037 -80755
rect 84081 -80799 84137 -80755
rect 84181 -80799 84237 -80755
rect 84281 -80799 84737 -80755
rect 84781 -80799 84837 -80755
rect 84881 -80799 84937 -80755
rect 84981 -80799 85037 -80755
rect 85081 -80799 85137 -80755
rect 85181 -80799 85237 -80755
rect 85281 -80799 85337 -80755
rect 85381 -80799 85437 -80755
rect 85481 -80799 85537 -80755
rect 85581 -80799 85637 -80755
rect 85681 -80799 85737 -80755
rect 85781 -80799 85837 -80755
rect 85881 -80799 85937 -80755
rect 85981 -80799 86037 -80755
rect 86081 -80799 86137 -80755
rect 86181 -80799 86237 -80755
rect 86281 -80799 86737 -80755
rect 86781 -80799 86837 -80755
rect 86881 -80799 86937 -80755
rect 86981 -80799 87037 -80755
rect 87081 -80799 87137 -80755
rect 87181 -80799 87237 -80755
rect 87281 -80799 87337 -80755
rect 87381 -80799 87437 -80755
rect 87481 -80799 87537 -80755
rect 87581 -80799 87637 -80755
rect 87681 -80799 87737 -80755
rect 87781 -80799 87837 -80755
rect 87881 -80799 87937 -80755
rect 87981 -80799 88037 -80755
rect 88081 -80799 88137 -80755
rect 88181 -80799 88237 -80755
rect 88281 -80799 89254 -80755
rect 79796 -80855 89254 -80799
rect 79796 -80899 80737 -80855
rect 80781 -80899 80837 -80855
rect 80881 -80899 80937 -80855
rect 80981 -80899 81037 -80855
rect 81081 -80899 81137 -80855
rect 81181 -80899 81237 -80855
rect 81281 -80899 81337 -80855
rect 81381 -80899 81437 -80855
rect 81481 -80899 81537 -80855
rect 81581 -80899 81637 -80855
rect 81681 -80899 81737 -80855
rect 81781 -80899 81837 -80855
rect 81881 -80899 81937 -80855
rect 81981 -80899 82037 -80855
rect 82081 -80899 82137 -80855
rect 82181 -80899 82237 -80855
rect 82281 -80899 82737 -80855
rect 82781 -80899 82837 -80855
rect 82881 -80899 82937 -80855
rect 82981 -80899 83037 -80855
rect 83081 -80899 83137 -80855
rect 83181 -80899 83237 -80855
rect 83281 -80899 83337 -80855
rect 83381 -80899 83437 -80855
rect 83481 -80899 83537 -80855
rect 83581 -80899 83637 -80855
rect 83681 -80899 83737 -80855
rect 83781 -80899 83837 -80855
rect 83881 -80899 83937 -80855
rect 83981 -80899 84037 -80855
rect 84081 -80899 84137 -80855
rect 84181 -80899 84237 -80855
rect 84281 -80899 84737 -80855
rect 84781 -80899 84837 -80855
rect 84881 -80899 84937 -80855
rect 84981 -80899 85037 -80855
rect 85081 -80899 85137 -80855
rect 85181 -80899 85237 -80855
rect 85281 -80899 85337 -80855
rect 85381 -80899 85437 -80855
rect 85481 -80899 85537 -80855
rect 85581 -80899 85637 -80855
rect 85681 -80899 85737 -80855
rect 85781 -80899 85837 -80855
rect 85881 -80899 85937 -80855
rect 85981 -80899 86037 -80855
rect 86081 -80899 86137 -80855
rect 86181 -80899 86237 -80855
rect 86281 -80899 86737 -80855
rect 86781 -80899 86837 -80855
rect 86881 -80899 86937 -80855
rect 86981 -80899 87037 -80855
rect 87081 -80899 87137 -80855
rect 87181 -80899 87237 -80855
rect 87281 -80899 87337 -80855
rect 87381 -80899 87437 -80855
rect 87481 -80899 87537 -80855
rect 87581 -80899 87637 -80855
rect 87681 -80899 87737 -80855
rect 87781 -80899 87837 -80855
rect 87881 -80899 87937 -80855
rect 87981 -80899 88037 -80855
rect 88081 -80899 88137 -80855
rect 88181 -80899 88237 -80855
rect 88281 -80899 89254 -80855
rect 79796 -80955 89254 -80899
rect 79796 -80999 80737 -80955
rect 80781 -80999 80837 -80955
rect 80881 -80999 80937 -80955
rect 80981 -80999 81037 -80955
rect 81081 -80999 81137 -80955
rect 81181 -80999 81237 -80955
rect 81281 -80999 81337 -80955
rect 81381 -80999 81437 -80955
rect 81481 -80999 81537 -80955
rect 81581 -80999 81637 -80955
rect 81681 -80999 81737 -80955
rect 81781 -80999 81837 -80955
rect 81881 -80999 81937 -80955
rect 81981 -80999 82037 -80955
rect 82081 -80999 82137 -80955
rect 82181 -80999 82237 -80955
rect 82281 -80999 82737 -80955
rect 82781 -80999 82837 -80955
rect 82881 -80999 82937 -80955
rect 82981 -80999 83037 -80955
rect 83081 -80999 83137 -80955
rect 83181 -80999 83237 -80955
rect 83281 -80999 83337 -80955
rect 83381 -80999 83437 -80955
rect 83481 -80999 83537 -80955
rect 83581 -80999 83637 -80955
rect 83681 -80999 83737 -80955
rect 83781 -80999 83837 -80955
rect 83881 -80999 83937 -80955
rect 83981 -80999 84037 -80955
rect 84081 -80999 84137 -80955
rect 84181 -80999 84237 -80955
rect 84281 -80999 84737 -80955
rect 84781 -80999 84837 -80955
rect 84881 -80999 84937 -80955
rect 84981 -80999 85037 -80955
rect 85081 -80999 85137 -80955
rect 85181 -80999 85237 -80955
rect 85281 -80999 85337 -80955
rect 85381 -80999 85437 -80955
rect 85481 -80999 85537 -80955
rect 85581 -80999 85637 -80955
rect 85681 -80999 85737 -80955
rect 85781 -80999 85837 -80955
rect 85881 -80999 85937 -80955
rect 85981 -80999 86037 -80955
rect 86081 -80999 86137 -80955
rect 86181 -80999 86237 -80955
rect 86281 -80999 86737 -80955
rect 86781 -80999 86837 -80955
rect 86881 -80999 86937 -80955
rect 86981 -80999 87037 -80955
rect 87081 -80999 87137 -80955
rect 87181 -80999 87237 -80955
rect 87281 -80999 87337 -80955
rect 87381 -80999 87437 -80955
rect 87481 -80999 87537 -80955
rect 87581 -80999 87637 -80955
rect 87681 -80999 87737 -80955
rect 87781 -80999 87837 -80955
rect 87881 -80999 87937 -80955
rect 87981 -80999 88037 -80955
rect 88081 -80999 88137 -80955
rect 88181 -80999 88237 -80955
rect 88281 -80999 89254 -80955
rect 79796 -81055 89254 -80999
rect 79796 -81099 80737 -81055
rect 80781 -81099 80837 -81055
rect 80881 -81099 80937 -81055
rect 80981 -81099 81037 -81055
rect 81081 -81099 81137 -81055
rect 81181 -81099 81237 -81055
rect 81281 -81099 81337 -81055
rect 81381 -81099 81437 -81055
rect 81481 -81099 81537 -81055
rect 81581 -81099 81637 -81055
rect 81681 -81099 81737 -81055
rect 81781 -81099 81837 -81055
rect 81881 -81099 81937 -81055
rect 81981 -81099 82037 -81055
rect 82081 -81099 82137 -81055
rect 82181 -81099 82237 -81055
rect 82281 -81099 82737 -81055
rect 82781 -81099 82837 -81055
rect 82881 -81099 82937 -81055
rect 82981 -81099 83037 -81055
rect 83081 -81099 83137 -81055
rect 83181 -81099 83237 -81055
rect 83281 -81099 83337 -81055
rect 83381 -81099 83437 -81055
rect 83481 -81099 83537 -81055
rect 83581 -81099 83637 -81055
rect 83681 -81099 83737 -81055
rect 83781 -81099 83837 -81055
rect 83881 -81099 83937 -81055
rect 83981 -81099 84037 -81055
rect 84081 -81099 84137 -81055
rect 84181 -81099 84237 -81055
rect 84281 -81099 84737 -81055
rect 84781 -81099 84837 -81055
rect 84881 -81099 84937 -81055
rect 84981 -81099 85037 -81055
rect 85081 -81099 85137 -81055
rect 85181 -81099 85237 -81055
rect 85281 -81099 85337 -81055
rect 85381 -81099 85437 -81055
rect 85481 -81099 85537 -81055
rect 85581 -81099 85637 -81055
rect 85681 -81099 85737 -81055
rect 85781 -81099 85837 -81055
rect 85881 -81099 85937 -81055
rect 85981 -81099 86037 -81055
rect 86081 -81099 86137 -81055
rect 86181 -81099 86237 -81055
rect 86281 -81099 86737 -81055
rect 86781 -81099 86837 -81055
rect 86881 -81099 86937 -81055
rect 86981 -81099 87037 -81055
rect 87081 -81099 87137 -81055
rect 87181 -81099 87237 -81055
rect 87281 -81099 87337 -81055
rect 87381 -81099 87437 -81055
rect 87481 -81099 87537 -81055
rect 87581 -81099 87637 -81055
rect 87681 -81099 87737 -81055
rect 87781 -81099 87837 -81055
rect 87881 -81099 87937 -81055
rect 87981 -81099 88037 -81055
rect 88081 -81099 88137 -81055
rect 88181 -81099 88237 -81055
rect 88281 -81099 89254 -81055
rect 79796 -81155 89254 -81099
rect 79796 -81199 80737 -81155
rect 80781 -81199 80837 -81155
rect 80881 -81199 80937 -81155
rect 80981 -81199 81037 -81155
rect 81081 -81199 81137 -81155
rect 81181 -81199 81237 -81155
rect 81281 -81199 81337 -81155
rect 81381 -81199 81437 -81155
rect 81481 -81199 81537 -81155
rect 81581 -81199 81637 -81155
rect 81681 -81199 81737 -81155
rect 81781 -81199 81837 -81155
rect 81881 -81199 81937 -81155
rect 81981 -81199 82037 -81155
rect 82081 -81199 82137 -81155
rect 82181 -81199 82237 -81155
rect 82281 -81199 82737 -81155
rect 82781 -81199 82837 -81155
rect 82881 -81199 82937 -81155
rect 82981 -81199 83037 -81155
rect 83081 -81199 83137 -81155
rect 83181 -81199 83237 -81155
rect 83281 -81199 83337 -81155
rect 83381 -81199 83437 -81155
rect 83481 -81199 83537 -81155
rect 83581 -81199 83637 -81155
rect 83681 -81199 83737 -81155
rect 83781 -81199 83837 -81155
rect 83881 -81199 83937 -81155
rect 83981 -81199 84037 -81155
rect 84081 -81199 84137 -81155
rect 84181 -81199 84237 -81155
rect 84281 -81199 84737 -81155
rect 84781 -81199 84837 -81155
rect 84881 -81199 84937 -81155
rect 84981 -81199 85037 -81155
rect 85081 -81199 85137 -81155
rect 85181 -81199 85237 -81155
rect 85281 -81199 85337 -81155
rect 85381 -81199 85437 -81155
rect 85481 -81199 85537 -81155
rect 85581 -81199 85637 -81155
rect 85681 -81199 85737 -81155
rect 85781 -81199 85837 -81155
rect 85881 -81199 85937 -81155
rect 85981 -81199 86037 -81155
rect 86081 -81199 86137 -81155
rect 86181 -81199 86237 -81155
rect 86281 -81199 86737 -81155
rect 86781 -81199 86837 -81155
rect 86881 -81199 86937 -81155
rect 86981 -81199 87037 -81155
rect 87081 -81199 87137 -81155
rect 87181 -81199 87237 -81155
rect 87281 -81199 87337 -81155
rect 87381 -81199 87437 -81155
rect 87481 -81199 87537 -81155
rect 87581 -81199 87637 -81155
rect 87681 -81199 87737 -81155
rect 87781 -81199 87837 -81155
rect 87881 -81199 87937 -81155
rect 87981 -81199 88037 -81155
rect 88081 -81199 88137 -81155
rect 88181 -81199 88237 -81155
rect 88281 -81199 89254 -81155
rect 79796 -81255 89254 -81199
rect 79796 -81299 80737 -81255
rect 80781 -81299 80837 -81255
rect 80881 -81299 80937 -81255
rect 80981 -81299 81037 -81255
rect 81081 -81299 81137 -81255
rect 81181 -81299 81237 -81255
rect 81281 -81299 81337 -81255
rect 81381 -81299 81437 -81255
rect 81481 -81299 81537 -81255
rect 81581 -81299 81637 -81255
rect 81681 -81299 81737 -81255
rect 81781 -81299 81837 -81255
rect 81881 -81299 81937 -81255
rect 81981 -81299 82037 -81255
rect 82081 -81299 82137 -81255
rect 82181 -81299 82237 -81255
rect 82281 -81299 82737 -81255
rect 82781 -81299 82837 -81255
rect 82881 -81299 82937 -81255
rect 82981 -81299 83037 -81255
rect 83081 -81299 83137 -81255
rect 83181 -81299 83237 -81255
rect 83281 -81299 83337 -81255
rect 83381 -81299 83437 -81255
rect 83481 -81299 83537 -81255
rect 83581 -81299 83637 -81255
rect 83681 -81299 83737 -81255
rect 83781 -81299 83837 -81255
rect 83881 -81299 83937 -81255
rect 83981 -81299 84037 -81255
rect 84081 -81299 84137 -81255
rect 84181 -81299 84237 -81255
rect 84281 -81299 84737 -81255
rect 84781 -81299 84837 -81255
rect 84881 -81299 84937 -81255
rect 84981 -81299 85037 -81255
rect 85081 -81299 85137 -81255
rect 85181 -81299 85237 -81255
rect 85281 -81299 85337 -81255
rect 85381 -81299 85437 -81255
rect 85481 -81299 85537 -81255
rect 85581 -81299 85637 -81255
rect 85681 -81299 85737 -81255
rect 85781 -81299 85837 -81255
rect 85881 -81299 85937 -81255
rect 85981 -81299 86037 -81255
rect 86081 -81299 86137 -81255
rect 86181 -81299 86237 -81255
rect 86281 -81299 86737 -81255
rect 86781 -81299 86837 -81255
rect 86881 -81299 86937 -81255
rect 86981 -81299 87037 -81255
rect 87081 -81299 87137 -81255
rect 87181 -81299 87237 -81255
rect 87281 -81299 87337 -81255
rect 87381 -81299 87437 -81255
rect 87481 -81299 87537 -81255
rect 87581 -81299 87637 -81255
rect 87681 -81299 87737 -81255
rect 87781 -81299 87837 -81255
rect 87881 -81299 87937 -81255
rect 87981 -81299 88037 -81255
rect 88081 -81299 88137 -81255
rect 88181 -81299 88237 -81255
rect 88281 -81299 89254 -81255
rect 79796 -81355 89254 -81299
rect 79796 -81399 80737 -81355
rect 80781 -81399 80837 -81355
rect 80881 -81399 80937 -81355
rect 80981 -81399 81037 -81355
rect 81081 -81399 81137 -81355
rect 81181 -81399 81237 -81355
rect 81281 -81399 81337 -81355
rect 81381 -81399 81437 -81355
rect 81481 -81399 81537 -81355
rect 81581 -81399 81637 -81355
rect 81681 -81399 81737 -81355
rect 81781 -81399 81837 -81355
rect 81881 -81399 81937 -81355
rect 81981 -81399 82037 -81355
rect 82081 -81399 82137 -81355
rect 82181 -81399 82237 -81355
rect 82281 -81399 82737 -81355
rect 82781 -81399 82837 -81355
rect 82881 -81399 82937 -81355
rect 82981 -81399 83037 -81355
rect 83081 -81399 83137 -81355
rect 83181 -81399 83237 -81355
rect 83281 -81399 83337 -81355
rect 83381 -81399 83437 -81355
rect 83481 -81399 83537 -81355
rect 83581 -81399 83637 -81355
rect 83681 -81399 83737 -81355
rect 83781 -81399 83837 -81355
rect 83881 -81399 83937 -81355
rect 83981 -81399 84037 -81355
rect 84081 -81399 84137 -81355
rect 84181 -81399 84237 -81355
rect 84281 -81399 84737 -81355
rect 84781 -81399 84837 -81355
rect 84881 -81399 84937 -81355
rect 84981 -81399 85037 -81355
rect 85081 -81399 85137 -81355
rect 85181 -81399 85237 -81355
rect 85281 -81399 85337 -81355
rect 85381 -81399 85437 -81355
rect 85481 -81399 85537 -81355
rect 85581 -81399 85637 -81355
rect 85681 -81399 85737 -81355
rect 85781 -81399 85837 -81355
rect 85881 -81399 85937 -81355
rect 85981 -81399 86037 -81355
rect 86081 -81399 86137 -81355
rect 86181 -81399 86237 -81355
rect 86281 -81399 86737 -81355
rect 86781 -81399 86837 -81355
rect 86881 -81399 86937 -81355
rect 86981 -81399 87037 -81355
rect 87081 -81399 87137 -81355
rect 87181 -81399 87237 -81355
rect 87281 -81399 87337 -81355
rect 87381 -81399 87437 -81355
rect 87481 -81399 87537 -81355
rect 87581 -81399 87637 -81355
rect 87681 -81399 87737 -81355
rect 87781 -81399 87837 -81355
rect 87881 -81399 87937 -81355
rect 87981 -81399 88037 -81355
rect 88081 -81399 88137 -81355
rect 88181 -81399 88237 -81355
rect 88281 -81399 89254 -81355
rect 79796 -81455 89254 -81399
rect 79796 -81499 80737 -81455
rect 80781 -81499 80837 -81455
rect 80881 -81499 80937 -81455
rect 80981 -81499 81037 -81455
rect 81081 -81499 81137 -81455
rect 81181 -81499 81237 -81455
rect 81281 -81499 81337 -81455
rect 81381 -81499 81437 -81455
rect 81481 -81499 81537 -81455
rect 81581 -81499 81637 -81455
rect 81681 -81499 81737 -81455
rect 81781 -81499 81837 -81455
rect 81881 -81499 81937 -81455
rect 81981 -81499 82037 -81455
rect 82081 -81499 82137 -81455
rect 82181 -81499 82237 -81455
rect 82281 -81499 82737 -81455
rect 82781 -81499 82837 -81455
rect 82881 -81499 82937 -81455
rect 82981 -81499 83037 -81455
rect 83081 -81499 83137 -81455
rect 83181 -81499 83237 -81455
rect 83281 -81499 83337 -81455
rect 83381 -81499 83437 -81455
rect 83481 -81499 83537 -81455
rect 83581 -81499 83637 -81455
rect 83681 -81499 83737 -81455
rect 83781 -81499 83837 -81455
rect 83881 -81499 83937 -81455
rect 83981 -81499 84037 -81455
rect 84081 -81499 84137 -81455
rect 84181 -81499 84237 -81455
rect 84281 -81499 84737 -81455
rect 84781 -81499 84837 -81455
rect 84881 -81499 84937 -81455
rect 84981 -81499 85037 -81455
rect 85081 -81499 85137 -81455
rect 85181 -81499 85237 -81455
rect 85281 -81499 85337 -81455
rect 85381 -81499 85437 -81455
rect 85481 -81499 85537 -81455
rect 85581 -81499 85637 -81455
rect 85681 -81499 85737 -81455
rect 85781 -81499 85837 -81455
rect 85881 -81499 85937 -81455
rect 85981 -81499 86037 -81455
rect 86081 -81499 86137 -81455
rect 86181 -81499 86237 -81455
rect 86281 -81499 86737 -81455
rect 86781 -81499 86837 -81455
rect 86881 -81499 86937 -81455
rect 86981 -81499 87037 -81455
rect 87081 -81499 87137 -81455
rect 87181 -81499 87237 -81455
rect 87281 -81499 87337 -81455
rect 87381 -81499 87437 -81455
rect 87481 -81499 87537 -81455
rect 87581 -81499 87637 -81455
rect 87681 -81499 87737 -81455
rect 87781 -81499 87837 -81455
rect 87881 -81499 87937 -81455
rect 87981 -81499 88037 -81455
rect 88081 -81499 88137 -81455
rect 88181 -81499 88237 -81455
rect 88281 -81499 89254 -81455
rect 79796 -81555 89254 -81499
rect 79796 -81599 80737 -81555
rect 80781 -81599 80837 -81555
rect 80881 -81599 80937 -81555
rect 80981 -81599 81037 -81555
rect 81081 -81599 81137 -81555
rect 81181 -81599 81237 -81555
rect 81281 -81599 81337 -81555
rect 81381 -81599 81437 -81555
rect 81481 -81599 81537 -81555
rect 81581 -81599 81637 -81555
rect 81681 -81599 81737 -81555
rect 81781 -81599 81837 -81555
rect 81881 -81599 81937 -81555
rect 81981 -81599 82037 -81555
rect 82081 -81599 82137 -81555
rect 82181 -81599 82237 -81555
rect 82281 -81599 82737 -81555
rect 82781 -81599 82837 -81555
rect 82881 -81599 82937 -81555
rect 82981 -81599 83037 -81555
rect 83081 -81599 83137 -81555
rect 83181 -81599 83237 -81555
rect 83281 -81599 83337 -81555
rect 83381 -81599 83437 -81555
rect 83481 -81599 83537 -81555
rect 83581 -81599 83637 -81555
rect 83681 -81599 83737 -81555
rect 83781 -81599 83837 -81555
rect 83881 -81599 83937 -81555
rect 83981 -81599 84037 -81555
rect 84081 -81599 84137 -81555
rect 84181 -81599 84237 -81555
rect 84281 -81599 84737 -81555
rect 84781 -81599 84837 -81555
rect 84881 -81599 84937 -81555
rect 84981 -81599 85037 -81555
rect 85081 -81599 85137 -81555
rect 85181 -81599 85237 -81555
rect 85281 -81599 85337 -81555
rect 85381 -81599 85437 -81555
rect 85481 -81599 85537 -81555
rect 85581 -81599 85637 -81555
rect 85681 -81599 85737 -81555
rect 85781 -81599 85837 -81555
rect 85881 -81599 85937 -81555
rect 85981 -81599 86037 -81555
rect 86081 -81599 86137 -81555
rect 86181 -81599 86237 -81555
rect 86281 -81599 86737 -81555
rect 86781 -81599 86837 -81555
rect 86881 -81599 86937 -81555
rect 86981 -81599 87037 -81555
rect 87081 -81599 87137 -81555
rect 87181 -81599 87237 -81555
rect 87281 -81599 87337 -81555
rect 87381 -81599 87437 -81555
rect 87481 -81599 87537 -81555
rect 87581 -81599 87637 -81555
rect 87681 -81599 87737 -81555
rect 87781 -81599 87837 -81555
rect 87881 -81599 87937 -81555
rect 87981 -81599 88037 -81555
rect 88081 -81599 88137 -81555
rect 88181 -81599 88237 -81555
rect 88281 -81599 89254 -81555
rect 79796 -81655 89254 -81599
rect 79796 -81699 80737 -81655
rect 80781 -81699 80837 -81655
rect 80881 -81699 80937 -81655
rect 80981 -81699 81037 -81655
rect 81081 -81699 81137 -81655
rect 81181 -81699 81237 -81655
rect 81281 -81699 81337 -81655
rect 81381 -81699 81437 -81655
rect 81481 -81699 81537 -81655
rect 81581 -81699 81637 -81655
rect 81681 -81699 81737 -81655
rect 81781 -81699 81837 -81655
rect 81881 -81699 81937 -81655
rect 81981 -81699 82037 -81655
rect 82081 -81699 82137 -81655
rect 82181 -81699 82237 -81655
rect 82281 -81699 82737 -81655
rect 82781 -81699 82837 -81655
rect 82881 -81699 82937 -81655
rect 82981 -81699 83037 -81655
rect 83081 -81699 83137 -81655
rect 83181 -81699 83237 -81655
rect 83281 -81699 83337 -81655
rect 83381 -81699 83437 -81655
rect 83481 -81699 83537 -81655
rect 83581 -81699 83637 -81655
rect 83681 -81699 83737 -81655
rect 83781 -81699 83837 -81655
rect 83881 -81699 83937 -81655
rect 83981 -81699 84037 -81655
rect 84081 -81699 84137 -81655
rect 84181 -81699 84237 -81655
rect 84281 -81699 84737 -81655
rect 84781 -81699 84837 -81655
rect 84881 -81699 84937 -81655
rect 84981 -81699 85037 -81655
rect 85081 -81699 85137 -81655
rect 85181 -81699 85237 -81655
rect 85281 -81699 85337 -81655
rect 85381 -81699 85437 -81655
rect 85481 -81699 85537 -81655
rect 85581 -81699 85637 -81655
rect 85681 -81699 85737 -81655
rect 85781 -81699 85837 -81655
rect 85881 -81699 85937 -81655
rect 85981 -81699 86037 -81655
rect 86081 -81699 86137 -81655
rect 86181 -81699 86237 -81655
rect 86281 -81699 86737 -81655
rect 86781 -81699 86837 -81655
rect 86881 -81699 86937 -81655
rect 86981 -81699 87037 -81655
rect 87081 -81699 87137 -81655
rect 87181 -81699 87237 -81655
rect 87281 -81699 87337 -81655
rect 87381 -81699 87437 -81655
rect 87481 -81699 87537 -81655
rect 87581 -81699 87637 -81655
rect 87681 -81699 87737 -81655
rect 87781 -81699 87837 -81655
rect 87881 -81699 87937 -81655
rect 87981 -81699 88037 -81655
rect 88081 -81699 88137 -81655
rect 88181 -81699 88237 -81655
rect 88281 -81699 89254 -81655
rect 79796 -81755 89254 -81699
rect 79796 -81799 80737 -81755
rect 80781 -81799 80837 -81755
rect 80881 -81799 80937 -81755
rect 80981 -81799 81037 -81755
rect 81081 -81799 81137 -81755
rect 81181 -81799 81237 -81755
rect 81281 -81799 81337 -81755
rect 81381 -81799 81437 -81755
rect 81481 -81799 81537 -81755
rect 81581 -81799 81637 -81755
rect 81681 -81799 81737 -81755
rect 81781 -81799 81837 -81755
rect 81881 -81799 81937 -81755
rect 81981 -81799 82037 -81755
rect 82081 -81799 82137 -81755
rect 82181 -81799 82237 -81755
rect 82281 -81799 82737 -81755
rect 82781 -81799 82837 -81755
rect 82881 -81799 82937 -81755
rect 82981 -81799 83037 -81755
rect 83081 -81799 83137 -81755
rect 83181 -81799 83237 -81755
rect 83281 -81799 83337 -81755
rect 83381 -81799 83437 -81755
rect 83481 -81799 83537 -81755
rect 83581 -81799 83637 -81755
rect 83681 -81799 83737 -81755
rect 83781 -81799 83837 -81755
rect 83881 -81799 83937 -81755
rect 83981 -81799 84037 -81755
rect 84081 -81799 84137 -81755
rect 84181 -81799 84237 -81755
rect 84281 -81799 84737 -81755
rect 84781 -81799 84837 -81755
rect 84881 -81799 84937 -81755
rect 84981 -81799 85037 -81755
rect 85081 -81799 85137 -81755
rect 85181 -81799 85237 -81755
rect 85281 -81799 85337 -81755
rect 85381 -81799 85437 -81755
rect 85481 -81799 85537 -81755
rect 85581 -81799 85637 -81755
rect 85681 -81799 85737 -81755
rect 85781 -81799 85837 -81755
rect 85881 -81799 85937 -81755
rect 85981 -81799 86037 -81755
rect 86081 -81799 86137 -81755
rect 86181 -81799 86237 -81755
rect 86281 -81799 86737 -81755
rect 86781 -81799 86837 -81755
rect 86881 -81799 86937 -81755
rect 86981 -81799 87037 -81755
rect 87081 -81799 87137 -81755
rect 87181 -81799 87237 -81755
rect 87281 -81799 87337 -81755
rect 87381 -81799 87437 -81755
rect 87481 -81799 87537 -81755
rect 87581 -81799 87637 -81755
rect 87681 -81799 87737 -81755
rect 87781 -81799 87837 -81755
rect 87881 -81799 87937 -81755
rect 87981 -81799 88037 -81755
rect 88081 -81799 88137 -81755
rect 88181 -81799 88237 -81755
rect 88281 -81799 89254 -81755
rect 79796 -81855 89254 -81799
rect 79796 -81899 80737 -81855
rect 80781 -81899 80837 -81855
rect 80881 -81899 80937 -81855
rect 80981 -81899 81037 -81855
rect 81081 -81899 81137 -81855
rect 81181 -81899 81237 -81855
rect 81281 -81899 81337 -81855
rect 81381 -81899 81437 -81855
rect 81481 -81899 81537 -81855
rect 81581 -81899 81637 -81855
rect 81681 -81899 81737 -81855
rect 81781 -81899 81837 -81855
rect 81881 -81899 81937 -81855
rect 81981 -81899 82037 -81855
rect 82081 -81899 82137 -81855
rect 82181 -81899 82237 -81855
rect 82281 -81899 82737 -81855
rect 82781 -81899 82837 -81855
rect 82881 -81899 82937 -81855
rect 82981 -81899 83037 -81855
rect 83081 -81899 83137 -81855
rect 83181 -81899 83237 -81855
rect 83281 -81899 83337 -81855
rect 83381 -81899 83437 -81855
rect 83481 -81899 83537 -81855
rect 83581 -81899 83637 -81855
rect 83681 -81899 83737 -81855
rect 83781 -81899 83837 -81855
rect 83881 -81899 83937 -81855
rect 83981 -81899 84037 -81855
rect 84081 -81899 84137 -81855
rect 84181 -81899 84237 -81855
rect 84281 -81899 84737 -81855
rect 84781 -81899 84837 -81855
rect 84881 -81899 84937 -81855
rect 84981 -81899 85037 -81855
rect 85081 -81899 85137 -81855
rect 85181 -81899 85237 -81855
rect 85281 -81899 85337 -81855
rect 85381 -81899 85437 -81855
rect 85481 -81899 85537 -81855
rect 85581 -81899 85637 -81855
rect 85681 -81899 85737 -81855
rect 85781 -81899 85837 -81855
rect 85881 -81899 85937 -81855
rect 85981 -81899 86037 -81855
rect 86081 -81899 86137 -81855
rect 86181 -81899 86237 -81855
rect 86281 -81899 86737 -81855
rect 86781 -81899 86837 -81855
rect 86881 -81899 86937 -81855
rect 86981 -81899 87037 -81855
rect 87081 -81899 87137 -81855
rect 87181 -81899 87237 -81855
rect 87281 -81899 87337 -81855
rect 87381 -81899 87437 -81855
rect 87481 -81899 87537 -81855
rect 87581 -81899 87637 -81855
rect 87681 -81899 87737 -81855
rect 87781 -81899 87837 -81855
rect 87881 -81899 87937 -81855
rect 87981 -81899 88037 -81855
rect 88081 -81899 88137 -81855
rect 88181 -81899 88237 -81855
rect 88281 -81899 89254 -81855
rect 79796 -81955 89254 -81899
rect 79796 -81999 80737 -81955
rect 80781 -81999 80837 -81955
rect 80881 -81999 80937 -81955
rect 80981 -81999 81037 -81955
rect 81081 -81999 81137 -81955
rect 81181 -81999 81237 -81955
rect 81281 -81999 81337 -81955
rect 81381 -81999 81437 -81955
rect 81481 -81999 81537 -81955
rect 81581 -81999 81637 -81955
rect 81681 -81999 81737 -81955
rect 81781 -81999 81837 -81955
rect 81881 -81999 81937 -81955
rect 81981 -81999 82037 -81955
rect 82081 -81999 82137 -81955
rect 82181 -81999 82237 -81955
rect 82281 -81999 82737 -81955
rect 82781 -81999 82837 -81955
rect 82881 -81999 82937 -81955
rect 82981 -81999 83037 -81955
rect 83081 -81999 83137 -81955
rect 83181 -81999 83237 -81955
rect 83281 -81999 83337 -81955
rect 83381 -81999 83437 -81955
rect 83481 -81999 83537 -81955
rect 83581 -81999 83637 -81955
rect 83681 -81999 83737 -81955
rect 83781 -81999 83837 -81955
rect 83881 -81999 83937 -81955
rect 83981 -81999 84037 -81955
rect 84081 -81999 84137 -81955
rect 84181 -81999 84237 -81955
rect 84281 -81999 84737 -81955
rect 84781 -81999 84837 -81955
rect 84881 -81999 84937 -81955
rect 84981 -81999 85037 -81955
rect 85081 -81999 85137 -81955
rect 85181 -81999 85237 -81955
rect 85281 -81999 85337 -81955
rect 85381 -81999 85437 -81955
rect 85481 -81999 85537 -81955
rect 85581 -81999 85637 -81955
rect 85681 -81999 85737 -81955
rect 85781 -81999 85837 -81955
rect 85881 -81999 85937 -81955
rect 85981 -81999 86037 -81955
rect 86081 -81999 86137 -81955
rect 86181 -81999 86237 -81955
rect 86281 -81999 86737 -81955
rect 86781 -81999 86837 -81955
rect 86881 -81999 86937 -81955
rect 86981 -81999 87037 -81955
rect 87081 -81999 87137 -81955
rect 87181 -81999 87237 -81955
rect 87281 -81999 87337 -81955
rect 87381 -81999 87437 -81955
rect 87481 -81999 87537 -81955
rect 87581 -81999 87637 -81955
rect 87681 -81999 87737 -81955
rect 87781 -81999 87837 -81955
rect 87881 -81999 87937 -81955
rect 87981 -81999 88037 -81955
rect 88081 -81999 88137 -81955
rect 88181 -81999 88237 -81955
rect 88281 -81999 89254 -81955
rect 79796 -83242 89254 -81999
rect 34207 -131429 37387 -131385
rect 37431 -131429 37487 -131385
rect 37531 -131429 37587 -131385
rect 37631 -131429 37687 -131385
rect 37731 -131429 37787 -131385
rect 37831 -131429 37887 -131385
rect 37931 -131429 37987 -131385
rect 38031 -131429 38087 -131385
rect 38131 -131429 38187 -131385
rect 38231 -131429 38287 -131385
rect 38331 -131429 38387 -131385
rect 38431 -131429 38487 -131385
rect 38531 -131429 38587 -131385
rect 38631 -131429 38687 -131385
rect 38731 -131429 38787 -131385
rect 38831 -131429 38887 -131385
rect 38931 -131429 39387 -131385
rect 39431 -131429 39487 -131385
rect 39531 -131429 39587 -131385
rect 39631 -131429 39687 -131385
rect 39731 -131429 39787 -131385
rect 39831 -131429 39887 -131385
rect 39931 -131429 39987 -131385
rect 40031 -131429 40087 -131385
rect 40131 -131429 40187 -131385
rect 40231 -131429 40287 -131385
rect 40331 -131429 40387 -131385
rect 40431 -131429 40487 -131385
rect 40531 -131429 40587 -131385
rect 40631 -131429 40687 -131385
rect 40731 -131429 40787 -131385
rect 40831 -131429 40887 -131385
rect 40931 -131429 41387 -131385
rect 41431 -131429 41487 -131385
rect 41531 -131429 41587 -131385
rect 41631 -131429 41687 -131385
rect 41731 -131429 41787 -131385
rect 41831 -131429 41887 -131385
rect 41931 -131429 41987 -131385
rect 42031 -131429 42087 -131385
rect 42131 -131429 42187 -131385
rect 42231 -131429 42287 -131385
rect 42331 -131429 42387 -131385
rect 42431 -131429 42487 -131385
rect 42531 -131429 42587 -131385
rect 42631 -131429 42687 -131385
rect 42731 -131429 42787 -131385
rect 42831 -131429 42887 -131385
rect 42931 -131429 43387 -131385
rect 43431 -131429 43487 -131385
rect 43531 -131429 43587 -131385
rect 43631 -131429 43687 -131385
rect 43731 -131429 43787 -131385
rect 43831 -131429 43887 -131385
rect 43931 -131429 43987 -131385
rect 44031 -131429 44087 -131385
rect 44131 -131429 44187 -131385
rect 44231 -131429 44287 -131385
rect 44331 -131429 44387 -131385
rect 44431 -131429 44487 -131385
rect 44531 -131429 44587 -131385
rect 44631 -131429 44687 -131385
rect 44731 -131429 44787 -131385
rect 44831 -131429 44887 -131385
rect 44931 -131429 47953 -131385
rect 34207 -131485 47953 -131429
rect 34207 -131529 37387 -131485
rect 37431 -131529 37487 -131485
rect 37531 -131529 37587 -131485
rect 37631 -131529 37687 -131485
rect 37731 -131529 37787 -131485
rect 37831 -131529 37887 -131485
rect 37931 -131529 37987 -131485
rect 38031 -131529 38087 -131485
rect 38131 -131529 38187 -131485
rect 38231 -131529 38287 -131485
rect 38331 -131529 38387 -131485
rect 38431 -131529 38487 -131485
rect 38531 -131529 38587 -131485
rect 38631 -131529 38687 -131485
rect 38731 -131529 38787 -131485
rect 38831 -131529 38887 -131485
rect 38931 -131529 39387 -131485
rect 39431 -131529 39487 -131485
rect 39531 -131529 39587 -131485
rect 39631 -131529 39687 -131485
rect 39731 -131529 39787 -131485
rect 39831 -131529 39887 -131485
rect 39931 -131529 39987 -131485
rect 40031 -131529 40087 -131485
rect 40131 -131529 40187 -131485
rect 40231 -131529 40287 -131485
rect 40331 -131529 40387 -131485
rect 40431 -131529 40487 -131485
rect 40531 -131529 40587 -131485
rect 40631 -131529 40687 -131485
rect 40731 -131529 40787 -131485
rect 40831 -131529 40887 -131485
rect 40931 -131529 41387 -131485
rect 41431 -131529 41487 -131485
rect 41531 -131529 41587 -131485
rect 41631 -131529 41687 -131485
rect 41731 -131529 41787 -131485
rect 41831 -131529 41887 -131485
rect 41931 -131529 41987 -131485
rect 42031 -131529 42087 -131485
rect 42131 -131529 42187 -131485
rect 42231 -131529 42287 -131485
rect 42331 -131529 42387 -131485
rect 42431 -131529 42487 -131485
rect 42531 -131529 42587 -131485
rect 42631 -131529 42687 -131485
rect 42731 -131529 42787 -131485
rect 42831 -131529 42887 -131485
rect 42931 -131529 43387 -131485
rect 43431 -131529 43487 -131485
rect 43531 -131529 43587 -131485
rect 43631 -131529 43687 -131485
rect 43731 -131529 43787 -131485
rect 43831 -131529 43887 -131485
rect 43931 -131529 43987 -131485
rect 44031 -131529 44087 -131485
rect 44131 -131529 44187 -131485
rect 44231 -131529 44287 -131485
rect 44331 -131529 44387 -131485
rect 44431 -131529 44487 -131485
rect 44531 -131529 44587 -131485
rect 44631 -131529 44687 -131485
rect 44731 -131529 44787 -131485
rect 44831 -131529 44887 -131485
rect 44931 -131529 47953 -131485
rect 34207 -131585 47953 -131529
rect 34207 -131629 37387 -131585
rect 37431 -131629 37487 -131585
rect 37531 -131629 37587 -131585
rect 37631 -131629 37687 -131585
rect 37731 -131629 37787 -131585
rect 37831 -131629 37887 -131585
rect 37931 -131629 37987 -131585
rect 38031 -131629 38087 -131585
rect 38131 -131629 38187 -131585
rect 38231 -131629 38287 -131585
rect 38331 -131629 38387 -131585
rect 38431 -131629 38487 -131585
rect 38531 -131629 38587 -131585
rect 38631 -131629 38687 -131585
rect 38731 -131629 38787 -131585
rect 38831 -131629 38887 -131585
rect 38931 -131629 39387 -131585
rect 39431 -131629 39487 -131585
rect 39531 -131629 39587 -131585
rect 39631 -131629 39687 -131585
rect 39731 -131629 39787 -131585
rect 39831 -131629 39887 -131585
rect 39931 -131629 39987 -131585
rect 40031 -131629 40087 -131585
rect 40131 -131629 40187 -131585
rect 40231 -131629 40287 -131585
rect 40331 -131629 40387 -131585
rect 40431 -131629 40487 -131585
rect 40531 -131629 40587 -131585
rect 40631 -131629 40687 -131585
rect 40731 -131629 40787 -131585
rect 40831 -131629 40887 -131585
rect 40931 -131629 41387 -131585
rect 41431 -131629 41487 -131585
rect 41531 -131629 41587 -131585
rect 41631 -131629 41687 -131585
rect 41731 -131629 41787 -131585
rect 41831 -131629 41887 -131585
rect 41931 -131629 41987 -131585
rect 42031 -131629 42087 -131585
rect 42131 -131629 42187 -131585
rect 42231 -131629 42287 -131585
rect 42331 -131629 42387 -131585
rect 42431 -131629 42487 -131585
rect 42531 -131629 42587 -131585
rect 42631 -131629 42687 -131585
rect 42731 -131629 42787 -131585
rect 42831 -131629 42887 -131585
rect 42931 -131629 43387 -131585
rect 43431 -131629 43487 -131585
rect 43531 -131629 43587 -131585
rect 43631 -131629 43687 -131585
rect 43731 -131629 43787 -131585
rect 43831 -131629 43887 -131585
rect 43931 -131629 43987 -131585
rect 44031 -131629 44087 -131585
rect 44131 -131629 44187 -131585
rect 44231 -131629 44287 -131585
rect 44331 -131629 44387 -131585
rect 44431 -131629 44487 -131585
rect 44531 -131629 44587 -131585
rect 44631 -131629 44687 -131585
rect 44731 -131629 44787 -131585
rect 44831 -131629 44887 -131585
rect 44931 -131629 47953 -131585
rect 34207 -131685 47953 -131629
rect 34207 -131729 37387 -131685
rect 37431 -131729 37487 -131685
rect 37531 -131729 37587 -131685
rect 37631 -131729 37687 -131685
rect 37731 -131729 37787 -131685
rect 37831 -131729 37887 -131685
rect 37931 -131729 37987 -131685
rect 38031 -131729 38087 -131685
rect 38131 -131729 38187 -131685
rect 38231 -131729 38287 -131685
rect 38331 -131729 38387 -131685
rect 38431 -131729 38487 -131685
rect 38531 -131729 38587 -131685
rect 38631 -131729 38687 -131685
rect 38731 -131729 38787 -131685
rect 38831 -131729 38887 -131685
rect 38931 -131729 39387 -131685
rect 39431 -131729 39487 -131685
rect 39531 -131729 39587 -131685
rect 39631 -131729 39687 -131685
rect 39731 -131729 39787 -131685
rect 39831 -131729 39887 -131685
rect 39931 -131729 39987 -131685
rect 40031 -131729 40087 -131685
rect 40131 -131729 40187 -131685
rect 40231 -131729 40287 -131685
rect 40331 -131729 40387 -131685
rect 40431 -131729 40487 -131685
rect 40531 -131729 40587 -131685
rect 40631 -131729 40687 -131685
rect 40731 -131729 40787 -131685
rect 40831 -131729 40887 -131685
rect 40931 -131729 41387 -131685
rect 41431 -131729 41487 -131685
rect 41531 -131729 41587 -131685
rect 41631 -131729 41687 -131685
rect 41731 -131729 41787 -131685
rect 41831 -131729 41887 -131685
rect 41931 -131729 41987 -131685
rect 42031 -131729 42087 -131685
rect 42131 -131729 42187 -131685
rect 42231 -131729 42287 -131685
rect 42331 -131729 42387 -131685
rect 42431 -131729 42487 -131685
rect 42531 -131729 42587 -131685
rect 42631 -131729 42687 -131685
rect 42731 -131729 42787 -131685
rect 42831 -131729 42887 -131685
rect 42931 -131729 43387 -131685
rect 43431 -131729 43487 -131685
rect 43531 -131729 43587 -131685
rect 43631 -131729 43687 -131685
rect 43731 -131729 43787 -131685
rect 43831 -131729 43887 -131685
rect 43931 -131729 43987 -131685
rect 44031 -131729 44087 -131685
rect 44131 -131729 44187 -131685
rect 44231 -131729 44287 -131685
rect 44331 -131729 44387 -131685
rect 44431 -131729 44487 -131685
rect 44531 -131729 44587 -131685
rect 44631 -131729 44687 -131685
rect 44731 -131729 44787 -131685
rect 44831 -131729 44887 -131685
rect 44931 -131729 47953 -131685
rect 34207 -131785 47953 -131729
rect 34207 -131829 37387 -131785
rect 37431 -131829 37487 -131785
rect 37531 -131829 37587 -131785
rect 37631 -131829 37687 -131785
rect 37731 -131829 37787 -131785
rect 37831 -131829 37887 -131785
rect 37931 -131829 37987 -131785
rect 38031 -131829 38087 -131785
rect 38131 -131829 38187 -131785
rect 38231 -131829 38287 -131785
rect 38331 -131829 38387 -131785
rect 38431 -131829 38487 -131785
rect 38531 -131829 38587 -131785
rect 38631 -131829 38687 -131785
rect 38731 -131829 38787 -131785
rect 38831 -131829 38887 -131785
rect 38931 -131829 39387 -131785
rect 39431 -131829 39487 -131785
rect 39531 -131829 39587 -131785
rect 39631 -131829 39687 -131785
rect 39731 -131829 39787 -131785
rect 39831 -131829 39887 -131785
rect 39931 -131829 39987 -131785
rect 40031 -131829 40087 -131785
rect 40131 -131829 40187 -131785
rect 40231 -131829 40287 -131785
rect 40331 -131829 40387 -131785
rect 40431 -131829 40487 -131785
rect 40531 -131829 40587 -131785
rect 40631 -131829 40687 -131785
rect 40731 -131829 40787 -131785
rect 40831 -131829 40887 -131785
rect 40931 -131829 41387 -131785
rect 41431 -131829 41487 -131785
rect 41531 -131829 41587 -131785
rect 41631 -131829 41687 -131785
rect 41731 -131829 41787 -131785
rect 41831 -131829 41887 -131785
rect 41931 -131829 41987 -131785
rect 42031 -131829 42087 -131785
rect 42131 -131829 42187 -131785
rect 42231 -131829 42287 -131785
rect 42331 -131829 42387 -131785
rect 42431 -131829 42487 -131785
rect 42531 -131829 42587 -131785
rect 42631 -131829 42687 -131785
rect 42731 -131829 42787 -131785
rect 42831 -131829 42887 -131785
rect 42931 -131829 43387 -131785
rect 43431 -131829 43487 -131785
rect 43531 -131829 43587 -131785
rect 43631 -131829 43687 -131785
rect 43731 -131829 43787 -131785
rect 43831 -131829 43887 -131785
rect 43931 -131829 43987 -131785
rect 44031 -131829 44087 -131785
rect 44131 -131829 44187 -131785
rect 44231 -131829 44287 -131785
rect 44331 -131829 44387 -131785
rect 44431 -131829 44487 -131785
rect 44531 -131829 44587 -131785
rect 44631 -131829 44687 -131785
rect 44731 -131829 44787 -131785
rect 44831 -131829 44887 -131785
rect 44931 -131829 47953 -131785
rect 34207 -131885 47953 -131829
rect 34207 -131929 37387 -131885
rect 37431 -131929 37487 -131885
rect 37531 -131929 37587 -131885
rect 37631 -131929 37687 -131885
rect 37731 -131929 37787 -131885
rect 37831 -131929 37887 -131885
rect 37931 -131929 37987 -131885
rect 38031 -131929 38087 -131885
rect 38131 -131929 38187 -131885
rect 38231 -131929 38287 -131885
rect 38331 -131929 38387 -131885
rect 38431 -131929 38487 -131885
rect 38531 -131929 38587 -131885
rect 38631 -131929 38687 -131885
rect 38731 -131929 38787 -131885
rect 38831 -131929 38887 -131885
rect 38931 -131929 39387 -131885
rect 39431 -131929 39487 -131885
rect 39531 -131929 39587 -131885
rect 39631 -131929 39687 -131885
rect 39731 -131929 39787 -131885
rect 39831 -131929 39887 -131885
rect 39931 -131929 39987 -131885
rect 40031 -131929 40087 -131885
rect 40131 -131929 40187 -131885
rect 40231 -131929 40287 -131885
rect 40331 -131929 40387 -131885
rect 40431 -131929 40487 -131885
rect 40531 -131929 40587 -131885
rect 40631 -131929 40687 -131885
rect 40731 -131929 40787 -131885
rect 40831 -131929 40887 -131885
rect 40931 -131929 41387 -131885
rect 41431 -131929 41487 -131885
rect 41531 -131929 41587 -131885
rect 41631 -131929 41687 -131885
rect 41731 -131929 41787 -131885
rect 41831 -131929 41887 -131885
rect 41931 -131929 41987 -131885
rect 42031 -131929 42087 -131885
rect 42131 -131929 42187 -131885
rect 42231 -131929 42287 -131885
rect 42331 -131929 42387 -131885
rect 42431 -131929 42487 -131885
rect 42531 -131929 42587 -131885
rect 42631 -131929 42687 -131885
rect 42731 -131929 42787 -131885
rect 42831 -131929 42887 -131885
rect 42931 -131929 43387 -131885
rect 43431 -131929 43487 -131885
rect 43531 -131929 43587 -131885
rect 43631 -131929 43687 -131885
rect 43731 -131929 43787 -131885
rect 43831 -131929 43887 -131885
rect 43931 -131929 43987 -131885
rect 44031 -131929 44087 -131885
rect 44131 -131929 44187 -131885
rect 44231 -131929 44287 -131885
rect 44331 -131929 44387 -131885
rect 44431 -131929 44487 -131885
rect 44531 -131929 44587 -131885
rect 44631 -131929 44687 -131885
rect 44731 -131929 44787 -131885
rect 44831 -131929 44887 -131885
rect 44931 -131929 47953 -131885
rect 34207 -131985 47953 -131929
rect 34207 -132029 37387 -131985
rect 37431 -132029 37487 -131985
rect 37531 -132029 37587 -131985
rect 37631 -132029 37687 -131985
rect 37731 -132029 37787 -131985
rect 37831 -132029 37887 -131985
rect 37931 -132029 37987 -131985
rect 38031 -132029 38087 -131985
rect 38131 -132029 38187 -131985
rect 38231 -132029 38287 -131985
rect 38331 -132029 38387 -131985
rect 38431 -132029 38487 -131985
rect 38531 -132029 38587 -131985
rect 38631 -132029 38687 -131985
rect 38731 -132029 38787 -131985
rect 38831 -132029 38887 -131985
rect 38931 -132029 39387 -131985
rect 39431 -132029 39487 -131985
rect 39531 -132029 39587 -131985
rect 39631 -132029 39687 -131985
rect 39731 -132029 39787 -131985
rect 39831 -132029 39887 -131985
rect 39931 -132029 39987 -131985
rect 40031 -132029 40087 -131985
rect 40131 -132029 40187 -131985
rect 40231 -132029 40287 -131985
rect 40331 -132029 40387 -131985
rect 40431 -132029 40487 -131985
rect 40531 -132029 40587 -131985
rect 40631 -132029 40687 -131985
rect 40731 -132029 40787 -131985
rect 40831 -132029 40887 -131985
rect 40931 -132029 41387 -131985
rect 41431 -132029 41487 -131985
rect 41531 -132029 41587 -131985
rect 41631 -132029 41687 -131985
rect 41731 -132029 41787 -131985
rect 41831 -132029 41887 -131985
rect 41931 -132029 41987 -131985
rect 42031 -132029 42087 -131985
rect 42131 -132029 42187 -131985
rect 42231 -132029 42287 -131985
rect 42331 -132029 42387 -131985
rect 42431 -132029 42487 -131985
rect 42531 -132029 42587 -131985
rect 42631 -132029 42687 -131985
rect 42731 -132029 42787 -131985
rect 42831 -132029 42887 -131985
rect 42931 -132029 43387 -131985
rect 43431 -132029 43487 -131985
rect 43531 -132029 43587 -131985
rect 43631 -132029 43687 -131985
rect 43731 -132029 43787 -131985
rect 43831 -132029 43887 -131985
rect 43931 -132029 43987 -131985
rect 44031 -132029 44087 -131985
rect 44131 -132029 44187 -131985
rect 44231 -132029 44287 -131985
rect 44331 -132029 44387 -131985
rect 44431 -132029 44487 -131985
rect 44531 -132029 44587 -131985
rect 44631 -132029 44687 -131985
rect 44731 -132029 44787 -131985
rect 44831 -132029 44887 -131985
rect 44931 -132029 47953 -131985
rect 34207 -132085 47953 -132029
rect 34207 -132129 37387 -132085
rect 37431 -132129 37487 -132085
rect 37531 -132129 37587 -132085
rect 37631 -132129 37687 -132085
rect 37731 -132129 37787 -132085
rect 37831 -132129 37887 -132085
rect 37931 -132129 37987 -132085
rect 38031 -132129 38087 -132085
rect 38131 -132129 38187 -132085
rect 38231 -132129 38287 -132085
rect 38331 -132129 38387 -132085
rect 38431 -132129 38487 -132085
rect 38531 -132129 38587 -132085
rect 38631 -132129 38687 -132085
rect 38731 -132129 38787 -132085
rect 38831 -132129 38887 -132085
rect 38931 -132129 39387 -132085
rect 39431 -132129 39487 -132085
rect 39531 -132129 39587 -132085
rect 39631 -132129 39687 -132085
rect 39731 -132129 39787 -132085
rect 39831 -132129 39887 -132085
rect 39931 -132129 39987 -132085
rect 40031 -132129 40087 -132085
rect 40131 -132129 40187 -132085
rect 40231 -132129 40287 -132085
rect 40331 -132129 40387 -132085
rect 40431 -132129 40487 -132085
rect 40531 -132129 40587 -132085
rect 40631 -132129 40687 -132085
rect 40731 -132129 40787 -132085
rect 40831 -132129 40887 -132085
rect 40931 -132129 41387 -132085
rect 41431 -132129 41487 -132085
rect 41531 -132129 41587 -132085
rect 41631 -132129 41687 -132085
rect 41731 -132129 41787 -132085
rect 41831 -132129 41887 -132085
rect 41931 -132129 41987 -132085
rect 42031 -132129 42087 -132085
rect 42131 -132129 42187 -132085
rect 42231 -132129 42287 -132085
rect 42331 -132129 42387 -132085
rect 42431 -132129 42487 -132085
rect 42531 -132129 42587 -132085
rect 42631 -132129 42687 -132085
rect 42731 -132129 42787 -132085
rect 42831 -132129 42887 -132085
rect 42931 -132129 43387 -132085
rect 43431 -132129 43487 -132085
rect 43531 -132129 43587 -132085
rect 43631 -132129 43687 -132085
rect 43731 -132129 43787 -132085
rect 43831 -132129 43887 -132085
rect 43931 -132129 43987 -132085
rect 44031 -132129 44087 -132085
rect 44131 -132129 44187 -132085
rect 44231 -132129 44287 -132085
rect 44331 -132129 44387 -132085
rect 44431 -132129 44487 -132085
rect 44531 -132129 44587 -132085
rect 44631 -132129 44687 -132085
rect 44731 -132129 44787 -132085
rect 44831 -132129 44887 -132085
rect 44931 -132129 47953 -132085
rect 34207 -132185 47953 -132129
rect 34207 -132229 37387 -132185
rect 37431 -132229 37487 -132185
rect 37531 -132229 37587 -132185
rect 37631 -132229 37687 -132185
rect 37731 -132229 37787 -132185
rect 37831 -132229 37887 -132185
rect 37931 -132229 37987 -132185
rect 38031 -132229 38087 -132185
rect 38131 -132229 38187 -132185
rect 38231 -132229 38287 -132185
rect 38331 -132229 38387 -132185
rect 38431 -132229 38487 -132185
rect 38531 -132229 38587 -132185
rect 38631 -132229 38687 -132185
rect 38731 -132229 38787 -132185
rect 38831 -132229 38887 -132185
rect 38931 -132229 39387 -132185
rect 39431 -132229 39487 -132185
rect 39531 -132229 39587 -132185
rect 39631 -132229 39687 -132185
rect 39731 -132229 39787 -132185
rect 39831 -132229 39887 -132185
rect 39931 -132229 39987 -132185
rect 40031 -132229 40087 -132185
rect 40131 -132229 40187 -132185
rect 40231 -132229 40287 -132185
rect 40331 -132229 40387 -132185
rect 40431 -132229 40487 -132185
rect 40531 -132229 40587 -132185
rect 40631 -132229 40687 -132185
rect 40731 -132229 40787 -132185
rect 40831 -132229 40887 -132185
rect 40931 -132229 41387 -132185
rect 41431 -132229 41487 -132185
rect 41531 -132229 41587 -132185
rect 41631 -132229 41687 -132185
rect 41731 -132229 41787 -132185
rect 41831 -132229 41887 -132185
rect 41931 -132229 41987 -132185
rect 42031 -132229 42087 -132185
rect 42131 -132229 42187 -132185
rect 42231 -132229 42287 -132185
rect 42331 -132229 42387 -132185
rect 42431 -132229 42487 -132185
rect 42531 -132229 42587 -132185
rect 42631 -132229 42687 -132185
rect 42731 -132229 42787 -132185
rect 42831 -132229 42887 -132185
rect 42931 -132229 43387 -132185
rect 43431 -132229 43487 -132185
rect 43531 -132229 43587 -132185
rect 43631 -132229 43687 -132185
rect 43731 -132229 43787 -132185
rect 43831 -132229 43887 -132185
rect 43931 -132229 43987 -132185
rect 44031 -132229 44087 -132185
rect 44131 -132229 44187 -132185
rect 44231 -132229 44287 -132185
rect 44331 -132229 44387 -132185
rect 44431 -132229 44487 -132185
rect 44531 -132229 44587 -132185
rect 44631 -132229 44687 -132185
rect 44731 -132229 44787 -132185
rect 44831 -132229 44887 -132185
rect 44931 -132229 47953 -132185
rect 34207 -132285 47953 -132229
rect 34207 -132329 37387 -132285
rect 37431 -132329 37487 -132285
rect 37531 -132329 37587 -132285
rect 37631 -132329 37687 -132285
rect 37731 -132329 37787 -132285
rect 37831 -132329 37887 -132285
rect 37931 -132329 37987 -132285
rect 38031 -132329 38087 -132285
rect 38131 -132329 38187 -132285
rect 38231 -132329 38287 -132285
rect 38331 -132329 38387 -132285
rect 38431 -132329 38487 -132285
rect 38531 -132329 38587 -132285
rect 38631 -132329 38687 -132285
rect 38731 -132329 38787 -132285
rect 38831 -132329 38887 -132285
rect 38931 -132329 39387 -132285
rect 39431 -132329 39487 -132285
rect 39531 -132329 39587 -132285
rect 39631 -132329 39687 -132285
rect 39731 -132329 39787 -132285
rect 39831 -132329 39887 -132285
rect 39931 -132329 39987 -132285
rect 40031 -132329 40087 -132285
rect 40131 -132329 40187 -132285
rect 40231 -132329 40287 -132285
rect 40331 -132329 40387 -132285
rect 40431 -132329 40487 -132285
rect 40531 -132329 40587 -132285
rect 40631 -132329 40687 -132285
rect 40731 -132329 40787 -132285
rect 40831 -132329 40887 -132285
rect 40931 -132329 41387 -132285
rect 41431 -132329 41487 -132285
rect 41531 -132329 41587 -132285
rect 41631 -132329 41687 -132285
rect 41731 -132329 41787 -132285
rect 41831 -132329 41887 -132285
rect 41931 -132329 41987 -132285
rect 42031 -132329 42087 -132285
rect 42131 -132329 42187 -132285
rect 42231 -132329 42287 -132285
rect 42331 -132329 42387 -132285
rect 42431 -132329 42487 -132285
rect 42531 -132329 42587 -132285
rect 42631 -132329 42687 -132285
rect 42731 -132329 42787 -132285
rect 42831 -132329 42887 -132285
rect 42931 -132329 43387 -132285
rect 43431 -132329 43487 -132285
rect 43531 -132329 43587 -132285
rect 43631 -132329 43687 -132285
rect 43731 -132329 43787 -132285
rect 43831 -132329 43887 -132285
rect 43931 -132329 43987 -132285
rect 44031 -132329 44087 -132285
rect 44131 -132329 44187 -132285
rect 44231 -132329 44287 -132285
rect 44331 -132329 44387 -132285
rect 44431 -132329 44487 -132285
rect 44531 -132329 44587 -132285
rect 44631 -132329 44687 -132285
rect 44731 -132329 44787 -132285
rect 44831 -132329 44887 -132285
rect 44931 -132329 47953 -132285
rect 34207 -132385 47953 -132329
rect 34207 -132429 37387 -132385
rect 37431 -132429 37487 -132385
rect 37531 -132429 37587 -132385
rect 37631 -132429 37687 -132385
rect 37731 -132429 37787 -132385
rect 37831 -132429 37887 -132385
rect 37931 -132429 37987 -132385
rect 38031 -132429 38087 -132385
rect 38131 -132429 38187 -132385
rect 38231 -132429 38287 -132385
rect 38331 -132429 38387 -132385
rect 38431 -132429 38487 -132385
rect 38531 -132429 38587 -132385
rect 38631 -132429 38687 -132385
rect 38731 -132429 38787 -132385
rect 38831 -132429 38887 -132385
rect 38931 -132429 39387 -132385
rect 39431 -132429 39487 -132385
rect 39531 -132429 39587 -132385
rect 39631 -132429 39687 -132385
rect 39731 -132429 39787 -132385
rect 39831 -132429 39887 -132385
rect 39931 -132429 39987 -132385
rect 40031 -132429 40087 -132385
rect 40131 -132429 40187 -132385
rect 40231 -132429 40287 -132385
rect 40331 -132429 40387 -132385
rect 40431 -132429 40487 -132385
rect 40531 -132429 40587 -132385
rect 40631 -132429 40687 -132385
rect 40731 -132429 40787 -132385
rect 40831 -132429 40887 -132385
rect 40931 -132429 41387 -132385
rect 41431 -132429 41487 -132385
rect 41531 -132429 41587 -132385
rect 41631 -132429 41687 -132385
rect 41731 -132429 41787 -132385
rect 41831 -132429 41887 -132385
rect 41931 -132429 41987 -132385
rect 42031 -132429 42087 -132385
rect 42131 -132429 42187 -132385
rect 42231 -132429 42287 -132385
rect 42331 -132429 42387 -132385
rect 42431 -132429 42487 -132385
rect 42531 -132429 42587 -132385
rect 42631 -132429 42687 -132385
rect 42731 -132429 42787 -132385
rect 42831 -132429 42887 -132385
rect 42931 -132429 43387 -132385
rect 43431 -132429 43487 -132385
rect 43531 -132429 43587 -132385
rect 43631 -132429 43687 -132385
rect 43731 -132429 43787 -132385
rect 43831 -132429 43887 -132385
rect 43931 -132429 43987 -132385
rect 44031 -132429 44087 -132385
rect 44131 -132429 44187 -132385
rect 44231 -132429 44287 -132385
rect 44331 -132429 44387 -132385
rect 44431 -132429 44487 -132385
rect 44531 -132429 44587 -132385
rect 44631 -132429 44687 -132385
rect 44731 -132429 44787 -132385
rect 44831 -132429 44887 -132385
rect 44931 -132429 47953 -132385
rect 34207 -132485 47953 -132429
rect 34207 -132529 37387 -132485
rect 37431 -132529 37487 -132485
rect 37531 -132529 37587 -132485
rect 37631 -132529 37687 -132485
rect 37731 -132529 37787 -132485
rect 37831 -132529 37887 -132485
rect 37931 -132529 37987 -132485
rect 38031 -132529 38087 -132485
rect 38131 -132529 38187 -132485
rect 38231 -132529 38287 -132485
rect 38331 -132529 38387 -132485
rect 38431 -132529 38487 -132485
rect 38531 -132529 38587 -132485
rect 38631 -132529 38687 -132485
rect 38731 -132529 38787 -132485
rect 38831 -132529 38887 -132485
rect 38931 -132529 39387 -132485
rect 39431 -132529 39487 -132485
rect 39531 -132529 39587 -132485
rect 39631 -132529 39687 -132485
rect 39731 -132529 39787 -132485
rect 39831 -132529 39887 -132485
rect 39931 -132529 39987 -132485
rect 40031 -132529 40087 -132485
rect 40131 -132529 40187 -132485
rect 40231 -132529 40287 -132485
rect 40331 -132529 40387 -132485
rect 40431 -132529 40487 -132485
rect 40531 -132529 40587 -132485
rect 40631 -132529 40687 -132485
rect 40731 -132529 40787 -132485
rect 40831 -132529 40887 -132485
rect 40931 -132529 41387 -132485
rect 41431 -132529 41487 -132485
rect 41531 -132529 41587 -132485
rect 41631 -132529 41687 -132485
rect 41731 -132529 41787 -132485
rect 41831 -132529 41887 -132485
rect 41931 -132529 41987 -132485
rect 42031 -132529 42087 -132485
rect 42131 -132529 42187 -132485
rect 42231 -132529 42287 -132485
rect 42331 -132529 42387 -132485
rect 42431 -132529 42487 -132485
rect 42531 -132529 42587 -132485
rect 42631 -132529 42687 -132485
rect 42731 -132529 42787 -132485
rect 42831 -132529 42887 -132485
rect 42931 -132529 43387 -132485
rect 43431 -132529 43487 -132485
rect 43531 -132529 43587 -132485
rect 43631 -132529 43687 -132485
rect 43731 -132529 43787 -132485
rect 43831 -132529 43887 -132485
rect 43931 -132529 43987 -132485
rect 44031 -132529 44087 -132485
rect 44131 -132529 44187 -132485
rect 44231 -132529 44287 -132485
rect 44331 -132529 44387 -132485
rect 44431 -132529 44487 -132485
rect 44531 -132529 44587 -132485
rect 44631 -132529 44687 -132485
rect 44731 -132529 44787 -132485
rect 44831 -132529 44887 -132485
rect 44931 -132529 47953 -132485
rect 34207 -132585 47953 -132529
rect 34207 -132629 37387 -132585
rect 37431 -132629 37487 -132585
rect 37531 -132629 37587 -132585
rect 37631 -132629 37687 -132585
rect 37731 -132629 37787 -132585
rect 37831 -132629 37887 -132585
rect 37931 -132629 37987 -132585
rect 38031 -132629 38087 -132585
rect 38131 -132629 38187 -132585
rect 38231 -132629 38287 -132585
rect 38331 -132629 38387 -132585
rect 38431 -132629 38487 -132585
rect 38531 -132629 38587 -132585
rect 38631 -132629 38687 -132585
rect 38731 -132629 38787 -132585
rect 38831 -132629 38887 -132585
rect 38931 -132629 39387 -132585
rect 39431 -132629 39487 -132585
rect 39531 -132629 39587 -132585
rect 39631 -132629 39687 -132585
rect 39731 -132629 39787 -132585
rect 39831 -132629 39887 -132585
rect 39931 -132629 39987 -132585
rect 40031 -132629 40087 -132585
rect 40131 -132629 40187 -132585
rect 40231 -132629 40287 -132585
rect 40331 -132629 40387 -132585
rect 40431 -132629 40487 -132585
rect 40531 -132629 40587 -132585
rect 40631 -132629 40687 -132585
rect 40731 -132629 40787 -132585
rect 40831 -132629 40887 -132585
rect 40931 -132629 41387 -132585
rect 41431 -132629 41487 -132585
rect 41531 -132629 41587 -132585
rect 41631 -132629 41687 -132585
rect 41731 -132629 41787 -132585
rect 41831 -132629 41887 -132585
rect 41931 -132629 41987 -132585
rect 42031 -132629 42087 -132585
rect 42131 -132629 42187 -132585
rect 42231 -132629 42287 -132585
rect 42331 -132629 42387 -132585
rect 42431 -132629 42487 -132585
rect 42531 -132629 42587 -132585
rect 42631 -132629 42687 -132585
rect 42731 -132629 42787 -132585
rect 42831 -132629 42887 -132585
rect 42931 -132629 43387 -132585
rect 43431 -132629 43487 -132585
rect 43531 -132629 43587 -132585
rect 43631 -132629 43687 -132585
rect 43731 -132629 43787 -132585
rect 43831 -132629 43887 -132585
rect 43931 -132629 43987 -132585
rect 44031 -132629 44087 -132585
rect 44131 -132629 44187 -132585
rect 44231 -132629 44287 -132585
rect 44331 -132629 44387 -132585
rect 44431 -132629 44487 -132585
rect 44531 -132629 44587 -132585
rect 44631 -132629 44687 -132585
rect 44731 -132629 44787 -132585
rect 44831 -132629 44887 -132585
rect 44931 -132629 47953 -132585
rect 34207 -132685 47953 -132629
rect 34207 -132729 37387 -132685
rect 37431 -132729 37487 -132685
rect 37531 -132729 37587 -132685
rect 37631 -132729 37687 -132685
rect 37731 -132729 37787 -132685
rect 37831 -132729 37887 -132685
rect 37931 -132729 37987 -132685
rect 38031 -132729 38087 -132685
rect 38131 -132729 38187 -132685
rect 38231 -132729 38287 -132685
rect 38331 -132729 38387 -132685
rect 38431 -132729 38487 -132685
rect 38531 -132729 38587 -132685
rect 38631 -132729 38687 -132685
rect 38731 -132729 38787 -132685
rect 38831 -132729 38887 -132685
rect 38931 -132729 39387 -132685
rect 39431 -132729 39487 -132685
rect 39531 -132729 39587 -132685
rect 39631 -132729 39687 -132685
rect 39731 -132729 39787 -132685
rect 39831 -132729 39887 -132685
rect 39931 -132729 39987 -132685
rect 40031 -132729 40087 -132685
rect 40131 -132729 40187 -132685
rect 40231 -132729 40287 -132685
rect 40331 -132729 40387 -132685
rect 40431 -132729 40487 -132685
rect 40531 -132729 40587 -132685
rect 40631 -132729 40687 -132685
rect 40731 -132729 40787 -132685
rect 40831 -132729 40887 -132685
rect 40931 -132729 41387 -132685
rect 41431 -132729 41487 -132685
rect 41531 -132729 41587 -132685
rect 41631 -132729 41687 -132685
rect 41731 -132729 41787 -132685
rect 41831 -132729 41887 -132685
rect 41931 -132729 41987 -132685
rect 42031 -132729 42087 -132685
rect 42131 -132729 42187 -132685
rect 42231 -132729 42287 -132685
rect 42331 -132729 42387 -132685
rect 42431 -132729 42487 -132685
rect 42531 -132729 42587 -132685
rect 42631 -132729 42687 -132685
rect 42731 -132729 42787 -132685
rect 42831 -132729 42887 -132685
rect 42931 -132729 43387 -132685
rect 43431 -132729 43487 -132685
rect 43531 -132729 43587 -132685
rect 43631 -132729 43687 -132685
rect 43731 -132729 43787 -132685
rect 43831 -132729 43887 -132685
rect 43931 -132729 43987 -132685
rect 44031 -132729 44087 -132685
rect 44131 -132729 44187 -132685
rect 44231 -132729 44287 -132685
rect 44331 -132729 44387 -132685
rect 44431 -132729 44487 -132685
rect 44531 -132729 44587 -132685
rect 44631 -132729 44687 -132685
rect 44731 -132729 44787 -132685
rect 44831 -132729 44887 -132685
rect 44931 -132729 47953 -132685
rect 34207 -132785 47953 -132729
rect 34207 -132829 37387 -132785
rect 37431 -132829 37487 -132785
rect 37531 -132829 37587 -132785
rect 37631 -132829 37687 -132785
rect 37731 -132829 37787 -132785
rect 37831 -132829 37887 -132785
rect 37931 -132829 37987 -132785
rect 38031 -132829 38087 -132785
rect 38131 -132829 38187 -132785
rect 38231 -132829 38287 -132785
rect 38331 -132829 38387 -132785
rect 38431 -132829 38487 -132785
rect 38531 -132829 38587 -132785
rect 38631 -132829 38687 -132785
rect 38731 -132829 38787 -132785
rect 38831 -132829 38887 -132785
rect 38931 -132829 39387 -132785
rect 39431 -132829 39487 -132785
rect 39531 -132829 39587 -132785
rect 39631 -132829 39687 -132785
rect 39731 -132829 39787 -132785
rect 39831 -132829 39887 -132785
rect 39931 -132829 39987 -132785
rect 40031 -132829 40087 -132785
rect 40131 -132829 40187 -132785
rect 40231 -132829 40287 -132785
rect 40331 -132829 40387 -132785
rect 40431 -132829 40487 -132785
rect 40531 -132829 40587 -132785
rect 40631 -132829 40687 -132785
rect 40731 -132829 40787 -132785
rect 40831 -132829 40887 -132785
rect 40931 -132829 41387 -132785
rect 41431 -132829 41487 -132785
rect 41531 -132829 41587 -132785
rect 41631 -132829 41687 -132785
rect 41731 -132829 41787 -132785
rect 41831 -132829 41887 -132785
rect 41931 -132829 41987 -132785
rect 42031 -132829 42087 -132785
rect 42131 -132829 42187 -132785
rect 42231 -132829 42287 -132785
rect 42331 -132829 42387 -132785
rect 42431 -132829 42487 -132785
rect 42531 -132829 42587 -132785
rect 42631 -132829 42687 -132785
rect 42731 -132829 42787 -132785
rect 42831 -132829 42887 -132785
rect 42931 -132829 43387 -132785
rect 43431 -132829 43487 -132785
rect 43531 -132829 43587 -132785
rect 43631 -132829 43687 -132785
rect 43731 -132829 43787 -132785
rect 43831 -132829 43887 -132785
rect 43931 -132829 43987 -132785
rect 44031 -132829 44087 -132785
rect 44131 -132829 44187 -132785
rect 44231 -132829 44287 -132785
rect 44331 -132829 44387 -132785
rect 44431 -132829 44487 -132785
rect 44531 -132829 44587 -132785
rect 44631 -132829 44687 -132785
rect 44731 -132829 44787 -132785
rect 44831 -132829 44887 -132785
rect 44931 -132829 47953 -132785
rect 34207 -132885 47953 -132829
rect 34207 -132929 37387 -132885
rect 37431 -132929 37487 -132885
rect 37531 -132929 37587 -132885
rect 37631 -132929 37687 -132885
rect 37731 -132929 37787 -132885
rect 37831 -132929 37887 -132885
rect 37931 -132929 37987 -132885
rect 38031 -132929 38087 -132885
rect 38131 -132929 38187 -132885
rect 38231 -132929 38287 -132885
rect 38331 -132929 38387 -132885
rect 38431 -132929 38487 -132885
rect 38531 -132929 38587 -132885
rect 38631 -132929 38687 -132885
rect 38731 -132929 38787 -132885
rect 38831 -132929 38887 -132885
rect 38931 -132929 39387 -132885
rect 39431 -132929 39487 -132885
rect 39531 -132929 39587 -132885
rect 39631 -132929 39687 -132885
rect 39731 -132929 39787 -132885
rect 39831 -132929 39887 -132885
rect 39931 -132929 39987 -132885
rect 40031 -132929 40087 -132885
rect 40131 -132929 40187 -132885
rect 40231 -132929 40287 -132885
rect 40331 -132929 40387 -132885
rect 40431 -132929 40487 -132885
rect 40531 -132929 40587 -132885
rect 40631 -132929 40687 -132885
rect 40731 -132929 40787 -132885
rect 40831 -132929 40887 -132885
rect 40931 -132929 41387 -132885
rect 41431 -132929 41487 -132885
rect 41531 -132929 41587 -132885
rect 41631 -132929 41687 -132885
rect 41731 -132929 41787 -132885
rect 41831 -132929 41887 -132885
rect 41931 -132929 41987 -132885
rect 42031 -132929 42087 -132885
rect 42131 -132929 42187 -132885
rect 42231 -132929 42287 -132885
rect 42331 -132929 42387 -132885
rect 42431 -132929 42487 -132885
rect 42531 -132929 42587 -132885
rect 42631 -132929 42687 -132885
rect 42731 -132929 42787 -132885
rect 42831 -132929 42887 -132885
rect 42931 -132929 43387 -132885
rect 43431 -132929 43487 -132885
rect 43531 -132929 43587 -132885
rect 43631 -132929 43687 -132885
rect 43731 -132929 43787 -132885
rect 43831 -132929 43887 -132885
rect 43931 -132929 43987 -132885
rect 44031 -132929 44087 -132885
rect 44131 -132929 44187 -132885
rect 44231 -132929 44287 -132885
rect 44331 -132929 44387 -132885
rect 44431 -132929 44487 -132885
rect 44531 -132929 44587 -132885
rect 44631 -132929 44687 -132885
rect 44731 -132929 44787 -132885
rect 44831 -132929 44887 -132885
rect 44931 -132929 47953 -132885
rect 34207 -133867 47953 -132929
rect -87194 -140275 -83265 -140231
rect -83221 -140275 -83165 -140231
rect -83121 -140275 -83065 -140231
rect -83021 -140275 -82965 -140231
rect -82921 -140275 -82865 -140231
rect -82821 -140275 -82765 -140231
rect -82721 -140275 -82665 -140231
rect -82621 -140275 -82565 -140231
rect -82521 -140275 -82465 -140231
rect -82421 -140275 -82365 -140231
rect -82321 -140275 -82265 -140231
rect -82221 -140275 -82165 -140231
rect -82121 -140275 -82065 -140231
rect -82021 -140275 -81965 -140231
rect -81921 -140275 -81865 -140231
rect -81821 -140275 -81765 -140231
rect -81721 -140275 -81265 -140231
rect -81221 -140275 -81165 -140231
rect -81121 -140275 -81065 -140231
rect -81021 -140275 -80965 -140231
rect -80921 -140275 -80865 -140231
rect -80821 -140275 -80765 -140231
rect -80721 -140275 -80665 -140231
rect -80621 -140275 -80565 -140231
rect -80521 -140275 -80465 -140231
rect -80421 -140275 -80365 -140231
rect -80321 -140275 -80265 -140231
rect -80221 -140275 -80165 -140231
rect -80121 -140275 -80065 -140231
rect -80021 -140275 -79965 -140231
rect -79921 -140275 -79865 -140231
rect -79821 -140275 -79765 -140231
rect -79721 -140275 -79265 -140231
rect -79221 -140275 -79165 -140231
rect -79121 -140275 -79065 -140231
rect -79021 -140275 -78965 -140231
rect -78921 -140275 -78865 -140231
rect -78821 -140275 -78765 -140231
rect -78721 -140275 -78665 -140231
rect -78621 -140275 -78565 -140231
rect -78521 -140275 -78465 -140231
rect -78421 -140275 -78365 -140231
rect -78321 -140275 -78265 -140231
rect -78221 -140275 -78165 -140231
rect -78121 -140275 -78065 -140231
rect -78021 -140275 -77965 -140231
rect -77921 -140275 -77865 -140231
rect -77821 -140275 -77765 -140231
rect -77721 -140275 -77265 -140231
rect -77221 -140275 -77165 -140231
rect -77121 -140275 -77065 -140231
rect -77021 -140275 -76965 -140231
rect -76921 -140275 -76865 -140231
rect -76821 -140275 -76765 -140231
rect -76721 -140275 -76665 -140231
rect -76621 -140275 -76565 -140231
rect -76521 -140275 -76465 -140231
rect -76421 -140275 -76365 -140231
rect -76321 -140275 -76265 -140231
rect -76221 -140275 -76165 -140231
rect -76121 -140275 -76065 -140231
rect -76021 -140275 -75965 -140231
rect -75921 -140275 -75865 -140231
rect -75821 -140275 -75765 -140231
rect -75721 -140275 -71799 -140231
rect -87194 -140331 -71799 -140275
rect -87194 -140375 -83265 -140331
rect -83221 -140375 -83165 -140331
rect -83121 -140375 -83065 -140331
rect -83021 -140375 -82965 -140331
rect -82921 -140375 -82865 -140331
rect -82821 -140375 -82765 -140331
rect -82721 -140375 -82665 -140331
rect -82621 -140375 -82565 -140331
rect -82521 -140375 -82465 -140331
rect -82421 -140375 -82365 -140331
rect -82321 -140375 -82265 -140331
rect -82221 -140375 -82165 -140331
rect -82121 -140375 -82065 -140331
rect -82021 -140375 -81965 -140331
rect -81921 -140375 -81865 -140331
rect -81821 -140375 -81765 -140331
rect -81721 -140375 -81265 -140331
rect -81221 -140375 -81165 -140331
rect -81121 -140375 -81065 -140331
rect -81021 -140375 -80965 -140331
rect -80921 -140375 -80865 -140331
rect -80821 -140375 -80765 -140331
rect -80721 -140375 -80665 -140331
rect -80621 -140375 -80565 -140331
rect -80521 -140375 -80465 -140331
rect -80421 -140375 -80365 -140331
rect -80321 -140375 -80265 -140331
rect -80221 -140375 -80165 -140331
rect -80121 -140375 -80065 -140331
rect -80021 -140375 -79965 -140331
rect -79921 -140375 -79865 -140331
rect -79821 -140375 -79765 -140331
rect -79721 -140375 -79265 -140331
rect -79221 -140375 -79165 -140331
rect -79121 -140375 -79065 -140331
rect -79021 -140375 -78965 -140331
rect -78921 -140375 -78865 -140331
rect -78821 -140375 -78765 -140331
rect -78721 -140375 -78665 -140331
rect -78621 -140375 -78565 -140331
rect -78521 -140375 -78465 -140331
rect -78421 -140375 -78365 -140331
rect -78321 -140375 -78265 -140331
rect -78221 -140375 -78165 -140331
rect -78121 -140375 -78065 -140331
rect -78021 -140375 -77965 -140331
rect -77921 -140375 -77865 -140331
rect -77821 -140375 -77765 -140331
rect -77721 -140375 -77265 -140331
rect -77221 -140375 -77165 -140331
rect -77121 -140375 -77065 -140331
rect -77021 -140375 -76965 -140331
rect -76921 -140375 -76865 -140331
rect -76821 -140375 -76765 -140331
rect -76721 -140375 -76665 -140331
rect -76621 -140375 -76565 -140331
rect -76521 -140375 -76465 -140331
rect -76421 -140375 -76365 -140331
rect -76321 -140375 -76265 -140331
rect -76221 -140375 -76165 -140331
rect -76121 -140375 -76065 -140331
rect -76021 -140375 -75965 -140331
rect -75921 -140375 -75865 -140331
rect -75821 -140375 -75765 -140331
rect -75721 -140375 -71799 -140331
rect -87194 -140431 -71799 -140375
rect -87194 -140475 -83265 -140431
rect -83221 -140475 -83165 -140431
rect -83121 -140475 -83065 -140431
rect -83021 -140475 -82965 -140431
rect -82921 -140475 -82865 -140431
rect -82821 -140475 -82765 -140431
rect -82721 -140475 -82665 -140431
rect -82621 -140475 -82565 -140431
rect -82521 -140475 -82465 -140431
rect -82421 -140475 -82365 -140431
rect -82321 -140475 -82265 -140431
rect -82221 -140475 -82165 -140431
rect -82121 -140475 -82065 -140431
rect -82021 -140475 -81965 -140431
rect -81921 -140475 -81865 -140431
rect -81821 -140475 -81765 -140431
rect -81721 -140475 -81265 -140431
rect -81221 -140475 -81165 -140431
rect -81121 -140475 -81065 -140431
rect -81021 -140475 -80965 -140431
rect -80921 -140475 -80865 -140431
rect -80821 -140475 -80765 -140431
rect -80721 -140475 -80665 -140431
rect -80621 -140475 -80565 -140431
rect -80521 -140475 -80465 -140431
rect -80421 -140475 -80365 -140431
rect -80321 -140475 -80265 -140431
rect -80221 -140475 -80165 -140431
rect -80121 -140475 -80065 -140431
rect -80021 -140475 -79965 -140431
rect -79921 -140475 -79865 -140431
rect -79821 -140475 -79765 -140431
rect -79721 -140475 -79265 -140431
rect -79221 -140475 -79165 -140431
rect -79121 -140475 -79065 -140431
rect -79021 -140475 -78965 -140431
rect -78921 -140475 -78865 -140431
rect -78821 -140475 -78765 -140431
rect -78721 -140475 -78665 -140431
rect -78621 -140475 -78565 -140431
rect -78521 -140475 -78465 -140431
rect -78421 -140475 -78365 -140431
rect -78321 -140475 -78265 -140431
rect -78221 -140475 -78165 -140431
rect -78121 -140475 -78065 -140431
rect -78021 -140475 -77965 -140431
rect -77921 -140475 -77865 -140431
rect -77821 -140475 -77765 -140431
rect -77721 -140475 -77265 -140431
rect -77221 -140475 -77165 -140431
rect -77121 -140475 -77065 -140431
rect -77021 -140475 -76965 -140431
rect -76921 -140475 -76865 -140431
rect -76821 -140475 -76765 -140431
rect -76721 -140475 -76665 -140431
rect -76621 -140475 -76565 -140431
rect -76521 -140475 -76465 -140431
rect -76421 -140475 -76365 -140431
rect -76321 -140475 -76265 -140431
rect -76221 -140475 -76165 -140431
rect -76121 -140475 -76065 -140431
rect -76021 -140475 -75965 -140431
rect -75921 -140475 -75865 -140431
rect -75821 -140475 -75765 -140431
rect -75721 -140475 -71799 -140431
rect -87194 -140531 -71799 -140475
rect -87194 -140575 -83265 -140531
rect -83221 -140575 -83165 -140531
rect -83121 -140575 -83065 -140531
rect -83021 -140575 -82965 -140531
rect -82921 -140575 -82865 -140531
rect -82821 -140575 -82765 -140531
rect -82721 -140575 -82665 -140531
rect -82621 -140575 -82565 -140531
rect -82521 -140575 -82465 -140531
rect -82421 -140575 -82365 -140531
rect -82321 -140575 -82265 -140531
rect -82221 -140575 -82165 -140531
rect -82121 -140575 -82065 -140531
rect -82021 -140575 -81965 -140531
rect -81921 -140575 -81865 -140531
rect -81821 -140575 -81765 -140531
rect -81721 -140575 -81265 -140531
rect -81221 -140575 -81165 -140531
rect -81121 -140575 -81065 -140531
rect -81021 -140575 -80965 -140531
rect -80921 -140575 -80865 -140531
rect -80821 -140575 -80765 -140531
rect -80721 -140575 -80665 -140531
rect -80621 -140575 -80565 -140531
rect -80521 -140575 -80465 -140531
rect -80421 -140575 -80365 -140531
rect -80321 -140575 -80265 -140531
rect -80221 -140575 -80165 -140531
rect -80121 -140575 -80065 -140531
rect -80021 -140575 -79965 -140531
rect -79921 -140575 -79865 -140531
rect -79821 -140575 -79765 -140531
rect -79721 -140575 -79265 -140531
rect -79221 -140575 -79165 -140531
rect -79121 -140575 -79065 -140531
rect -79021 -140575 -78965 -140531
rect -78921 -140575 -78865 -140531
rect -78821 -140575 -78765 -140531
rect -78721 -140575 -78665 -140531
rect -78621 -140575 -78565 -140531
rect -78521 -140575 -78465 -140531
rect -78421 -140575 -78365 -140531
rect -78321 -140575 -78265 -140531
rect -78221 -140575 -78165 -140531
rect -78121 -140575 -78065 -140531
rect -78021 -140575 -77965 -140531
rect -77921 -140575 -77865 -140531
rect -77821 -140575 -77765 -140531
rect -77721 -140575 -77265 -140531
rect -77221 -140575 -77165 -140531
rect -77121 -140575 -77065 -140531
rect -77021 -140575 -76965 -140531
rect -76921 -140575 -76865 -140531
rect -76821 -140575 -76765 -140531
rect -76721 -140575 -76665 -140531
rect -76621 -140575 -76565 -140531
rect -76521 -140575 -76465 -140531
rect -76421 -140575 -76365 -140531
rect -76321 -140575 -76265 -140531
rect -76221 -140575 -76165 -140531
rect -76121 -140575 -76065 -140531
rect -76021 -140575 -75965 -140531
rect -75921 -140575 -75865 -140531
rect -75821 -140575 -75765 -140531
rect -75721 -140575 -71799 -140531
rect -87194 -140631 -71799 -140575
rect -87194 -140675 -83265 -140631
rect -83221 -140675 -83165 -140631
rect -83121 -140675 -83065 -140631
rect -83021 -140675 -82965 -140631
rect -82921 -140675 -82865 -140631
rect -82821 -140675 -82765 -140631
rect -82721 -140675 -82665 -140631
rect -82621 -140675 -82565 -140631
rect -82521 -140675 -82465 -140631
rect -82421 -140675 -82365 -140631
rect -82321 -140675 -82265 -140631
rect -82221 -140675 -82165 -140631
rect -82121 -140675 -82065 -140631
rect -82021 -140675 -81965 -140631
rect -81921 -140675 -81865 -140631
rect -81821 -140675 -81765 -140631
rect -81721 -140675 -81265 -140631
rect -81221 -140675 -81165 -140631
rect -81121 -140675 -81065 -140631
rect -81021 -140675 -80965 -140631
rect -80921 -140675 -80865 -140631
rect -80821 -140675 -80765 -140631
rect -80721 -140675 -80665 -140631
rect -80621 -140675 -80565 -140631
rect -80521 -140675 -80465 -140631
rect -80421 -140675 -80365 -140631
rect -80321 -140675 -80265 -140631
rect -80221 -140675 -80165 -140631
rect -80121 -140675 -80065 -140631
rect -80021 -140675 -79965 -140631
rect -79921 -140675 -79865 -140631
rect -79821 -140675 -79765 -140631
rect -79721 -140675 -79265 -140631
rect -79221 -140675 -79165 -140631
rect -79121 -140675 -79065 -140631
rect -79021 -140675 -78965 -140631
rect -78921 -140675 -78865 -140631
rect -78821 -140675 -78765 -140631
rect -78721 -140675 -78665 -140631
rect -78621 -140675 -78565 -140631
rect -78521 -140675 -78465 -140631
rect -78421 -140675 -78365 -140631
rect -78321 -140675 -78265 -140631
rect -78221 -140675 -78165 -140631
rect -78121 -140675 -78065 -140631
rect -78021 -140675 -77965 -140631
rect -77921 -140675 -77865 -140631
rect -77821 -140675 -77765 -140631
rect -77721 -140675 -77265 -140631
rect -77221 -140675 -77165 -140631
rect -77121 -140675 -77065 -140631
rect -77021 -140675 -76965 -140631
rect -76921 -140675 -76865 -140631
rect -76821 -140675 -76765 -140631
rect -76721 -140675 -76665 -140631
rect -76621 -140675 -76565 -140631
rect -76521 -140675 -76465 -140631
rect -76421 -140675 -76365 -140631
rect -76321 -140675 -76265 -140631
rect -76221 -140675 -76165 -140631
rect -76121 -140675 -76065 -140631
rect -76021 -140675 -75965 -140631
rect -75921 -140675 -75865 -140631
rect -75821 -140675 -75765 -140631
rect -75721 -140675 -71799 -140631
rect -87194 -140731 -71799 -140675
rect -87194 -140775 -83265 -140731
rect -83221 -140775 -83165 -140731
rect -83121 -140775 -83065 -140731
rect -83021 -140775 -82965 -140731
rect -82921 -140775 -82865 -140731
rect -82821 -140775 -82765 -140731
rect -82721 -140775 -82665 -140731
rect -82621 -140775 -82565 -140731
rect -82521 -140775 -82465 -140731
rect -82421 -140775 -82365 -140731
rect -82321 -140775 -82265 -140731
rect -82221 -140775 -82165 -140731
rect -82121 -140775 -82065 -140731
rect -82021 -140775 -81965 -140731
rect -81921 -140775 -81865 -140731
rect -81821 -140775 -81765 -140731
rect -81721 -140775 -81265 -140731
rect -81221 -140775 -81165 -140731
rect -81121 -140775 -81065 -140731
rect -81021 -140775 -80965 -140731
rect -80921 -140775 -80865 -140731
rect -80821 -140775 -80765 -140731
rect -80721 -140775 -80665 -140731
rect -80621 -140775 -80565 -140731
rect -80521 -140775 -80465 -140731
rect -80421 -140775 -80365 -140731
rect -80321 -140775 -80265 -140731
rect -80221 -140775 -80165 -140731
rect -80121 -140775 -80065 -140731
rect -80021 -140775 -79965 -140731
rect -79921 -140775 -79865 -140731
rect -79821 -140775 -79765 -140731
rect -79721 -140775 -79265 -140731
rect -79221 -140775 -79165 -140731
rect -79121 -140775 -79065 -140731
rect -79021 -140775 -78965 -140731
rect -78921 -140775 -78865 -140731
rect -78821 -140775 -78765 -140731
rect -78721 -140775 -78665 -140731
rect -78621 -140775 -78565 -140731
rect -78521 -140775 -78465 -140731
rect -78421 -140775 -78365 -140731
rect -78321 -140775 -78265 -140731
rect -78221 -140775 -78165 -140731
rect -78121 -140775 -78065 -140731
rect -78021 -140775 -77965 -140731
rect -77921 -140775 -77865 -140731
rect -77821 -140775 -77765 -140731
rect -77721 -140775 -77265 -140731
rect -77221 -140775 -77165 -140731
rect -77121 -140775 -77065 -140731
rect -77021 -140775 -76965 -140731
rect -76921 -140775 -76865 -140731
rect -76821 -140775 -76765 -140731
rect -76721 -140775 -76665 -140731
rect -76621 -140775 -76565 -140731
rect -76521 -140775 -76465 -140731
rect -76421 -140775 -76365 -140731
rect -76321 -140775 -76265 -140731
rect -76221 -140775 -76165 -140731
rect -76121 -140775 -76065 -140731
rect -76021 -140775 -75965 -140731
rect -75921 -140775 -75865 -140731
rect -75821 -140775 -75765 -140731
rect -75721 -140775 -71799 -140731
rect -87194 -140831 -71799 -140775
rect -87194 -140875 -83265 -140831
rect -83221 -140875 -83165 -140831
rect -83121 -140875 -83065 -140831
rect -83021 -140875 -82965 -140831
rect -82921 -140875 -82865 -140831
rect -82821 -140875 -82765 -140831
rect -82721 -140875 -82665 -140831
rect -82621 -140875 -82565 -140831
rect -82521 -140875 -82465 -140831
rect -82421 -140875 -82365 -140831
rect -82321 -140875 -82265 -140831
rect -82221 -140875 -82165 -140831
rect -82121 -140875 -82065 -140831
rect -82021 -140875 -81965 -140831
rect -81921 -140875 -81865 -140831
rect -81821 -140875 -81765 -140831
rect -81721 -140875 -81265 -140831
rect -81221 -140875 -81165 -140831
rect -81121 -140875 -81065 -140831
rect -81021 -140875 -80965 -140831
rect -80921 -140875 -80865 -140831
rect -80821 -140875 -80765 -140831
rect -80721 -140875 -80665 -140831
rect -80621 -140875 -80565 -140831
rect -80521 -140875 -80465 -140831
rect -80421 -140875 -80365 -140831
rect -80321 -140875 -80265 -140831
rect -80221 -140875 -80165 -140831
rect -80121 -140875 -80065 -140831
rect -80021 -140875 -79965 -140831
rect -79921 -140875 -79865 -140831
rect -79821 -140875 -79765 -140831
rect -79721 -140875 -79265 -140831
rect -79221 -140875 -79165 -140831
rect -79121 -140875 -79065 -140831
rect -79021 -140875 -78965 -140831
rect -78921 -140875 -78865 -140831
rect -78821 -140875 -78765 -140831
rect -78721 -140875 -78665 -140831
rect -78621 -140875 -78565 -140831
rect -78521 -140875 -78465 -140831
rect -78421 -140875 -78365 -140831
rect -78321 -140875 -78265 -140831
rect -78221 -140875 -78165 -140831
rect -78121 -140875 -78065 -140831
rect -78021 -140875 -77965 -140831
rect -77921 -140875 -77865 -140831
rect -77821 -140875 -77765 -140831
rect -77721 -140875 -77265 -140831
rect -77221 -140875 -77165 -140831
rect -77121 -140875 -77065 -140831
rect -77021 -140875 -76965 -140831
rect -76921 -140875 -76865 -140831
rect -76821 -140875 -76765 -140831
rect -76721 -140875 -76665 -140831
rect -76621 -140875 -76565 -140831
rect -76521 -140875 -76465 -140831
rect -76421 -140875 -76365 -140831
rect -76321 -140875 -76265 -140831
rect -76221 -140875 -76165 -140831
rect -76121 -140875 -76065 -140831
rect -76021 -140875 -75965 -140831
rect -75921 -140875 -75865 -140831
rect -75821 -140875 -75765 -140831
rect -75721 -140875 -71799 -140831
rect -87194 -140931 -71799 -140875
rect -87194 -140975 -83265 -140931
rect -83221 -140975 -83165 -140931
rect -83121 -140975 -83065 -140931
rect -83021 -140975 -82965 -140931
rect -82921 -140975 -82865 -140931
rect -82821 -140975 -82765 -140931
rect -82721 -140975 -82665 -140931
rect -82621 -140975 -82565 -140931
rect -82521 -140975 -82465 -140931
rect -82421 -140975 -82365 -140931
rect -82321 -140975 -82265 -140931
rect -82221 -140975 -82165 -140931
rect -82121 -140975 -82065 -140931
rect -82021 -140975 -81965 -140931
rect -81921 -140975 -81865 -140931
rect -81821 -140975 -81765 -140931
rect -81721 -140975 -81265 -140931
rect -81221 -140975 -81165 -140931
rect -81121 -140975 -81065 -140931
rect -81021 -140975 -80965 -140931
rect -80921 -140975 -80865 -140931
rect -80821 -140975 -80765 -140931
rect -80721 -140975 -80665 -140931
rect -80621 -140975 -80565 -140931
rect -80521 -140975 -80465 -140931
rect -80421 -140975 -80365 -140931
rect -80321 -140975 -80265 -140931
rect -80221 -140975 -80165 -140931
rect -80121 -140975 -80065 -140931
rect -80021 -140975 -79965 -140931
rect -79921 -140975 -79865 -140931
rect -79821 -140975 -79765 -140931
rect -79721 -140975 -79265 -140931
rect -79221 -140975 -79165 -140931
rect -79121 -140975 -79065 -140931
rect -79021 -140975 -78965 -140931
rect -78921 -140975 -78865 -140931
rect -78821 -140975 -78765 -140931
rect -78721 -140975 -78665 -140931
rect -78621 -140975 -78565 -140931
rect -78521 -140975 -78465 -140931
rect -78421 -140975 -78365 -140931
rect -78321 -140975 -78265 -140931
rect -78221 -140975 -78165 -140931
rect -78121 -140975 -78065 -140931
rect -78021 -140975 -77965 -140931
rect -77921 -140975 -77865 -140931
rect -77821 -140975 -77765 -140931
rect -77721 -140975 -77265 -140931
rect -77221 -140975 -77165 -140931
rect -77121 -140975 -77065 -140931
rect -77021 -140975 -76965 -140931
rect -76921 -140975 -76865 -140931
rect -76821 -140975 -76765 -140931
rect -76721 -140975 -76665 -140931
rect -76621 -140975 -76565 -140931
rect -76521 -140975 -76465 -140931
rect -76421 -140975 -76365 -140931
rect -76321 -140975 -76265 -140931
rect -76221 -140975 -76165 -140931
rect -76121 -140975 -76065 -140931
rect -76021 -140975 -75965 -140931
rect -75921 -140975 -75865 -140931
rect -75821 -140975 -75765 -140931
rect -75721 -140975 -71799 -140931
rect -87194 -141031 -71799 -140975
rect -87194 -141075 -83265 -141031
rect -83221 -141075 -83165 -141031
rect -83121 -141075 -83065 -141031
rect -83021 -141075 -82965 -141031
rect -82921 -141075 -82865 -141031
rect -82821 -141075 -82765 -141031
rect -82721 -141075 -82665 -141031
rect -82621 -141075 -82565 -141031
rect -82521 -141075 -82465 -141031
rect -82421 -141075 -82365 -141031
rect -82321 -141075 -82265 -141031
rect -82221 -141075 -82165 -141031
rect -82121 -141075 -82065 -141031
rect -82021 -141075 -81965 -141031
rect -81921 -141075 -81865 -141031
rect -81821 -141075 -81765 -141031
rect -81721 -141075 -81265 -141031
rect -81221 -141075 -81165 -141031
rect -81121 -141075 -81065 -141031
rect -81021 -141075 -80965 -141031
rect -80921 -141075 -80865 -141031
rect -80821 -141075 -80765 -141031
rect -80721 -141075 -80665 -141031
rect -80621 -141075 -80565 -141031
rect -80521 -141075 -80465 -141031
rect -80421 -141075 -80365 -141031
rect -80321 -141075 -80265 -141031
rect -80221 -141075 -80165 -141031
rect -80121 -141075 -80065 -141031
rect -80021 -141075 -79965 -141031
rect -79921 -141075 -79865 -141031
rect -79821 -141075 -79765 -141031
rect -79721 -141075 -79265 -141031
rect -79221 -141075 -79165 -141031
rect -79121 -141075 -79065 -141031
rect -79021 -141075 -78965 -141031
rect -78921 -141075 -78865 -141031
rect -78821 -141075 -78765 -141031
rect -78721 -141075 -78665 -141031
rect -78621 -141075 -78565 -141031
rect -78521 -141075 -78465 -141031
rect -78421 -141075 -78365 -141031
rect -78321 -141075 -78265 -141031
rect -78221 -141075 -78165 -141031
rect -78121 -141075 -78065 -141031
rect -78021 -141075 -77965 -141031
rect -77921 -141075 -77865 -141031
rect -77821 -141075 -77765 -141031
rect -77721 -141075 -77265 -141031
rect -77221 -141075 -77165 -141031
rect -77121 -141075 -77065 -141031
rect -77021 -141075 -76965 -141031
rect -76921 -141075 -76865 -141031
rect -76821 -141075 -76765 -141031
rect -76721 -141075 -76665 -141031
rect -76621 -141075 -76565 -141031
rect -76521 -141075 -76465 -141031
rect -76421 -141075 -76365 -141031
rect -76321 -141075 -76265 -141031
rect -76221 -141075 -76165 -141031
rect -76121 -141075 -76065 -141031
rect -76021 -141075 -75965 -141031
rect -75921 -141075 -75865 -141031
rect -75821 -141075 -75765 -141031
rect -75721 -141075 -71799 -141031
rect -87194 -141131 -71799 -141075
rect -87194 -141175 -83265 -141131
rect -83221 -141175 -83165 -141131
rect -83121 -141175 -83065 -141131
rect -83021 -141175 -82965 -141131
rect -82921 -141175 -82865 -141131
rect -82821 -141175 -82765 -141131
rect -82721 -141175 -82665 -141131
rect -82621 -141175 -82565 -141131
rect -82521 -141175 -82465 -141131
rect -82421 -141175 -82365 -141131
rect -82321 -141175 -82265 -141131
rect -82221 -141175 -82165 -141131
rect -82121 -141175 -82065 -141131
rect -82021 -141175 -81965 -141131
rect -81921 -141175 -81865 -141131
rect -81821 -141175 -81765 -141131
rect -81721 -141175 -81265 -141131
rect -81221 -141175 -81165 -141131
rect -81121 -141175 -81065 -141131
rect -81021 -141175 -80965 -141131
rect -80921 -141175 -80865 -141131
rect -80821 -141175 -80765 -141131
rect -80721 -141175 -80665 -141131
rect -80621 -141175 -80565 -141131
rect -80521 -141175 -80465 -141131
rect -80421 -141175 -80365 -141131
rect -80321 -141175 -80265 -141131
rect -80221 -141175 -80165 -141131
rect -80121 -141175 -80065 -141131
rect -80021 -141175 -79965 -141131
rect -79921 -141175 -79865 -141131
rect -79821 -141175 -79765 -141131
rect -79721 -141175 -79265 -141131
rect -79221 -141175 -79165 -141131
rect -79121 -141175 -79065 -141131
rect -79021 -141175 -78965 -141131
rect -78921 -141175 -78865 -141131
rect -78821 -141175 -78765 -141131
rect -78721 -141175 -78665 -141131
rect -78621 -141175 -78565 -141131
rect -78521 -141175 -78465 -141131
rect -78421 -141175 -78365 -141131
rect -78321 -141175 -78265 -141131
rect -78221 -141175 -78165 -141131
rect -78121 -141175 -78065 -141131
rect -78021 -141175 -77965 -141131
rect -77921 -141175 -77865 -141131
rect -77821 -141175 -77765 -141131
rect -77721 -141175 -77265 -141131
rect -77221 -141175 -77165 -141131
rect -77121 -141175 -77065 -141131
rect -77021 -141175 -76965 -141131
rect -76921 -141175 -76865 -141131
rect -76821 -141175 -76765 -141131
rect -76721 -141175 -76665 -141131
rect -76621 -141175 -76565 -141131
rect -76521 -141175 -76465 -141131
rect -76421 -141175 -76365 -141131
rect -76321 -141175 -76265 -141131
rect -76221 -141175 -76165 -141131
rect -76121 -141175 -76065 -141131
rect -76021 -141175 -75965 -141131
rect -75921 -141175 -75865 -141131
rect -75821 -141175 -75765 -141131
rect -75721 -141175 -71799 -141131
rect -87194 -141231 -71799 -141175
rect -87194 -141275 -83265 -141231
rect -83221 -141275 -83165 -141231
rect -83121 -141275 -83065 -141231
rect -83021 -141275 -82965 -141231
rect -82921 -141275 -82865 -141231
rect -82821 -141275 -82765 -141231
rect -82721 -141275 -82665 -141231
rect -82621 -141275 -82565 -141231
rect -82521 -141275 -82465 -141231
rect -82421 -141275 -82365 -141231
rect -82321 -141275 -82265 -141231
rect -82221 -141275 -82165 -141231
rect -82121 -141275 -82065 -141231
rect -82021 -141275 -81965 -141231
rect -81921 -141275 -81865 -141231
rect -81821 -141275 -81765 -141231
rect -81721 -141275 -81265 -141231
rect -81221 -141275 -81165 -141231
rect -81121 -141275 -81065 -141231
rect -81021 -141275 -80965 -141231
rect -80921 -141275 -80865 -141231
rect -80821 -141275 -80765 -141231
rect -80721 -141275 -80665 -141231
rect -80621 -141275 -80565 -141231
rect -80521 -141275 -80465 -141231
rect -80421 -141275 -80365 -141231
rect -80321 -141275 -80265 -141231
rect -80221 -141275 -80165 -141231
rect -80121 -141275 -80065 -141231
rect -80021 -141275 -79965 -141231
rect -79921 -141275 -79865 -141231
rect -79821 -141275 -79765 -141231
rect -79721 -141275 -79265 -141231
rect -79221 -141275 -79165 -141231
rect -79121 -141275 -79065 -141231
rect -79021 -141275 -78965 -141231
rect -78921 -141275 -78865 -141231
rect -78821 -141275 -78765 -141231
rect -78721 -141275 -78665 -141231
rect -78621 -141275 -78565 -141231
rect -78521 -141275 -78465 -141231
rect -78421 -141275 -78365 -141231
rect -78321 -141275 -78265 -141231
rect -78221 -141275 -78165 -141231
rect -78121 -141275 -78065 -141231
rect -78021 -141275 -77965 -141231
rect -77921 -141275 -77865 -141231
rect -77821 -141275 -77765 -141231
rect -77721 -141275 -77265 -141231
rect -77221 -141275 -77165 -141231
rect -77121 -141275 -77065 -141231
rect -77021 -141275 -76965 -141231
rect -76921 -141275 -76865 -141231
rect -76821 -141275 -76765 -141231
rect -76721 -141275 -76665 -141231
rect -76621 -141275 -76565 -141231
rect -76521 -141275 -76465 -141231
rect -76421 -141275 -76365 -141231
rect -76321 -141275 -76265 -141231
rect -76221 -141275 -76165 -141231
rect -76121 -141275 -76065 -141231
rect -76021 -141275 -75965 -141231
rect -75921 -141275 -75865 -141231
rect -75821 -141275 -75765 -141231
rect -75721 -141275 -71799 -141231
rect -87194 -141331 -71799 -141275
rect -87194 -141375 -83265 -141331
rect -83221 -141375 -83165 -141331
rect -83121 -141375 -83065 -141331
rect -83021 -141375 -82965 -141331
rect -82921 -141375 -82865 -141331
rect -82821 -141375 -82765 -141331
rect -82721 -141375 -82665 -141331
rect -82621 -141375 -82565 -141331
rect -82521 -141375 -82465 -141331
rect -82421 -141375 -82365 -141331
rect -82321 -141375 -82265 -141331
rect -82221 -141375 -82165 -141331
rect -82121 -141375 -82065 -141331
rect -82021 -141375 -81965 -141331
rect -81921 -141375 -81865 -141331
rect -81821 -141375 -81765 -141331
rect -81721 -141375 -81265 -141331
rect -81221 -141375 -81165 -141331
rect -81121 -141375 -81065 -141331
rect -81021 -141375 -80965 -141331
rect -80921 -141375 -80865 -141331
rect -80821 -141375 -80765 -141331
rect -80721 -141375 -80665 -141331
rect -80621 -141375 -80565 -141331
rect -80521 -141375 -80465 -141331
rect -80421 -141375 -80365 -141331
rect -80321 -141375 -80265 -141331
rect -80221 -141375 -80165 -141331
rect -80121 -141375 -80065 -141331
rect -80021 -141375 -79965 -141331
rect -79921 -141375 -79865 -141331
rect -79821 -141375 -79765 -141331
rect -79721 -141375 -79265 -141331
rect -79221 -141375 -79165 -141331
rect -79121 -141375 -79065 -141331
rect -79021 -141375 -78965 -141331
rect -78921 -141375 -78865 -141331
rect -78821 -141375 -78765 -141331
rect -78721 -141375 -78665 -141331
rect -78621 -141375 -78565 -141331
rect -78521 -141375 -78465 -141331
rect -78421 -141375 -78365 -141331
rect -78321 -141375 -78265 -141331
rect -78221 -141375 -78165 -141331
rect -78121 -141375 -78065 -141331
rect -78021 -141375 -77965 -141331
rect -77921 -141375 -77865 -141331
rect -77821 -141375 -77765 -141331
rect -77721 -141375 -77265 -141331
rect -77221 -141375 -77165 -141331
rect -77121 -141375 -77065 -141331
rect -77021 -141375 -76965 -141331
rect -76921 -141375 -76865 -141331
rect -76821 -141375 -76765 -141331
rect -76721 -141375 -76665 -141331
rect -76621 -141375 -76565 -141331
rect -76521 -141375 -76465 -141331
rect -76421 -141375 -76365 -141331
rect -76321 -141375 -76265 -141331
rect -76221 -141375 -76165 -141331
rect -76121 -141375 -76065 -141331
rect -76021 -141375 -75965 -141331
rect -75921 -141375 -75865 -141331
rect -75821 -141375 -75765 -141331
rect -75721 -141375 -71799 -141331
rect -87194 -141431 -71799 -141375
rect -87194 -141475 -83265 -141431
rect -83221 -141475 -83165 -141431
rect -83121 -141475 -83065 -141431
rect -83021 -141475 -82965 -141431
rect -82921 -141475 -82865 -141431
rect -82821 -141475 -82765 -141431
rect -82721 -141475 -82665 -141431
rect -82621 -141475 -82565 -141431
rect -82521 -141475 -82465 -141431
rect -82421 -141475 -82365 -141431
rect -82321 -141475 -82265 -141431
rect -82221 -141475 -82165 -141431
rect -82121 -141475 -82065 -141431
rect -82021 -141475 -81965 -141431
rect -81921 -141475 -81865 -141431
rect -81821 -141475 -81765 -141431
rect -81721 -141475 -81265 -141431
rect -81221 -141475 -81165 -141431
rect -81121 -141475 -81065 -141431
rect -81021 -141475 -80965 -141431
rect -80921 -141475 -80865 -141431
rect -80821 -141475 -80765 -141431
rect -80721 -141475 -80665 -141431
rect -80621 -141475 -80565 -141431
rect -80521 -141475 -80465 -141431
rect -80421 -141475 -80365 -141431
rect -80321 -141475 -80265 -141431
rect -80221 -141475 -80165 -141431
rect -80121 -141475 -80065 -141431
rect -80021 -141475 -79965 -141431
rect -79921 -141475 -79865 -141431
rect -79821 -141475 -79765 -141431
rect -79721 -141475 -79265 -141431
rect -79221 -141475 -79165 -141431
rect -79121 -141475 -79065 -141431
rect -79021 -141475 -78965 -141431
rect -78921 -141475 -78865 -141431
rect -78821 -141475 -78765 -141431
rect -78721 -141475 -78665 -141431
rect -78621 -141475 -78565 -141431
rect -78521 -141475 -78465 -141431
rect -78421 -141475 -78365 -141431
rect -78321 -141475 -78265 -141431
rect -78221 -141475 -78165 -141431
rect -78121 -141475 -78065 -141431
rect -78021 -141475 -77965 -141431
rect -77921 -141475 -77865 -141431
rect -77821 -141475 -77765 -141431
rect -77721 -141475 -77265 -141431
rect -77221 -141475 -77165 -141431
rect -77121 -141475 -77065 -141431
rect -77021 -141475 -76965 -141431
rect -76921 -141475 -76865 -141431
rect -76821 -141475 -76765 -141431
rect -76721 -141475 -76665 -141431
rect -76621 -141475 -76565 -141431
rect -76521 -141475 -76465 -141431
rect -76421 -141475 -76365 -141431
rect -76321 -141475 -76265 -141431
rect -76221 -141475 -76165 -141431
rect -76121 -141475 -76065 -141431
rect -76021 -141475 -75965 -141431
rect -75921 -141475 -75865 -141431
rect -75821 -141475 -75765 -141431
rect -75721 -141475 -71799 -141431
rect -87194 -141531 -71799 -141475
rect -87194 -141575 -83265 -141531
rect -83221 -141575 -83165 -141531
rect -83121 -141575 -83065 -141531
rect -83021 -141575 -82965 -141531
rect -82921 -141575 -82865 -141531
rect -82821 -141575 -82765 -141531
rect -82721 -141575 -82665 -141531
rect -82621 -141575 -82565 -141531
rect -82521 -141575 -82465 -141531
rect -82421 -141575 -82365 -141531
rect -82321 -141575 -82265 -141531
rect -82221 -141575 -82165 -141531
rect -82121 -141575 -82065 -141531
rect -82021 -141575 -81965 -141531
rect -81921 -141575 -81865 -141531
rect -81821 -141575 -81765 -141531
rect -81721 -141575 -81265 -141531
rect -81221 -141575 -81165 -141531
rect -81121 -141575 -81065 -141531
rect -81021 -141575 -80965 -141531
rect -80921 -141575 -80865 -141531
rect -80821 -141575 -80765 -141531
rect -80721 -141575 -80665 -141531
rect -80621 -141575 -80565 -141531
rect -80521 -141575 -80465 -141531
rect -80421 -141575 -80365 -141531
rect -80321 -141575 -80265 -141531
rect -80221 -141575 -80165 -141531
rect -80121 -141575 -80065 -141531
rect -80021 -141575 -79965 -141531
rect -79921 -141575 -79865 -141531
rect -79821 -141575 -79765 -141531
rect -79721 -141575 -79265 -141531
rect -79221 -141575 -79165 -141531
rect -79121 -141575 -79065 -141531
rect -79021 -141575 -78965 -141531
rect -78921 -141575 -78865 -141531
rect -78821 -141575 -78765 -141531
rect -78721 -141575 -78665 -141531
rect -78621 -141575 -78565 -141531
rect -78521 -141575 -78465 -141531
rect -78421 -141575 -78365 -141531
rect -78321 -141575 -78265 -141531
rect -78221 -141575 -78165 -141531
rect -78121 -141575 -78065 -141531
rect -78021 -141575 -77965 -141531
rect -77921 -141575 -77865 -141531
rect -77821 -141575 -77765 -141531
rect -77721 -141575 -77265 -141531
rect -77221 -141575 -77165 -141531
rect -77121 -141575 -77065 -141531
rect -77021 -141575 -76965 -141531
rect -76921 -141575 -76865 -141531
rect -76821 -141575 -76765 -141531
rect -76721 -141575 -76665 -141531
rect -76621 -141575 -76565 -141531
rect -76521 -141575 -76465 -141531
rect -76421 -141575 -76365 -141531
rect -76321 -141575 -76265 -141531
rect -76221 -141575 -76165 -141531
rect -76121 -141575 -76065 -141531
rect -76021 -141575 -75965 -141531
rect -75921 -141575 -75865 -141531
rect -75821 -141575 -75765 -141531
rect -75721 -141575 -71799 -141531
rect -87194 -141631 -71799 -141575
rect -87194 -141675 -83265 -141631
rect -83221 -141675 -83165 -141631
rect -83121 -141675 -83065 -141631
rect -83021 -141675 -82965 -141631
rect -82921 -141675 -82865 -141631
rect -82821 -141675 -82765 -141631
rect -82721 -141675 -82665 -141631
rect -82621 -141675 -82565 -141631
rect -82521 -141675 -82465 -141631
rect -82421 -141675 -82365 -141631
rect -82321 -141675 -82265 -141631
rect -82221 -141675 -82165 -141631
rect -82121 -141675 -82065 -141631
rect -82021 -141675 -81965 -141631
rect -81921 -141675 -81865 -141631
rect -81821 -141675 -81765 -141631
rect -81721 -141675 -81265 -141631
rect -81221 -141675 -81165 -141631
rect -81121 -141675 -81065 -141631
rect -81021 -141675 -80965 -141631
rect -80921 -141675 -80865 -141631
rect -80821 -141675 -80765 -141631
rect -80721 -141675 -80665 -141631
rect -80621 -141675 -80565 -141631
rect -80521 -141675 -80465 -141631
rect -80421 -141675 -80365 -141631
rect -80321 -141675 -80265 -141631
rect -80221 -141675 -80165 -141631
rect -80121 -141675 -80065 -141631
rect -80021 -141675 -79965 -141631
rect -79921 -141675 -79865 -141631
rect -79821 -141675 -79765 -141631
rect -79721 -141675 -79265 -141631
rect -79221 -141675 -79165 -141631
rect -79121 -141675 -79065 -141631
rect -79021 -141675 -78965 -141631
rect -78921 -141675 -78865 -141631
rect -78821 -141675 -78765 -141631
rect -78721 -141675 -78665 -141631
rect -78621 -141675 -78565 -141631
rect -78521 -141675 -78465 -141631
rect -78421 -141675 -78365 -141631
rect -78321 -141675 -78265 -141631
rect -78221 -141675 -78165 -141631
rect -78121 -141675 -78065 -141631
rect -78021 -141675 -77965 -141631
rect -77921 -141675 -77865 -141631
rect -77821 -141675 -77765 -141631
rect -77721 -141675 -77265 -141631
rect -77221 -141675 -77165 -141631
rect -77121 -141675 -77065 -141631
rect -77021 -141675 -76965 -141631
rect -76921 -141675 -76865 -141631
rect -76821 -141675 -76765 -141631
rect -76721 -141675 -76665 -141631
rect -76621 -141675 -76565 -141631
rect -76521 -141675 -76465 -141631
rect -76421 -141675 -76365 -141631
rect -76321 -141675 -76265 -141631
rect -76221 -141675 -76165 -141631
rect -76121 -141675 -76065 -141631
rect -76021 -141675 -75965 -141631
rect -75921 -141675 -75865 -141631
rect -75821 -141675 -75765 -141631
rect -75721 -141675 -71799 -141631
rect -87194 -141731 -71799 -141675
rect -87194 -141775 -83265 -141731
rect -83221 -141775 -83165 -141731
rect -83121 -141775 -83065 -141731
rect -83021 -141775 -82965 -141731
rect -82921 -141775 -82865 -141731
rect -82821 -141775 -82765 -141731
rect -82721 -141775 -82665 -141731
rect -82621 -141775 -82565 -141731
rect -82521 -141775 -82465 -141731
rect -82421 -141775 -82365 -141731
rect -82321 -141775 -82265 -141731
rect -82221 -141775 -82165 -141731
rect -82121 -141775 -82065 -141731
rect -82021 -141775 -81965 -141731
rect -81921 -141775 -81865 -141731
rect -81821 -141775 -81765 -141731
rect -81721 -141775 -81265 -141731
rect -81221 -141775 -81165 -141731
rect -81121 -141775 -81065 -141731
rect -81021 -141775 -80965 -141731
rect -80921 -141775 -80865 -141731
rect -80821 -141775 -80765 -141731
rect -80721 -141775 -80665 -141731
rect -80621 -141775 -80565 -141731
rect -80521 -141775 -80465 -141731
rect -80421 -141775 -80365 -141731
rect -80321 -141775 -80265 -141731
rect -80221 -141775 -80165 -141731
rect -80121 -141775 -80065 -141731
rect -80021 -141775 -79965 -141731
rect -79921 -141775 -79865 -141731
rect -79821 -141775 -79765 -141731
rect -79721 -141775 -79265 -141731
rect -79221 -141775 -79165 -141731
rect -79121 -141775 -79065 -141731
rect -79021 -141775 -78965 -141731
rect -78921 -141775 -78865 -141731
rect -78821 -141775 -78765 -141731
rect -78721 -141775 -78665 -141731
rect -78621 -141775 -78565 -141731
rect -78521 -141775 -78465 -141731
rect -78421 -141775 -78365 -141731
rect -78321 -141775 -78265 -141731
rect -78221 -141775 -78165 -141731
rect -78121 -141775 -78065 -141731
rect -78021 -141775 -77965 -141731
rect -77921 -141775 -77865 -141731
rect -77821 -141775 -77765 -141731
rect -77721 -141775 -77265 -141731
rect -77221 -141775 -77165 -141731
rect -77121 -141775 -77065 -141731
rect -77021 -141775 -76965 -141731
rect -76921 -141775 -76865 -141731
rect -76821 -141775 -76765 -141731
rect -76721 -141775 -76665 -141731
rect -76621 -141775 -76565 -141731
rect -76521 -141775 -76465 -141731
rect -76421 -141775 -76365 -141731
rect -76321 -141775 -76265 -141731
rect -76221 -141775 -76165 -141731
rect -76121 -141775 -76065 -141731
rect -76021 -141775 -75965 -141731
rect -75921 -141775 -75865 -141731
rect -75821 -141775 -75765 -141731
rect -75721 -141775 -71799 -141731
rect -87194 -144989 -71799 -141775
rect 81061 -137966 89740 -136015
rect 81061 -138010 81632 -137966
rect 81676 -138010 81732 -137966
rect 81776 -138010 81832 -137966
rect 81876 -138010 81932 -137966
rect 81976 -138010 82032 -137966
rect 82076 -138010 82132 -137966
rect 82176 -138010 82232 -137966
rect 82276 -138010 82332 -137966
rect 82376 -138010 82432 -137966
rect 82476 -138010 82532 -137966
rect 82576 -138010 82632 -137966
rect 82676 -138010 82732 -137966
rect 82776 -138010 82832 -137966
rect 82876 -138010 82932 -137966
rect 82976 -138010 83032 -137966
rect 83076 -138010 83132 -137966
rect 83176 -138010 83632 -137966
rect 83676 -138010 83732 -137966
rect 83776 -138010 83832 -137966
rect 83876 -138010 83932 -137966
rect 83976 -138010 84032 -137966
rect 84076 -138010 84132 -137966
rect 84176 -138010 84232 -137966
rect 84276 -138010 84332 -137966
rect 84376 -138010 84432 -137966
rect 84476 -138010 84532 -137966
rect 84576 -138010 84632 -137966
rect 84676 -138010 84732 -137966
rect 84776 -138010 84832 -137966
rect 84876 -138010 84932 -137966
rect 84976 -138010 85032 -137966
rect 85076 -138010 85132 -137966
rect 85176 -138010 85632 -137966
rect 85676 -138010 85732 -137966
rect 85776 -138010 85832 -137966
rect 85876 -138010 85932 -137966
rect 85976 -138010 86032 -137966
rect 86076 -138010 86132 -137966
rect 86176 -138010 86232 -137966
rect 86276 -138010 86332 -137966
rect 86376 -138010 86432 -137966
rect 86476 -138010 86532 -137966
rect 86576 -138010 86632 -137966
rect 86676 -138010 86732 -137966
rect 86776 -138010 86832 -137966
rect 86876 -138010 86932 -137966
rect 86976 -138010 87032 -137966
rect 87076 -138010 87132 -137966
rect 87176 -138010 87632 -137966
rect 87676 -138010 87732 -137966
rect 87776 -138010 87832 -137966
rect 87876 -138010 87932 -137966
rect 87976 -138010 88032 -137966
rect 88076 -138010 88132 -137966
rect 88176 -138010 88232 -137966
rect 88276 -138010 88332 -137966
rect 88376 -138010 88432 -137966
rect 88476 -138010 88532 -137966
rect 88576 -138010 88632 -137966
rect 88676 -138010 88732 -137966
rect 88776 -138010 88832 -137966
rect 88876 -138010 88932 -137966
rect 88976 -138010 89032 -137966
rect 89076 -138010 89132 -137966
rect 89176 -138010 89740 -137966
rect 81061 -138066 89740 -138010
rect 81061 -138110 81632 -138066
rect 81676 -138110 81732 -138066
rect 81776 -138110 81832 -138066
rect 81876 -138110 81932 -138066
rect 81976 -138110 82032 -138066
rect 82076 -138110 82132 -138066
rect 82176 -138110 82232 -138066
rect 82276 -138110 82332 -138066
rect 82376 -138110 82432 -138066
rect 82476 -138110 82532 -138066
rect 82576 -138110 82632 -138066
rect 82676 -138110 82732 -138066
rect 82776 -138110 82832 -138066
rect 82876 -138110 82932 -138066
rect 82976 -138110 83032 -138066
rect 83076 -138110 83132 -138066
rect 83176 -138110 83632 -138066
rect 83676 -138110 83732 -138066
rect 83776 -138110 83832 -138066
rect 83876 -138110 83932 -138066
rect 83976 -138110 84032 -138066
rect 84076 -138110 84132 -138066
rect 84176 -138110 84232 -138066
rect 84276 -138110 84332 -138066
rect 84376 -138110 84432 -138066
rect 84476 -138110 84532 -138066
rect 84576 -138110 84632 -138066
rect 84676 -138110 84732 -138066
rect 84776 -138110 84832 -138066
rect 84876 -138110 84932 -138066
rect 84976 -138110 85032 -138066
rect 85076 -138110 85132 -138066
rect 85176 -138110 85632 -138066
rect 85676 -138110 85732 -138066
rect 85776 -138110 85832 -138066
rect 85876 -138110 85932 -138066
rect 85976 -138110 86032 -138066
rect 86076 -138110 86132 -138066
rect 86176 -138110 86232 -138066
rect 86276 -138110 86332 -138066
rect 86376 -138110 86432 -138066
rect 86476 -138110 86532 -138066
rect 86576 -138110 86632 -138066
rect 86676 -138110 86732 -138066
rect 86776 -138110 86832 -138066
rect 86876 -138110 86932 -138066
rect 86976 -138110 87032 -138066
rect 87076 -138110 87132 -138066
rect 87176 -138110 87632 -138066
rect 87676 -138110 87732 -138066
rect 87776 -138110 87832 -138066
rect 87876 -138110 87932 -138066
rect 87976 -138110 88032 -138066
rect 88076 -138110 88132 -138066
rect 88176 -138110 88232 -138066
rect 88276 -138110 88332 -138066
rect 88376 -138110 88432 -138066
rect 88476 -138110 88532 -138066
rect 88576 -138110 88632 -138066
rect 88676 -138110 88732 -138066
rect 88776 -138110 88832 -138066
rect 88876 -138110 88932 -138066
rect 88976 -138110 89032 -138066
rect 89076 -138110 89132 -138066
rect 89176 -138110 89740 -138066
rect 81061 -138166 89740 -138110
rect 81061 -138210 81632 -138166
rect 81676 -138210 81732 -138166
rect 81776 -138210 81832 -138166
rect 81876 -138210 81932 -138166
rect 81976 -138210 82032 -138166
rect 82076 -138210 82132 -138166
rect 82176 -138210 82232 -138166
rect 82276 -138210 82332 -138166
rect 82376 -138210 82432 -138166
rect 82476 -138210 82532 -138166
rect 82576 -138210 82632 -138166
rect 82676 -138210 82732 -138166
rect 82776 -138210 82832 -138166
rect 82876 -138210 82932 -138166
rect 82976 -138210 83032 -138166
rect 83076 -138210 83132 -138166
rect 83176 -138210 83632 -138166
rect 83676 -138210 83732 -138166
rect 83776 -138210 83832 -138166
rect 83876 -138210 83932 -138166
rect 83976 -138210 84032 -138166
rect 84076 -138210 84132 -138166
rect 84176 -138210 84232 -138166
rect 84276 -138210 84332 -138166
rect 84376 -138210 84432 -138166
rect 84476 -138210 84532 -138166
rect 84576 -138210 84632 -138166
rect 84676 -138210 84732 -138166
rect 84776 -138210 84832 -138166
rect 84876 -138210 84932 -138166
rect 84976 -138210 85032 -138166
rect 85076 -138210 85132 -138166
rect 85176 -138210 85632 -138166
rect 85676 -138210 85732 -138166
rect 85776 -138210 85832 -138166
rect 85876 -138210 85932 -138166
rect 85976 -138210 86032 -138166
rect 86076 -138210 86132 -138166
rect 86176 -138210 86232 -138166
rect 86276 -138210 86332 -138166
rect 86376 -138210 86432 -138166
rect 86476 -138210 86532 -138166
rect 86576 -138210 86632 -138166
rect 86676 -138210 86732 -138166
rect 86776 -138210 86832 -138166
rect 86876 -138210 86932 -138166
rect 86976 -138210 87032 -138166
rect 87076 -138210 87132 -138166
rect 87176 -138210 87632 -138166
rect 87676 -138210 87732 -138166
rect 87776 -138210 87832 -138166
rect 87876 -138210 87932 -138166
rect 87976 -138210 88032 -138166
rect 88076 -138210 88132 -138166
rect 88176 -138210 88232 -138166
rect 88276 -138210 88332 -138166
rect 88376 -138210 88432 -138166
rect 88476 -138210 88532 -138166
rect 88576 -138210 88632 -138166
rect 88676 -138210 88732 -138166
rect 88776 -138210 88832 -138166
rect 88876 -138210 88932 -138166
rect 88976 -138210 89032 -138166
rect 89076 -138210 89132 -138166
rect 89176 -138210 89740 -138166
rect 81061 -138266 89740 -138210
rect 81061 -138310 81632 -138266
rect 81676 -138310 81732 -138266
rect 81776 -138310 81832 -138266
rect 81876 -138310 81932 -138266
rect 81976 -138310 82032 -138266
rect 82076 -138310 82132 -138266
rect 82176 -138310 82232 -138266
rect 82276 -138310 82332 -138266
rect 82376 -138310 82432 -138266
rect 82476 -138310 82532 -138266
rect 82576 -138310 82632 -138266
rect 82676 -138310 82732 -138266
rect 82776 -138310 82832 -138266
rect 82876 -138310 82932 -138266
rect 82976 -138310 83032 -138266
rect 83076 -138310 83132 -138266
rect 83176 -138310 83632 -138266
rect 83676 -138310 83732 -138266
rect 83776 -138310 83832 -138266
rect 83876 -138310 83932 -138266
rect 83976 -138310 84032 -138266
rect 84076 -138310 84132 -138266
rect 84176 -138310 84232 -138266
rect 84276 -138310 84332 -138266
rect 84376 -138310 84432 -138266
rect 84476 -138310 84532 -138266
rect 84576 -138310 84632 -138266
rect 84676 -138310 84732 -138266
rect 84776 -138310 84832 -138266
rect 84876 -138310 84932 -138266
rect 84976 -138310 85032 -138266
rect 85076 -138310 85132 -138266
rect 85176 -138310 85632 -138266
rect 85676 -138310 85732 -138266
rect 85776 -138310 85832 -138266
rect 85876 -138310 85932 -138266
rect 85976 -138310 86032 -138266
rect 86076 -138310 86132 -138266
rect 86176 -138310 86232 -138266
rect 86276 -138310 86332 -138266
rect 86376 -138310 86432 -138266
rect 86476 -138310 86532 -138266
rect 86576 -138310 86632 -138266
rect 86676 -138310 86732 -138266
rect 86776 -138310 86832 -138266
rect 86876 -138310 86932 -138266
rect 86976 -138310 87032 -138266
rect 87076 -138310 87132 -138266
rect 87176 -138310 87632 -138266
rect 87676 -138310 87732 -138266
rect 87776 -138310 87832 -138266
rect 87876 -138310 87932 -138266
rect 87976 -138310 88032 -138266
rect 88076 -138310 88132 -138266
rect 88176 -138310 88232 -138266
rect 88276 -138310 88332 -138266
rect 88376 -138310 88432 -138266
rect 88476 -138310 88532 -138266
rect 88576 -138310 88632 -138266
rect 88676 -138310 88732 -138266
rect 88776 -138310 88832 -138266
rect 88876 -138310 88932 -138266
rect 88976 -138310 89032 -138266
rect 89076 -138310 89132 -138266
rect 89176 -138310 89740 -138266
rect 81061 -138366 89740 -138310
rect 81061 -138410 81632 -138366
rect 81676 -138410 81732 -138366
rect 81776 -138410 81832 -138366
rect 81876 -138410 81932 -138366
rect 81976 -138410 82032 -138366
rect 82076 -138410 82132 -138366
rect 82176 -138410 82232 -138366
rect 82276 -138410 82332 -138366
rect 82376 -138410 82432 -138366
rect 82476 -138410 82532 -138366
rect 82576 -138410 82632 -138366
rect 82676 -138410 82732 -138366
rect 82776 -138410 82832 -138366
rect 82876 -138410 82932 -138366
rect 82976 -138410 83032 -138366
rect 83076 -138410 83132 -138366
rect 83176 -138410 83632 -138366
rect 83676 -138410 83732 -138366
rect 83776 -138410 83832 -138366
rect 83876 -138410 83932 -138366
rect 83976 -138410 84032 -138366
rect 84076 -138410 84132 -138366
rect 84176 -138410 84232 -138366
rect 84276 -138410 84332 -138366
rect 84376 -138410 84432 -138366
rect 84476 -138410 84532 -138366
rect 84576 -138410 84632 -138366
rect 84676 -138410 84732 -138366
rect 84776 -138410 84832 -138366
rect 84876 -138410 84932 -138366
rect 84976 -138410 85032 -138366
rect 85076 -138410 85132 -138366
rect 85176 -138410 85632 -138366
rect 85676 -138410 85732 -138366
rect 85776 -138410 85832 -138366
rect 85876 -138410 85932 -138366
rect 85976 -138410 86032 -138366
rect 86076 -138410 86132 -138366
rect 86176 -138410 86232 -138366
rect 86276 -138410 86332 -138366
rect 86376 -138410 86432 -138366
rect 86476 -138410 86532 -138366
rect 86576 -138410 86632 -138366
rect 86676 -138410 86732 -138366
rect 86776 -138410 86832 -138366
rect 86876 -138410 86932 -138366
rect 86976 -138410 87032 -138366
rect 87076 -138410 87132 -138366
rect 87176 -138410 87632 -138366
rect 87676 -138410 87732 -138366
rect 87776 -138410 87832 -138366
rect 87876 -138410 87932 -138366
rect 87976 -138410 88032 -138366
rect 88076 -138410 88132 -138366
rect 88176 -138410 88232 -138366
rect 88276 -138410 88332 -138366
rect 88376 -138410 88432 -138366
rect 88476 -138410 88532 -138366
rect 88576 -138410 88632 -138366
rect 88676 -138410 88732 -138366
rect 88776 -138410 88832 -138366
rect 88876 -138410 88932 -138366
rect 88976 -138410 89032 -138366
rect 89076 -138410 89132 -138366
rect 89176 -138410 89740 -138366
rect 81061 -138466 89740 -138410
rect 81061 -138510 81632 -138466
rect 81676 -138510 81732 -138466
rect 81776 -138510 81832 -138466
rect 81876 -138510 81932 -138466
rect 81976 -138510 82032 -138466
rect 82076 -138510 82132 -138466
rect 82176 -138510 82232 -138466
rect 82276 -138510 82332 -138466
rect 82376 -138510 82432 -138466
rect 82476 -138510 82532 -138466
rect 82576 -138510 82632 -138466
rect 82676 -138510 82732 -138466
rect 82776 -138510 82832 -138466
rect 82876 -138510 82932 -138466
rect 82976 -138510 83032 -138466
rect 83076 -138510 83132 -138466
rect 83176 -138510 83632 -138466
rect 83676 -138510 83732 -138466
rect 83776 -138510 83832 -138466
rect 83876 -138510 83932 -138466
rect 83976 -138510 84032 -138466
rect 84076 -138510 84132 -138466
rect 84176 -138510 84232 -138466
rect 84276 -138510 84332 -138466
rect 84376 -138510 84432 -138466
rect 84476 -138510 84532 -138466
rect 84576 -138510 84632 -138466
rect 84676 -138510 84732 -138466
rect 84776 -138510 84832 -138466
rect 84876 -138510 84932 -138466
rect 84976 -138510 85032 -138466
rect 85076 -138510 85132 -138466
rect 85176 -138510 85632 -138466
rect 85676 -138510 85732 -138466
rect 85776 -138510 85832 -138466
rect 85876 -138510 85932 -138466
rect 85976 -138510 86032 -138466
rect 86076 -138510 86132 -138466
rect 86176 -138510 86232 -138466
rect 86276 -138510 86332 -138466
rect 86376 -138510 86432 -138466
rect 86476 -138510 86532 -138466
rect 86576 -138510 86632 -138466
rect 86676 -138510 86732 -138466
rect 86776 -138510 86832 -138466
rect 86876 -138510 86932 -138466
rect 86976 -138510 87032 -138466
rect 87076 -138510 87132 -138466
rect 87176 -138510 87632 -138466
rect 87676 -138510 87732 -138466
rect 87776 -138510 87832 -138466
rect 87876 -138510 87932 -138466
rect 87976 -138510 88032 -138466
rect 88076 -138510 88132 -138466
rect 88176 -138510 88232 -138466
rect 88276 -138510 88332 -138466
rect 88376 -138510 88432 -138466
rect 88476 -138510 88532 -138466
rect 88576 -138510 88632 -138466
rect 88676 -138510 88732 -138466
rect 88776 -138510 88832 -138466
rect 88876 -138510 88932 -138466
rect 88976 -138510 89032 -138466
rect 89076 -138510 89132 -138466
rect 89176 -138510 89740 -138466
rect 81061 -138566 89740 -138510
rect 81061 -138610 81632 -138566
rect 81676 -138610 81732 -138566
rect 81776 -138610 81832 -138566
rect 81876 -138610 81932 -138566
rect 81976 -138610 82032 -138566
rect 82076 -138610 82132 -138566
rect 82176 -138610 82232 -138566
rect 82276 -138610 82332 -138566
rect 82376 -138610 82432 -138566
rect 82476 -138610 82532 -138566
rect 82576 -138610 82632 -138566
rect 82676 -138610 82732 -138566
rect 82776 -138610 82832 -138566
rect 82876 -138610 82932 -138566
rect 82976 -138610 83032 -138566
rect 83076 -138610 83132 -138566
rect 83176 -138610 83632 -138566
rect 83676 -138610 83732 -138566
rect 83776 -138610 83832 -138566
rect 83876 -138610 83932 -138566
rect 83976 -138610 84032 -138566
rect 84076 -138610 84132 -138566
rect 84176 -138610 84232 -138566
rect 84276 -138610 84332 -138566
rect 84376 -138610 84432 -138566
rect 84476 -138610 84532 -138566
rect 84576 -138610 84632 -138566
rect 84676 -138610 84732 -138566
rect 84776 -138610 84832 -138566
rect 84876 -138610 84932 -138566
rect 84976 -138610 85032 -138566
rect 85076 -138610 85132 -138566
rect 85176 -138610 85632 -138566
rect 85676 -138610 85732 -138566
rect 85776 -138610 85832 -138566
rect 85876 -138610 85932 -138566
rect 85976 -138610 86032 -138566
rect 86076 -138610 86132 -138566
rect 86176 -138610 86232 -138566
rect 86276 -138610 86332 -138566
rect 86376 -138610 86432 -138566
rect 86476 -138610 86532 -138566
rect 86576 -138610 86632 -138566
rect 86676 -138610 86732 -138566
rect 86776 -138610 86832 -138566
rect 86876 -138610 86932 -138566
rect 86976 -138610 87032 -138566
rect 87076 -138610 87132 -138566
rect 87176 -138610 87632 -138566
rect 87676 -138610 87732 -138566
rect 87776 -138610 87832 -138566
rect 87876 -138610 87932 -138566
rect 87976 -138610 88032 -138566
rect 88076 -138610 88132 -138566
rect 88176 -138610 88232 -138566
rect 88276 -138610 88332 -138566
rect 88376 -138610 88432 -138566
rect 88476 -138610 88532 -138566
rect 88576 -138610 88632 -138566
rect 88676 -138610 88732 -138566
rect 88776 -138610 88832 -138566
rect 88876 -138610 88932 -138566
rect 88976 -138610 89032 -138566
rect 89076 -138610 89132 -138566
rect 89176 -138610 89740 -138566
rect 81061 -138666 89740 -138610
rect 81061 -138710 81632 -138666
rect 81676 -138710 81732 -138666
rect 81776 -138710 81832 -138666
rect 81876 -138710 81932 -138666
rect 81976 -138710 82032 -138666
rect 82076 -138710 82132 -138666
rect 82176 -138710 82232 -138666
rect 82276 -138710 82332 -138666
rect 82376 -138710 82432 -138666
rect 82476 -138710 82532 -138666
rect 82576 -138710 82632 -138666
rect 82676 -138710 82732 -138666
rect 82776 -138710 82832 -138666
rect 82876 -138710 82932 -138666
rect 82976 -138710 83032 -138666
rect 83076 -138710 83132 -138666
rect 83176 -138710 83632 -138666
rect 83676 -138710 83732 -138666
rect 83776 -138710 83832 -138666
rect 83876 -138710 83932 -138666
rect 83976 -138710 84032 -138666
rect 84076 -138710 84132 -138666
rect 84176 -138710 84232 -138666
rect 84276 -138710 84332 -138666
rect 84376 -138710 84432 -138666
rect 84476 -138710 84532 -138666
rect 84576 -138710 84632 -138666
rect 84676 -138710 84732 -138666
rect 84776 -138710 84832 -138666
rect 84876 -138710 84932 -138666
rect 84976 -138710 85032 -138666
rect 85076 -138710 85132 -138666
rect 85176 -138710 85632 -138666
rect 85676 -138710 85732 -138666
rect 85776 -138710 85832 -138666
rect 85876 -138710 85932 -138666
rect 85976 -138710 86032 -138666
rect 86076 -138710 86132 -138666
rect 86176 -138710 86232 -138666
rect 86276 -138710 86332 -138666
rect 86376 -138710 86432 -138666
rect 86476 -138710 86532 -138666
rect 86576 -138710 86632 -138666
rect 86676 -138710 86732 -138666
rect 86776 -138710 86832 -138666
rect 86876 -138710 86932 -138666
rect 86976 -138710 87032 -138666
rect 87076 -138710 87132 -138666
rect 87176 -138710 87632 -138666
rect 87676 -138710 87732 -138666
rect 87776 -138710 87832 -138666
rect 87876 -138710 87932 -138666
rect 87976 -138710 88032 -138666
rect 88076 -138710 88132 -138666
rect 88176 -138710 88232 -138666
rect 88276 -138710 88332 -138666
rect 88376 -138710 88432 -138666
rect 88476 -138710 88532 -138666
rect 88576 -138710 88632 -138666
rect 88676 -138710 88732 -138666
rect 88776 -138710 88832 -138666
rect 88876 -138710 88932 -138666
rect 88976 -138710 89032 -138666
rect 89076 -138710 89132 -138666
rect 89176 -138710 89740 -138666
rect 81061 -138766 89740 -138710
rect 81061 -138810 81632 -138766
rect 81676 -138810 81732 -138766
rect 81776 -138810 81832 -138766
rect 81876 -138810 81932 -138766
rect 81976 -138810 82032 -138766
rect 82076 -138810 82132 -138766
rect 82176 -138810 82232 -138766
rect 82276 -138810 82332 -138766
rect 82376 -138810 82432 -138766
rect 82476 -138810 82532 -138766
rect 82576 -138810 82632 -138766
rect 82676 -138810 82732 -138766
rect 82776 -138810 82832 -138766
rect 82876 -138810 82932 -138766
rect 82976 -138810 83032 -138766
rect 83076 -138810 83132 -138766
rect 83176 -138810 83632 -138766
rect 83676 -138810 83732 -138766
rect 83776 -138810 83832 -138766
rect 83876 -138810 83932 -138766
rect 83976 -138810 84032 -138766
rect 84076 -138810 84132 -138766
rect 84176 -138810 84232 -138766
rect 84276 -138810 84332 -138766
rect 84376 -138810 84432 -138766
rect 84476 -138810 84532 -138766
rect 84576 -138810 84632 -138766
rect 84676 -138810 84732 -138766
rect 84776 -138810 84832 -138766
rect 84876 -138810 84932 -138766
rect 84976 -138810 85032 -138766
rect 85076 -138810 85132 -138766
rect 85176 -138810 85632 -138766
rect 85676 -138810 85732 -138766
rect 85776 -138810 85832 -138766
rect 85876 -138810 85932 -138766
rect 85976 -138810 86032 -138766
rect 86076 -138810 86132 -138766
rect 86176 -138810 86232 -138766
rect 86276 -138810 86332 -138766
rect 86376 -138810 86432 -138766
rect 86476 -138810 86532 -138766
rect 86576 -138810 86632 -138766
rect 86676 -138810 86732 -138766
rect 86776 -138810 86832 -138766
rect 86876 -138810 86932 -138766
rect 86976 -138810 87032 -138766
rect 87076 -138810 87132 -138766
rect 87176 -138810 87632 -138766
rect 87676 -138810 87732 -138766
rect 87776 -138810 87832 -138766
rect 87876 -138810 87932 -138766
rect 87976 -138810 88032 -138766
rect 88076 -138810 88132 -138766
rect 88176 -138810 88232 -138766
rect 88276 -138810 88332 -138766
rect 88376 -138810 88432 -138766
rect 88476 -138810 88532 -138766
rect 88576 -138810 88632 -138766
rect 88676 -138810 88732 -138766
rect 88776 -138810 88832 -138766
rect 88876 -138810 88932 -138766
rect 88976 -138810 89032 -138766
rect 89076 -138810 89132 -138766
rect 89176 -138810 89740 -138766
rect 81061 -138866 89740 -138810
rect 81061 -138910 81632 -138866
rect 81676 -138910 81732 -138866
rect 81776 -138910 81832 -138866
rect 81876 -138910 81932 -138866
rect 81976 -138910 82032 -138866
rect 82076 -138910 82132 -138866
rect 82176 -138910 82232 -138866
rect 82276 -138910 82332 -138866
rect 82376 -138910 82432 -138866
rect 82476 -138910 82532 -138866
rect 82576 -138910 82632 -138866
rect 82676 -138910 82732 -138866
rect 82776 -138910 82832 -138866
rect 82876 -138910 82932 -138866
rect 82976 -138910 83032 -138866
rect 83076 -138910 83132 -138866
rect 83176 -138910 83632 -138866
rect 83676 -138910 83732 -138866
rect 83776 -138910 83832 -138866
rect 83876 -138910 83932 -138866
rect 83976 -138910 84032 -138866
rect 84076 -138910 84132 -138866
rect 84176 -138910 84232 -138866
rect 84276 -138910 84332 -138866
rect 84376 -138910 84432 -138866
rect 84476 -138910 84532 -138866
rect 84576 -138910 84632 -138866
rect 84676 -138910 84732 -138866
rect 84776 -138910 84832 -138866
rect 84876 -138910 84932 -138866
rect 84976 -138910 85032 -138866
rect 85076 -138910 85132 -138866
rect 85176 -138910 85632 -138866
rect 85676 -138910 85732 -138866
rect 85776 -138910 85832 -138866
rect 85876 -138910 85932 -138866
rect 85976 -138910 86032 -138866
rect 86076 -138910 86132 -138866
rect 86176 -138910 86232 -138866
rect 86276 -138910 86332 -138866
rect 86376 -138910 86432 -138866
rect 86476 -138910 86532 -138866
rect 86576 -138910 86632 -138866
rect 86676 -138910 86732 -138866
rect 86776 -138910 86832 -138866
rect 86876 -138910 86932 -138866
rect 86976 -138910 87032 -138866
rect 87076 -138910 87132 -138866
rect 87176 -138910 87632 -138866
rect 87676 -138910 87732 -138866
rect 87776 -138910 87832 -138866
rect 87876 -138910 87932 -138866
rect 87976 -138910 88032 -138866
rect 88076 -138910 88132 -138866
rect 88176 -138910 88232 -138866
rect 88276 -138910 88332 -138866
rect 88376 -138910 88432 -138866
rect 88476 -138910 88532 -138866
rect 88576 -138910 88632 -138866
rect 88676 -138910 88732 -138866
rect 88776 -138910 88832 -138866
rect 88876 -138910 88932 -138866
rect 88976 -138910 89032 -138866
rect 89076 -138910 89132 -138866
rect 89176 -138910 89740 -138866
rect 81061 -138966 89740 -138910
rect 81061 -139010 81632 -138966
rect 81676 -139010 81732 -138966
rect 81776 -139010 81832 -138966
rect 81876 -139010 81932 -138966
rect 81976 -139010 82032 -138966
rect 82076 -139010 82132 -138966
rect 82176 -139010 82232 -138966
rect 82276 -139010 82332 -138966
rect 82376 -139010 82432 -138966
rect 82476 -139010 82532 -138966
rect 82576 -139010 82632 -138966
rect 82676 -139010 82732 -138966
rect 82776 -139010 82832 -138966
rect 82876 -139010 82932 -138966
rect 82976 -139010 83032 -138966
rect 83076 -139010 83132 -138966
rect 83176 -139010 83632 -138966
rect 83676 -139010 83732 -138966
rect 83776 -139010 83832 -138966
rect 83876 -139010 83932 -138966
rect 83976 -139010 84032 -138966
rect 84076 -139010 84132 -138966
rect 84176 -139010 84232 -138966
rect 84276 -139010 84332 -138966
rect 84376 -139010 84432 -138966
rect 84476 -139010 84532 -138966
rect 84576 -139010 84632 -138966
rect 84676 -139010 84732 -138966
rect 84776 -139010 84832 -138966
rect 84876 -139010 84932 -138966
rect 84976 -139010 85032 -138966
rect 85076 -139010 85132 -138966
rect 85176 -139010 85632 -138966
rect 85676 -139010 85732 -138966
rect 85776 -139010 85832 -138966
rect 85876 -139010 85932 -138966
rect 85976 -139010 86032 -138966
rect 86076 -139010 86132 -138966
rect 86176 -139010 86232 -138966
rect 86276 -139010 86332 -138966
rect 86376 -139010 86432 -138966
rect 86476 -139010 86532 -138966
rect 86576 -139010 86632 -138966
rect 86676 -139010 86732 -138966
rect 86776 -139010 86832 -138966
rect 86876 -139010 86932 -138966
rect 86976 -139010 87032 -138966
rect 87076 -139010 87132 -138966
rect 87176 -139010 87632 -138966
rect 87676 -139010 87732 -138966
rect 87776 -139010 87832 -138966
rect 87876 -139010 87932 -138966
rect 87976 -139010 88032 -138966
rect 88076 -139010 88132 -138966
rect 88176 -139010 88232 -138966
rect 88276 -139010 88332 -138966
rect 88376 -139010 88432 -138966
rect 88476 -139010 88532 -138966
rect 88576 -139010 88632 -138966
rect 88676 -139010 88732 -138966
rect 88776 -139010 88832 -138966
rect 88876 -139010 88932 -138966
rect 88976 -139010 89032 -138966
rect 89076 -139010 89132 -138966
rect 89176 -139010 89740 -138966
rect 81061 -139066 89740 -139010
rect 81061 -139110 81632 -139066
rect 81676 -139110 81732 -139066
rect 81776 -139110 81832 -139066
rect 81876 -139110 81932 -139066
rect 81976 -139110 82032 -139066
rect 82076 -139110 82132 -139066
rect 82176 -139110 82232 -139066
rect 82276 -139110 82332 -139066
rect 82376 -139110 82432 -139066
rect 82476 -139110 82532 -139066
rect 82576 -139110 82632 -139066
rect 82676 -139110 82732 -139066
rect 82776 -139110 82832 -139066
rect 82876 -139110 82932 -139066
rect 82976 -139110 83032 -139066
rect 83076 -139110 83132 -139066
rect 83176 -139110 83632 -139066
rect 83676 -139110 83732 -139066
rect 83776 -139110 83832 -139066
rect 83876 -139110 83932 -139066
rect 83976 -139110 84032 -139066
rect 84076 -139110 84132 -139066
rect 84176 -139110 84232 -139066
rect 84276 -139110 84332 -139066
rect 84376 -139110 84432 -139066
rect 84476 -139110 84532 -139066
rect 84576 -139110 84632 -139066
rect 84676 -139110 84732 -139066
rect 84776 -139110 84832 -139066
rect 84876 -139110 84932 -139066
rect 84976 -139110 85032 -139066
rect 85076 -139110 85132 -139066
rect 85176 -139110 85632 -139066
rect 85676 -139110 85732 -139066
rect 85776 -139110 85832 -139066
rect 85876 -139110 85932 -139066
rect 85976 -139110 86032 -139066
rect 86076 -139110 86132 -139066
rect 86176 -139110 86232 -139066
rect 86276 -139110 86332 -139066
rect 86376 -139110 86432 -139066
rect 86476 -139110 86532 -139066
rect 86576 -139110 86632 -139066
rect 86676 -139110 86732 -139066
rect 86776 -139110 86832 -139066
rect 86876 -139110 86932 -139066
rect 86976 -139110 87032 -139066
rect 87076 -139110 87132 -139066
rect 87176 -139110 87632 -139066
rect 87676 -139110 87732 -139066
rect 87776 -139110 87832 -139066
rect 87876 -139110 87932 -139066
rect 87976 -139110 88032 -139066
rect 88076 -139110 88132 -139066
rect 88176 -139110 88232 -139066
rect 88276 -139110 88332 -139066
rect 88376 -139110 88432 -139066
rect 88476 -139110 88532 -139066
rect 88576 -139110 88632 -139066
rect 88676 -139110 88732 -139066
rect 88776 -139110 88832 -139066
rect 88876 -139110 88932 -139066
rect 88976 -139110 89032 -139066
rect 89076 -139110 89132 -139066
rect 89176 -139110 89740 -139066
rect 81061 -139166 89740 -139110
rect 81061 -139210 81632 -139166
rect 81676 -139210 81732 -139166
rect 81776 -139210 81832 -139166
rect 81876 -139210 81932 -139166
rect 81976 -139210 82032 -139166
rect 82076 -139210 82132 -139166
rect 82176 -139210 82232 -139166
rect 82276 -139210 82332 -139166
rect 82376 -139210 82432 -139166
rect 82476 -139210 82532 -139166
rect 82576 -139210 82632 -139166
rect 82676 -139210 82732 -139166
rect 82776 -139210 82832 -139166
rect 82876 -139210 82932 -139166
rect 82976 -139210 83032 -139166
rect 83076 -139210 83132 -139166
rect 83176 -139210 83632 -139166
rect 83676 -139210 83732 -139166
rect 83776 -139210 83832 -139166
rect 83876 -139210 83932 -139166
rect 83976 -139210 84032 -139166
rect 84076 -139210 84132 -139166
rect 84176 -139210 84232 -139166
rect 84276 -139210 84332 -139166
rect 84376 -139210 84432 -139166
rect 84476 -139210 84532 -139166
rect 84576 -139210 84632 -139166
rect 84676 -139210 84732 -139166
rect 84776 -139210 84832 -139166
rect 84876 -139210 84932 -139166
rect 84976 -139210 85032 -139166
rect 85076 -139210 85132 -139166
rect 85176 -139210 85632 -139166
rect 85676 -139210 85732 -139166
rect 85776 -139210 85832 -139166
rect 85876 -139210 85932 -139166
rect 85976 -139210 86032 -139166
rect 86076 -139210 86132 -139166
rect 86176 -139210 86232 -139166
rect 86276 -139210 86332 -139166
rect 86376 -139210 86432 -139166
rect 86476 -139210 86532 -139166
rect 86576 -139210 86632 -139166
rect 86676 -139210 86732 -139166
rect 86776 -139210 86832 -139166
rect 86876 -139210 86932 -139166
rect 86976 -139210 87032 -139166
rect 87076 -139210 87132 -139166
rect 87176 -139210 87632 -139166
rect 87676 -139210 87732 -139166
rect 87776 -139210 87832 -139166
rect 87876 -139210 87932 -139166
rect 87976 -139210 88032 -139166
rect 88076 -139210 88132 -139166
rect 88176 -139210 88232 -139166
rect 88276 -139210 88332 -139166
rect 88376 -139210 88432 -139166
rect 88476 -139210 88532 -139166
rect 88576 -139210 88632 -139166
rect 88676 -139210 88732 -139166
rect 88776 -139210 88832 -139166
rect 88876 -139210 88932 -139166
rect 88976 -139210 89032 -139166
rect 89076 -139210 89132 -139166
rect 89176 -139210 89740 -139166
rect 81061 -139266 89740 -139210
rect 81061 -139310 81632 -139266
rect 81676 -139310 81732 -139266
rect 81776 -139310 81832 -139266
rect 81876 -139310 81932 -139266
rect 81976 -139310 82032 -139266
rect 82076 -139310 82132 -139266
rect 82176 -139310 82232 -139266
rect 82276 -139310 82332 -139266
rect 82376 -139310 82432 -139266
rect 82476 -139310 82532 -139266
rect 82576 -139310 82632 -139266
rect 82676 -139310 82732 -139266
rect 82776 -139310 82832 -139266
rect 82876 -139310 82932 -139266
rect 82976 -139310 83032 -139266
rect 83076 -139310 83132 -139266
rect 83176 -139310 83632 -139266
rect 83676 -139310 83732 -139266
rect 83776 -139310 83832 -139266
rect 83876 -139310 83932 -139266
rect 83976 -139310 84032 -139266
rect 84076 -139310 84132 -139266
rect 84176 -139310 84232 -139266
rect 84276 -139310 84332 -139266
rect 84376 -139310 84432 -139266
rect 84476 -139310 84532 -139266
rect 84576 -139310 84632 -139266
rect 84676 -139310 84732 -139266
rect 84776 -139310 84832 -139266
rect 84876 -139310 84932 -139266
rect 84976 -139310 85032 -139266
rect 85076 -139310 85132 -139266
rect 85176 -139310 85632 -139266
rect 85676 -139310 85732 -139266
rect 85776 -139310 85832 -139266
rect 85876 -139310 85932 -139266
rect 85976 -139310 86032 -139266
rect 86076 -139310 86132 -139266
rect 86176 -139310 86232 -139266
rect 86276 -139310 86332 -139266
rect 86376 -139310 86432 -139266
rect 86476 -139310 86532 -139266
rect 86576 -139310 86632 -139266
rect 86676 -139310 86732 -139266
rect 86776 -139310 86832 -139266
rect 86876 -139310 86932 -139266
rect 86976 -139310 87032 -139266
rect 87076 -139310 87132 -139266
rect 87176 -139310 87632 -139266
rect 87676 -139310 87732 -139266
rect 87776 -139310 87832 -139266
rect 87876 -139310 87932 -139266
rect 87976 -139310 88032 -139266
rect 88076 -139310 88132 -139266
rect 88176 -139310 88232 -139266
rect 88276 -139310 88332 -139266
rect 88376 -139310 88432 -139266
rect 88476 -139310 88532 -139266
rect 88576 -139310 88632 -139266
rect 88676 -139310 88732 -139266
rect 88776 -139310 88832 -139266
rect 88876 -139310 88932 -139266
rect 88976 -139310 89032 -139266
rect 89076 -139310 89132 -139266
rect 89176 -139310 89740 -139266
rect 81061 -139366 89740 -139310
rect 81061 -139410 81632 -139366
rect 81676 -139410 81732 -139366
rect 81776 -139410 81832 -139366
rect 81876 -139410 81932 -139366
rect 81976 -139410 82032 -139366
rect 82076 -139410 82132 -139366
rect 82176 -139410 82232 -139366
rect 82276 -139410 82332 -139366
rect 82376 -139410 82432 -139366
rect 82476 -139410 82532 -139366
rect 82576 -139410 82632 -139366
rect 82676 -139410 82732 -139366
rect 82776 -139410 82832 -139366
rect 82876 -139410 82932 -139366
rect 82976 -139410 83032 -139366
rect 83076 -139410 83132 -139366
rect 83176 -139410 83632 -139366
rect 83676 -139410 83732 -139366
rect 83776 -139410 83832 -139366
rect 83876 -139410 83932 -139366
rect 83976 -139410 84032 -139366
rect 84076 -139410 84132 -139366
rect 84176 -139410 84232 -139366
rect 84276 -139410 84332 -139366
rect 84376 -139410 84432 -139366
rect 84476 -139410 84532 -139366
rect 84576 -139410 84632 -139366
rect 84676 -139410 84732 -139366
rect 84776 -139410 84832 -139366
rect 84876 -139410 84932 -139366
rect 84976 -139410 85032 -139366
rect 85076 -139410 85132 -139366
rect 85176 -139410 85632 -139366
rect 85676 -139410 85732 -139366
rect 85776 -139410 85832 -139366
rect 85876 -139410 85932 -139366
rect 85976 -139410 86032 -139366
rect 86076 -139410 86132 -139366
rect 86176 -139410 86232 -139366
rect 86276 -139410 86332 -139366
rect 86376 -139410 86432 -139366
rect 86476 -139410 86532 -139366
rect 86576 -139410 86632 -139366
rect 86676 -139410 86732 -139366
rect 86776 -139410 86832 -139366
rect 86876 -139410 86932 -139366
rect 86976 -139410 87032 -139366
rect 87076 -139410 87132 -139366
rect 87176 -139410 87632 -139366
rect 87676 -139410 87732 -139366
rect 87776 -139410 87832 -139366
rect 87876 -139410 87932 -139366
rect 87976 -139410 88032 -139366
rect 88076 -139410 88132 -139366
rect 88176 -139410 88232 -139366
rect 88276 -139410 88332 -139366
rect 88376 -139410 88432 -139366
rect 88476 -139410 88532 -139366
rect 88576 -139410 88632 -139366
rect 88676 -139410 88732 -139366
rect 88776 -139410 88832 -139366
rect 88876 -139410 88932 -139366
rect 88976 -139410 89032 -139366
rect 89076 -139410 89132 -139366
rect 89176 -139410 89740 -139366
rect 81061 -139466 89740 -139410
rect 81061 -139510 81632 -139466
rect 81676 -139510 81732 -139466
rect 81776 -139510 81832 -139466
rect 81876 -139510 81932 -139466
rect 81976 -139510 82032 -139466
rect 82076 -139510 82132 -139466
rect 82176 -139510 82232 -139466
rect 82276 -139510 82332 -139466
rect 82376 -139510 82432 -139466
rect 82476 -139510 82532 -139466
rect 82576 -139510 82632 -139466
rect 82676 -139510 82732 -139466
rect 82776 -139510 82832 -139466
rect 82876 -139510 82932 -139466
rect 82976 -139510 83032 -139466
rect 83076 -139510 83132 -139466
rect 83176 -139510 83632 -139466
rect 83676 -139510 83732 -139466
rect 83776 -139510 83832 -139466
rect 83876 -139510 83932 -139466
rect 83976 -139510 84032 -139466
rect 84076 -139510 84132 -139466
rect 84176 -139510 84232 -139466
rect 84276 -139510 84332 -139466
rect 84376 -139510 84432 -139466
rect 84476 -139510 84532 -139466
rect 84576 -139510 84632 -139466
rect 84676 -139510 84732 -139466
rect 84776 -139510 84832 -139466
rect 84876 -139510 84932 -139466
rect 84976 -139510 85032 -139466
rect 85076 -139510 85132 -139466
rect 85176 -139510 85632 -139466
rect 85676 -139510 85732 -139466
rect 85776 -139510 85832 -139466
rect 85876 -139510 85932 -139466
rect 85976 -139510 86032 -139466
rect 86076 -139510 86132 -139466
rect 86176 -139510 86232 -139466
rect 86276 -139510 86332 -139466
rect 86376 -139510 86432 -139466
rect 86476 -139510 86532 -139466
rect 86576 -139510 86632 -139466
rect 86676 -139510 86732 -139466
rect 86776 -139510 86832 -139466
rect 86876 -139510 86932 -139466
rect 86976 -139510 87032 -139466
rect 87076 -139510 87132 -139466
rect 87176 -139510 87632 -139466
rect 87676 -139510 87732 -139466
rect 87776 -139510 87832 -139466
rect 87876 -139510 87932 -139466
rect 87976 -139510 88032 -139466
rect 88076 -139510 88132 -139466
rect 88176 -139510 88232 -139466
rect 88276 -139510 88332 -139466
rect 88376 -139510 88432 -139466
rect 88476 -139510 88532 -139466
rect 88576 -139510 88632 -139466
rect 88676 -139510 88732 -139466
rect 88776 -139510 88832 -139466
rect 88876 -139510 88932 -139466
rect 88976 -139510 89032 -139466
rect 89076 -139510 89132 -139466
rect 89176 -139510 89740 -139466
rect 81061 -173049 89740 -139510
rect 142660 -165615 154949 -18989
rect 142660 -165659 145268 -165615
rect 145312 -165659 145368 -165615
rect 145412 -165659 145468 -165615
rect 145512 -165659 145568 -165615
rect 145612 -165659 145668 -165615
rect 145712 -165659 145768 -165615
rect 145812 -165659 145868 -165615
rect 145912 -165659 145968 -165615
rect 146012 -165659 146068 -165615
rect 146112 -165659 146168 -165615
rect 146212 -165659 146268 -165615
rect 146312 -165659 146368 -165615
rect 146412 -165659 146468 -165615
rect 146512 -165659 146568 -165615
rect 146612 -165659 146668 -165615
rect 146712 -165659 146768 -165615
rect 146812 -165659 147268 -165615
rect 147312 -165659 147368 -165615
rect 147412 -165659 147468 -165615
rect 147512 -165659 147568 -165615
rect 147612 -165659 147668 -165615
rect 147712 -165659 147768 -165615
rect 147812 -165659 147868 -165615
rect 147912 -165659 147968 -165615
rect 148012 -165659 148068 -165615
rect 148112 -165659 148168 -165615
rect 148212 -165659 148268 -165615
rect 148312 -165659 148368 -165615
rect 148412 -165659 148468 -165615
rect 148512 -165659 148568 -165615
rect 148612 -165659 148668 -165615
rect 148712 -165659 148768 -165615
rect 148812 -165659 149268 -165615
rect 149312 -165659 149368 -165615
rect 149412 -165659 149468 -165615
rect 149512 -165659 149568 -165615
rect 149612 -165659 149668 -165615
rect 149712 -165659 149768 -165615
rect 149812 -165659 149868 -165615
rect 149912 -165659 149968 -165615
rect 150012 -165659 150068 -165615
rect 150112 -165659 150168 -165615
rect 150212 -165659 150268 -165615
rect 150312 -165659 150368 -165615
rect 150412 -165659 150468 -165615
rect 150512 -165659 150568 -165615
rect 150612 -165659 150668 -165615
rect 150712 -165659 150768 -165615
rect 150812 -165659 151268 -165615
rect 151312 -165659 151368 -165615
rect 151412 -165659 151468 -165615
rect 151512 -165659 151568 -165615
rect 151612 -165659 151668 -165615
rect 151712 -165659 151768 -165615
rect 151812 -165659 151868 -165615
rect 151912 -165659 151968 -165615
rect 152012 -165659 152068 -165615
rect 152112 -165659 152168 -165615
rect 152212 -165659 152268 -165615
rect 152312 -165659 152368 -165615
rect 152412 -165659 152468 -165615
rect 152512 -165659 152568 -165615
rect 152612 -165659 152668 -165615
rect 152712 -165659 152768 -165615
rect 152812 -165659 154949 -165615
rect 142660 -165715 154949 -165659
rect 142660 -165759 145268 -165715
rect 145312 -165759 145368 -165715
rect 145412 -165759 145468 -165715
rect 145512 -165759 145568 -165715
rect 145612 -165759 145668 -165715
rect 145712 -165759 145768 -165715
rect 145812 -165759 145868 -165715
rect 145912 -165759 145968 -165715
rect 146012 -165759 146068 -165715
rect 146112 -165759 146168 -165715
rect 146212 -165759 146268 -165715
rect 146312 -165759 146368 -165715
rect 146412 -165759 146468 -165715
rect 146512 -165759 146568 -165715
rect 146612 -165759 146668 -165715
rect 146712 -165759 146768 -165715
rect 146812 -165759 147268 -165715
rect 147312 -165759 147368 -165715
rect 147412 -165759 147468 -165715
rect 147512 -165759 147568 -165715
rect 147612 -165759 147668 -165715
rect 147712 -165759 147768 -165715
rect 147812 -165759 147868 -165715
rect 147912 -165759 147968 -165715
rect 148012 -165759 148068 -165715
rect 148112 -165759 148168 -165715
rect 148212 -165759 148268 -165715
rect 148312 -165759 148368 -165715
rect 148412 -165759 148468 -165715
rect 148512 -165759 148568 -165715
rect 148612 -165759 148668 -165715
rect 148712 -165759 148768 -165715
rect 148812 -165759 149268 -165715
rect 149312 -165759 149368 -165715
rect 149412 -165759 149468 -165715
rect 149512 -165759 149568 -165715
rect 149612 -165759 149668 -165715
rect 149712 -165759 149768 -165715
rect 149812 -165759 149868 -165715
rect 149912 -165759 149968 -165715
rect 150012 -165759 150068 -165715
rect 150112 -165759 150168 -165715
rect 150212 -165759 150268 -165715
rect 150312 -165759 150368 -165715
rect 150412 -165759 150468 -165715
rect 150512 -165759 150568 -165715
rect 150612 -165759 150668 -165715
rect 150712 -165759 150768 -165715
rect 150812 -165759 151268 -165715
rect 151312 -165759 151368 -165715
rect 151412 -165759 151468 -165715
rect 151512 -165759 151568 -165715
rect 151612 -165759 151668 -165715
rect 151712 -165759 151768 -165715
rect 151812 -165759 151868 -165715
rect 151912 -165759 151968 -165715
rect 152012 -165759 152068 -165715
rect 152112 -165759 152168 -165715
rect 152212 -165759 152268 -165715
rect 152312 -165759 152368 -165715
rect 152412 -165759 152468 -165715
rect 152512 -165759 152568 -165715
rect 152612 -165759 152668 -165715
rect 152712 -165759 152768 -165715
rect 152812 -165759 154949 -165715
rect 142660 -165815 154949 -165759
rect 142660 -165859 145268 -165815
rect 145312 -165859 145368 -165815
rect 145412 -165859 145468 -165815
rect 145512 -165859 145568 -165815
rect 145612 -165859 145668 -165815
rect 145712 -165859 145768 -165815
rect 145812 -165859 145868 -165815
rect 145912 -165859 145968 -165815
rect 146012 -165859 146068 -165815
rect 146112 -165859 146168 -165815
rect 146212 -165859 146268 -165815
rect 146312 -165859 146368 -165815
rect 146412 -165859 146468 -165815
rect 146512 -165859 146568 -165815
rect 146612 -165859 146668 -165815
rect 146712 -165859 146768 -165815
rect 146812 -165859 147268 -165815
rect 147312 -165859 147368 -165815
rect 147412 -165859 147468 -165815
rect 147512 -165859 147568 -165815
rect 147612 -165859 147668 -165815
rect 147712 -165859 147768 -165815
rect 147812 -165859 147868 -165815
rect 147912 -165859 147968 -165815
rect 148012 -165859 148068 -165815
rect 148112 -165859 148168 -165815
rect 148212 -165859 148268 -165815
rect 148312 -165859 148368 -165815
rect 148412 -165859 148468 -165815
rect 148512 -165859 148568 -165815
rect 148612 -165859 148668 -165815
rect 148712 -165859 148768 -165815
rect 148812 -165859 149268 -165815
rect 149312 -165859 149368 -165815
rect 149412 -165859 149468 -165815
rect 149512 -165859 149568 -165815
rect 149612 -165859 149668 -165815
rect 149712 -165859 149768 -165815
rect 149812 -165859 149868 -165815
rect 149912 -165859 149968 -165815
rect 150012 -165859 150068 -165815
rect 150112 -165859 150168 -165815
rect 150212 -165859 150268 -165815
rect 150312 -165859 150368 -165815
rect 150412 -165859 150468 -165815
rect 150512 -165859 150568 -165815
rect 150612 -165859 150668 -165815
rect 150712 -165859 150768 -165815
rect 150812 -165859 151268 -165815
rect 151312 -165859 151368 -165815
rect 151412 -165859 151468 -165815
rect 151512 -165859 151568 -165815
rect 151612 -165859 151668 -165815
rect 151712 -165859 151768 -165815
rect 151812 -165859 151868 -165815
rect 151912 -165859 151968 -165815
rect 152012 -165859 152068 -165815
rect 152112 -165859 152168 -165815
rect 152212 -165859 152268 -165815
rect 152312 -165859 152368 -165815
rect 152412 -165859 152468 -165815
rect 152512 -165859 152568 -165815
rect 152612 -165859 152668 -165815
rect 152712 -165859 152768 -165815
rect 152812 -165859 154949 -165815
rect 142660 -165915 154949 -165859
rect 142660 -165959 145268 -165915
rect 145312 -165959 145368 -165915
rect 145412 -165959 145468 -165915
rect 145512 -165959 145568 -165915
rect 145612 -165959 145668 -165915
rect 145712 -165959 145768 -165915
rect 145812 -165959 145868 -165915
rect 145912 -165959 145968 -165915
rect 146012 -165959 146068 -165915
rect 146112 -165959 146168 -165915
rect 146212 -165959 146268 -165915
rect 146312 -165959 146368 -165915
rect 146412 -165959 146468 -165915
rect 146512 -165959 146568 -165915
rect 146612 -165959 146668 -165915
rect 146712 -165959 146768 -165915
rect 146812 -165959 147268 -165915
rect 147312 -165959 147368 -165915
rect 147412 -165959 147468 -165915
rect 147512 -165959 147568 -165915
rect 147612 -165959 147668 -165915
rect 147712 -165959 147768 -165915
rect 147812 -165959 147868 -165915
rect 147912 -165959 147968 -165915
rect 148012 -165959 148068 -165915
rect 148112 -165959 148168 -165915
rect 148212 -165959 148268 -165915
rect 148312 -165959 148368 -165915
rect 148412 -165959 148468 -165915
rect 148512 -165959 148568 -165915
rect 148612 -165959 148668 -165915
rect 148712 -165959 148768 -165915
rect 148812 -165959 149268 -165915
rect 149312 -165959 149368 -165915
rect 149412 -165959 149468 -165915
rect 149512 -165959 149568 -165915
rect 149612 -165959 149668 -165915
rect 149712 -165959 149768 -165915
rect 149812 -165959 149868 -165915
rect 149912 -165959 149968 -165915
rect 150012 -165959 150068 -165915
rect 150112 -165959 150168 -165915
rect 150212 -165959 150268 -165915
rect 150312 -165959 150368 -165915
rect 150412 -165959 150468 -165915
rect 150512 -165959 150568 -165915
rect 150612 -165959 150668 -165915
rect 150712 -165959 150768 -165915
rect 150812 -165959 151268 -165915
rect 151312 -165959 151368 -165915
rect 151412 -165959 151468 -165915
rect 151512 -165959 151568 -165915
rect 151612 -165959 151668 -165915
rect 151712 -165959 151768 -165915
rect 151812 -165959 151868 -165915
rect 151912 -165959 151968 -165915
rect 152012 -165959 152068 -165915
rect 152112 -165959 152168 -165915
rect 152212 -165959 152268 -165915
rect 152312 -165959 152368 -165915
rect 152412 -165959 152468 -165915
rect 152512 -165959 152568 -165915
rect 152612 -165959 152668 -165915
rect 152712 -165959 152768 -165915
rect 152812 -165959 154949 -165915
rect 142660 -166015 154949 -165959
rect 142660 -166059 145268 -166015
rect 145312 -166059 145368 -166015
rect 145412 -166059 145468 -166015
rect 145512 -166059 145568 -166015
rect 145612 -166059 145668 -166015
rect 145712 -166059 145768 -166015
rect 145812 -166059 145868 -166015
rect 145912 -166059 145968 -166015
rect 146012 -166059 146068 -166015
rect 146112 -166059 146168 -166015
rect 146212 -166059 146268 -166015
rect 146312 -166059 146368 -166015
rect 146412 -166059 146468 -166015
rect 146512 -166059 146568 -166015
rect 146612 -166059 146668 -166015
rect 146712 -166059 146768 -166015
rect 146812 -166059 147268 -166015
rect 147312 -166059 147368 -166015
rect 147412 -166059 147468 -166015
rect 147512 -166059 147568 -166015
rect 147612 -166059 147668 -166015
rect 147712 -166059 147768 -166015
rect 147812 -166059 147868 -166015
rect 147912 -166059 147968 -166015
rect 148012 -166059 148068 -166015
rect 148112 -166059 148168 -166015
rect 148212 -166059 148268 -166015
rect 148312 -166059 148368 -166015
rect 148412 -166059 148468 -166015
rect 148512 -166059 148568 -166015
rect 148612 -166059 148668 -166015
rect 148712 -166059 148768 -166015
rect 148812 -166059 149268 -166015
rect 149312 -166059 149368 -166015
rect 149412 -166059 149468 -166015
rect 149512 -166059 149568 -166015
rect 149612 -166059 149668 -166015
rect 149712 -166059 149768 -166015
rect 149812 -166059 149868 -166015
rect 149912 -166059 149968 -166015
rect 150012 -166059 150068 -166015
rect 150112 -166059 150168 -166015
rect 150212 -166059 150268 -166015
rect 150312 -166059 150368 -166015
rect 150412 -166059 150468 -166015
rect 150512 -166059 150568 -166015
rect 150612 -166059 150668 -166015
rect 150712 -166059 150768 -166015
rect 150812 -166059 151268 -166015
rect 151312 -166059 151368 -166015
rect 151412 -166059 151468 -166015
rect 151512 -166059 151568 -166015
rect 151612 -166059 151668 -166015
rect 151712 -166059 151768 -166015
rect 151812 -166059 151868 -166015
rect 151912 -166059 151968 -166015
rect 152012 -166059 152068 -166015
rect 152112 -166059 152168 -166015
rect 152212 -166059 152268 -166015
rect 152312 -166059 152368 -166015
rect 152412 -166059 152468 -166015
rect 152512 -166059 152568 -166015
rect 152612 -166059 152668 -166015
rect 152712 -166059 152768 -166015
rect 152812 -166059 154949 -166015
rect 142660 -166115 154949 -166059
rect 142660 -166159 145268 -166115
rect 145312 -166159 145368 -166115
rect 145412 -166159 145468 -166115
rect 145512 -166159 145568 -166115
rect 145612 -166159 145668 -166115
rect 145712 -166159 145768 -166115
rect 145812 -166159 145868 -166115
rect 145912 -166159 145968 -166115
rect 146012 -166159 146068 -166115
rect 146112 -166159 146168 -166115
rect 146212 -166159 146268 -166115
rect 146312 -166159 146368 -166115
rect 146412 -166159 146468 -166115
rect 146512 -166159 146568 -166115
rect 146612 -166159 146668 -166115
rect 146712 -166159 146768 -166115
rect 146812 -166159 147268 -166115
rect 147312 -166159 147368 -166115
rect 147412 -166159 147468 -166115
rect 147512 -166159 147568 -166115
rect 147612 -166159 147668 -166115
rect 147712 -166159 147768 -166115
rect 147812 -166159 147868 -166115
rect 147912 -166159 147968 -166115
rect 148012 -166159 148068 -166115
rect 148112 -166159 148168 -166115
rect 148212 -166159 148268 -166115
rect 148312 -166159 148368 -166115
rect 148412 -166159 148468 -166115
rect 148512 -166159 148568 -166115
rect 148612 -166159 148668 -166115
rect 148712 -166159 148768 -166115
rect 148812 -166159 149268 -166115
rect 149312 -166159 149368 -166115
rect 149412 -166159 149468 -166115
rect 149512 -166159 149568 -166115
rect 149612 -166159 149668 -166115
rect 149712 -166159 149768 -166115
rect 149812 -166159 149868 -166115
rect 149912 -166159 149968 -166115
rect 150012 -166159 150068 -166115
rect 150112 -166159 150168 -166115
rect 150212 -166159 150268 -166115
rect 150312 -166159 150368 -166115
rect 150412 -166159 150468 -166115
rect 150512 -166159 150568 -166115
rect 150612 -166159 150668 -166115
rect 150712 -166159 150768 -166115
rect 150812 -166159 151268 -166115
rect 151312 -166159 151368 -166115
rect 151412 -166159 151468 -166115
rect 151512 -166159 151568 -166115
rect 151612 -166159 151668 -166115
rect 151712 -166159 151768 -166115
rect 151812 -166159 151868 -166115
rect 151912 -166159 151968 -166115
rect 152012 -166159 152068 -166115
rect 152112 -166159 152168 -166115
rect 152212 -166159 152268 -166115
rect 152312 -166159 152368 -166115
rect 152412 -166159 152468 -166115
rect 152512 -166159 152568 -166115
rect 152612 -166159 152668 -166115
rect 152712 -166159 152768 -166115
rect 152812 -166159 154949 -166115
rect 142660 -166215 154949 -166159
rect 142660 -166259 145268 -166215
rect 145312 -166259 145368 -166215
rect 145412 -166259 145468 -166215
rect 145512 -166259 145568 -166215
rect 145612 -166259 145668 -166215
rect 145712 -166259 145768 -166215
rect 145812 -166259 145868 -166215
rect 145912 -166259 145968 -166215
rect 146012 -166259 146068 -166215
rect 146112 -166259 146168 -166215
rect 146212 -166259 146268 -166215
rect 146312 -166259 146368 -166215
rect 146412 -166259 146468 -166215
rect 146512 -166259 146568 -166215
rect 146612 -166259 146668 -166215
rect 146712 -166259 146768 -166215
rect 146812 -166259 147268 -166215
rect 147312 -166259 147368 -166215
rect 147412 -166259 147468 -166215
rect 147512 -166259 147568 -166215
rect 147612 -166259 147668 -166215
rect 147712 -166259 147768 -166215
rect 147812 -166259 147868 -166215
rect 147912 -166259 147968 -166215
rect 148012 -166259 148068 -166215
rect 148112 -166259 148168 -166215
rect 148212 -166259 148268 -166215
rect 148312 -166259 148368 -166215
rect 148412 -166259 148468 -166215
rect 148512 -166259 148568 -166215
rect 148612 -166259 148668 -166215
rect 148712 -166259 148768 -166215
rect 148812 -166259 149268 -166215
rect 149312 -166259 149368 -166215
rect 149412 -166259 149468 -166215
rect 149512 -166259 149568 -166215
rect 149612 -166259 149668 -166215
rect 149712 -166259 149768 -166215
rect 149812 -166259 149868 -166215
rect 149912 -166259 149968 -166215
rect 150012 -166259 150068 -166215
rect 150112 -166259 150168 -166215
rect 150212 -166259 150268 -166215
rect 150312 -166259 150368 -166215
rect 150412 -166259 150468 -166215
rect 150512 -166259 150568 -166215
rect 150612 -166259 150668 -166215
rect 150712 -166259 150768 -166215
rect 150812 -166259 151268 -166215
rect 151312 -166259 151368 -166215
rect 151412 -166259 151468 -166215
rect 151512 -166259 151568 -166215
rect 151612 -166259 151668 -166215
rect 151712 -166259 151768 -166215
rect 151812 -166259 151868 -166215
rect 151912 -166259 151968 -166215
rect 152012 -166259 152068 -166215
rect 152112 -166259 152168 -166215
rect 152212 -166259 152268 -166215
rect 152312 -166259 152368 -166215
rect 152412 -166259 152468 -166215
rect 152512 -166259 152568 -166215
rect 152612 -166259 152668 -166215
rect 152712 -166259 152768 -166215
rect 152812 -166259 154949 -166215
rect 142660 -166315 154949 -166259
rect 142660 -166359 145268 -166315
rect 145312 -166359 145368 -166315
rect 145412 -166359 145468 -166315
rect 145512 -166359 145568 -166315
rect 145612 -166359 145668 -166315
rect 145712 -166359 145768 -166315
rect 145812 -166359 145868 -166315
rect 145912 -166359 145968 -166315
rect 146012 -166359 146068 -166315
rect 146112 -166359 146168 -166315
rect 146212 -166359 146268 -166315
rect 146312 -166359 146368 -166315
rect 146412 -166359 146468 -166315
rect 146512 -166359 146568 -166315
rect 146612 -166359 146668 -166315
rect 146712 -166359 146768 -166315
rect 146812 -166359 147268 -166315
rect 147312 -166359 147368 -166315
rect 147412 -166359 147468 -166315
rect 147512 -166359 147568 -166315
rect 147612 -166359 147668 -166315
rect 147712 -166359 147768 -166315
rect 147812 -166359 147868 -166315
rect 147912 -166359 147968 -166315
rect 148012 -166359 148068 -166315
rect 148112 -166359 148168 -166315
rect 148212 -166359 148268 -166315
rect 148312 -166359 148368 -166315
rect 148412 -166359 148468 -166315
rect 148512 -166359 148568 -166315
rect 148612 -166359 148668 -166315
rect 148712 -166359 148768 -166315
rect 148812 -166359 149268 -166315
rect 149312 -166359 149368 -166315
rect 149412 -166359 149468 -166315
rect 149512 -166359 149568 -166315
rect 149612 -166359 149668 -166315
rect 149712 -166359 149768 -166315
rect 149812 -166359 149868 -166315
rect 149912 -166359 149968 -166315
rect 150012 -166359 150068 -166315
rect 150112 -166359 150168 -166315
rect 150212 -166359 150268 -166315
rect 150312 -166359 150368 -166315
rect 150412 -166359 150468 -166315
rect 150512 -166359 150568 -166315
rect 150612 -166359 150668 -166315
rect 150712 -166359 150768 -166315
rect 150812 -166359 151268 -166315
rect 151312 -166359 151368 -166315
rect 151412 -166359 151468 -166315
rect 151512 -166359 151568 -166315
rect 151612 -166359 151668 -166315
rect 151712 -166359 151768 -166315
rect 151812 -166359 151868 -166315
rect 151912 -166359 151968 -166315
rect 152012 -166359 152068 -166315
rect 152112 -166359 152168 -166315
rect 152212 -166359 152268 -166315
rect 152312 -166359 152368 -166315
rect 152412 -166359 152468 -166315
rect 152512 -166359 152568 -166315
rect 152612 -166359 152668 -166315
rect 152712 -166359 152768 -166315
rect 152812 -166359 154949 -166315
rect 142660 -166415 154949 -166359
rect 142660 -166459 145268 -166415
rect 145312 -166459 145368 -166415
rect 145412 -166459 145468 -166415
rect 145512 -166459 145568 -166415
rect 145612 -166459 145668 -166415
rect 145712 -166459 145768 -166415
rect 145812 -166459 145868 -166415
rect 145912 -166459 145968 -166415
rect 146012 -166459 146068 -166415
rect 146112 -166459 146168 -166415
rect 146212 -166459 146268 -166415
rect 146312 -166459 146368 -166415
rect 146412 -166459 146468 -166415
rect 146512 -166459 146568 -166415
rect 146612 -166459 146668 -166415
rect 146712 -166459 146768 -166415
rect 146812 -166459 147268 -166415
rect 147312 -166459 147368 -166415
rect 147412 -166459 147468 -166415
rect 147512 -166459 147568 -166415
rect 147612 -166459 147668 -166415
rect 147712 -166459 147768 -166415
rect 147812 -166459 147868 -166415
rect 147912 -166459 147968 -166415
rect 148012 -166459 148068 -166415
rect 148112 -166459 148168 -166415
rect 148212 -166459 148268 -166415
rect 148312 -166459 148368 -166415
rect 148412 -166459 148468 -166415
rect 148512 -166459 148568 -166415
rect 148612 -166459 148668 -166415
rect 148712 -166459 148768 -166415
rect 148812 -166459 149268 -166415
rect 149312 -166459 149368 -166415
rect 149412 -166459 149468 -166415
rect 149512 -166459 149568 -166415
rect 149612 -166459 149668 -166415
rect 149712 -166459 149768 -166415
rect 149812 -166459 149868 -166415
rect 149912 -166459 149968 -166415
rect 150012 -166459 150068 -166415
rect 150112 -166459 150168 -166415
rect 150212 -166459 150268 -166415
rect 150312 -166459 150368 -166415
rect 150412 -166459 150468 -166415
rect 150512 -166459 150568 -166415
rect 150612 -166459 150668 -166415
rect 150712 -166459 150768 -166415
rect 150812 -166459 151268 -166415
rect 151312 -166459 151368 -166415
rect 151412 -166459 151468 -166415
rect 151512 -166459 151568 -166415
rect 151612 -166459 151668 -166415
rect 151712 -166459 151768 -166415
rect 151812 -166459 151868 -166415
rect 151912 -166459 151968 -166415
rect 152012 -166459 152068 -166415
rect 152112 -166459 152168 -166415
rect 152212 -166459 152268 -166415
rect 152312 -166459 152368 -166415
rect 152412 -166459 152468 -166415
rect 152512 -166459 152568 -166415
rect 152612 -166459 152668 -166415
rect 152712 -166459 152768 -166415
rect 152812 -166459 154949 -166415
rect 142660 -166515 154949 -166459
rect 142660 -166559 145268 -166515
rect 145312 -166559 145368 -166515
rect 145412 -166559 145468 -166515
rect 145512 -166559 145568 -166515
rect 145612 -166559 145668 -166515
rect 145712 -166559 145768 -166515
rect 145812 -166559 145868 -166515
rect 145912 -166559 145968 -166515
rect 146012 -166559 146068 -166515
rect 146112 -166559 146168 -166515
rect 146212 -166559 146268 -166515
rect 146312 -166559 146368 -166515
rect 146412 -166559 146468 -166515
rect 146512 -166559 146568 -166515
rect 146612 -166559 146668 -166515
rect 146712 -166559 146768 -166515
rect 146812 -166559 147268 -166515
rect 147312 -166559 147368 -166515
rect 147412 -166559 147468 -166515
rect 147512 -166559 147568 -166515
rect 147612 -166559 147668 -166515
rect 147712 -166559 147768 -166515
rect 147812 -166559 147868 -166515
rect 147912 -166559 147968 -166515
rect 148012 -166559 148068 -166515
rect 148112 -166559 148168 -166515
rect 148212 -166559 148268 -166515
rect 148312 -166559 148368 -166515
rect 148412 -166559 148468 -166515
rect 148512 -166559 148568 -166515
rect 148612 -166559 148668 -166515
rect 148712 -166559 148768 -166515
rect 148812 -166559 149268 -166515
rect 149312 -166559 149368 -166515
rect 149412 -166559 149468 -166515
rect 149512 -166559 149568 -166515
rect 149612 -166559 149668 -166515
rect 149712 -166559 149768 -166515
rect 149812 -166559 149868 -166515
rect 149912 -166559 149968 -166515
rect 150012 -166559 150068 -166515
rect 150112 -166559 150168 -166515
rect 150212 -166559 150268 -166515
rect 150312 -166559 150368 -166515
rect 150412 -166559 150468 -166515
rect 150512 -166559 150568 -166515
rect 150612 -166559 150668 -166515
rect 150712 -166559 150768 -166515
rect 150812 -166559 151268 -166515
rect 151312 -166559 151368 -166515
rect 151412 -166559 151468 -166515
rect 151512 -166559 151568 -166515
rect 151612 -166559 151668 -166515
rect 151712 -166559 151768 -166515
rect 151812 -166559 151868 -166515
rect 151912 -166559 151968 -166515
rect 152012 -166559 152068 -166515
rect 152112 -166559 152168 -166515
rect 152212 -166559 152268 -166515
rect 152312 -166559 152368 -166515
rect 152412 -166559 152468 -166515
rect 152512 -166559 152568 -166515
rect 152612 -166559 152668 -166515
rect 152712 -166559 152768 -166515
rect 152812 -166559 154949 -166515
rect 142660 -166615 154949 -166559
rect 142660 -166659 145268 -166615
rect 145312 -166659 145368 -166615
rect 145412 -166659 145468 -166615
rect 145512 -166659 145568 -166615
rect 145612 -166659 145668 -166615
rect 145712 -166659 145768 -166615
rect 145812 -166659 145868 -166615
rect 145912 -166659 145968 -166615
rect 146012 -166659 146068 -166615
rect 146112 -166659 146168 -166615
rect 146212 -166659 146268 -166615
rect 146312 -166659 146368 -166615
rect 146412 -166659 146468 -166615
rect 146512 -166659 146568 -166615
rect 146612 -166659 146668 -166615
rect 146712 -166659 146768 -166615
rect 146812 -166659 147268 -166615
rect 147312 -166659 147368 -166615
rect 147412 -166659 147468 -166615
rect 147512 -166659 147568 -166615
rect 147612 -166659 147668 -166615
rect 147712 -166659 147768 -166615
rect 147812 -166659 147868 -166615
rect 147912 -166659 147968 -166615
rect 148012 -166659 148068 -166615
rect 148112 -166659 148168 -166615
rect 148212 -166659 148268 -166615
rect 148312 -166659 148368 -166615
rect 148412 -166659 148468 -166615
rect 148512 -166659 148568 -166615
rect 148612 -166659 148668 -166615
rect 148712 -166659 148768 -166615
rect 148812 -166659 149268 -166615
rect 149312 -166659 149368 -166615
rect 149412 -166659 149468 -166615
rect 149512 -166659 149568 -166615
rect 149612 -166659 149668 -166615
rect 149712 -166659 149768 -166615
rect 149812 -166659 149868 -166615
rect 149912 -166659 149968 -166615
rect 150012 -166659 150068 -166615
rect 150112 -166659 150168 -166615
rect 150212 -166659 150268 -166615
rect 150312 -166659 150368 -166615
rect 150412 -166659 150468 -166615
rect 150512 -166659 150568 -166615
rect 150612 -166659 150668 -166615
rect 150712 -166659 150768 -166615
rect 150812 -166659 151268 -166615
rect 151312 -166659 151368 -166615
rect 151412 -166659 151468 -166615
rect 151512 -166659 151568 -166615
rect 151612 -166659 151668 -166615
rect 151712 -166659 151768 -166615
rect 151812 -166659 151868 -166615
rect 151912 -166659 151968 -166615
rect 152012 -166659 152068 -166615
rect 152112 -166659 152168 -166615
rect 152212 -166659 152268 -166615
rect 152312 -166659 152368 -166615
rect 152412 -166659 152468 -166615
rect 152512 -166659 152568 -166615
rect 152612 -166659 152668 -166615
rect 152712 -166659 152768 -166615
rect 152812 -166659 154949 -166615
rect 142660 -166715 154949 -166659
rect 142660 -166759 145268 -166715
rect 145312 -166759 145368 -166715
rect 145412 -166759 145468 -166715
rect 145512 -166759 145568 -166715
rect 145612 -166759 145668 -166715
rect 145712 -166759 145768 -166715
rect 145812 -166759 145868 -166715
rect 145912 -166759 145968 -166715
rect 146012 -166759 146068 -166715
rect 146112 -166759 146168 -166715
rect 146212 -166759 146268 -166715
rect 146312 -166759 146368 -166715
rect 146412 -166759 146468 -166715
rect 146512 -166759 146568 -166715
rect 146612 -166759 146668 -166715
rect 146712 -166759 146768 -166715
rect 146812 -166759 147268 -166715
rect 147312 -166759 147368 -166715
rect 147412 -166759 147468 -166715
rect 147512 -166759 147568 -166715
rect 147612 -166759 147668 -166715
rect 147712 -166759 147768 -166715
rect 147812 -166759 147868 -166715
rect 147912 -166759 147968 -166715
rect 148012 -166759 148068 -166715
rect 148112 -166759 148168 -166715
rect 148212 -166759 148268 -166715
rect 148312 -166759 148368 -166715
rect 148412 -166759 148468 -166715
rect 148512 -166759 148568 -166715
rect 148612 -166759 148668 -166715
rect 148712 -166759 148768 -166715
rect 148812 -166759 149268 -166715
rect 149312 -166759 149368 -166715
rect 149412 -166759 149468 -166715
rect 149512 -166759 149568 -166715
rect 149612 -166759 149668 -166715
rect 149712 -166759 149768 -166715
rect 149812 -166759 149868 -166715
rect 149912 -166759 149968 -166715
rect 150012 -166759 150068 -166715
rect 150112 -166759 150168 -166715
rect 150212 -166759 150268 -166715
rect 150312 -166759 150368 -166715
rect 150412 -166759 150468 -166715
rect 150512 -166759 150568 -166715
rect 150612 -166759 150668 -166715
rect 150712 -166759 150768 -166715
rect 150812 -166759 151268 -166715
rect 151312 -166759 151368 -166715
rect 151412 -166759 151468 -166715
rect 151512 -166759 151568 -166715
rect 151612 -166759 151668 -166715
rect 151712 -166759 151768 -166715
rect 151812 -166759 151868 -166715
rect 151912 -166759 151968 -166715
rect 152012 -166759 152068 -166715
rect 152112 -166759 152168 -166715
rect 152212 -166759 152268 -166715
rect 152312 -166759 152368 -166715
rect 152412 -166759 152468 -166715
rect 152512 -166759 152568 -166715
rect 152612 -166759 152668 -166715
rect 152712 -166759 152768 -166715
rect 152812 -166759 154949 -166715
rect 142660 -166815 154949 -166759
rect 142660 -166859 145268 -166815
rect 145312 -166859 145368 -166815
rect 145412 -166859 145468 -166815
rect 145512 -166859 145568 -166815
rect 145612 -166859 145668 -166815
rect 145712 -166859 145768 -166815
rect 145812 -166859 145868 -166815
rect 145912 -166859 145968 -166815
rect 146012 -166859 146068 -166815
rect 146112 -166859 146168 -166815
rect 146212 -166859 146268 -166815
rect 146312 -166859 146368 -166815
rect 146412 -166859 146468 -166815
rect 146512 -166859 146568 -166815
rect 146612 -166859 146668 -166815
rect 146712 -166859 146768 -166815
rect 146812 -166859 147268 -166815
rect 147312 -166859 147368 -166815
rect 147412 -166859 147468 -166815
rect 147512 -166859 147568 -166815
rect 147612 -166859 147668 -166815
rect 147712 -166859 147768 -166815
rect 147812 -166859 147868 -166815
rect 147912 -166859 147968 -166815
rect 148012 -166859 148068 -166815
rect 148112 -166859 148168 -166815
rect 148212 -166859 148268 -166815
rect 148312 -166859 148368 -166815
rect 148412 -166859 148468 -166815
rect 148512 -166859 148568 -166815
rect 148612 -166859 148668 -166815
rect 148712 -166859 148768 -166815
rect 148812 -166859 149268 -166815
rect 149312 -166859 149368 -166815
rect 149412 -166859 149468 -166815
rect 149512 -166859 149568 -166815
rect 149612 -166859 149668 -166815
rect 149712 -166859 149768 -166815
rect 149812 -166859 149868 -166815
rect 149912 -166859 149968 -166815
rect 150012 -166859 150068 -166815
rect 150112 -166859 150168 -166815
rect 150212 -166859 150268 -166815
rect 150312 -166859 150368 -166815
rect 150412 -166859 150468 -166815
rect 150512 -166859 150568 -166815
rect 150612 -166859 150668 -166815
rect 150712 -166859 150768 -166815
rect 150812 -166859 151268 -166815
rect 151312 -166859 151368 -166815
rect 151412 -166859 151468 -166815
rect 151512 -166859 151568 -166815
rect 151612 -166859 151668 -166815
rect 151712 -166859 151768 -166815
rect 151812 -166859 151868 -166815
rect 151912 -166859 151968 -166815
rect 152012 -166859 152068 -166815
rect 152112 -166859 152168 -166815
rect 152212 -166859 152268 -166815
rect 152312 -166859 152368 -166815
rect 152412 -166859 152468 -166815
rect 152512 -166859 152568 -166815
rect 152612 -166859 152668 -166815
rect 152712 -166859 152768 -166815
rect 152812 -166859 154949 -166815
rect 142660 -166915 154949 -166859
rect 142660 -166959 145268 -166915
rect 145312 -166959 145368 -166915
rect 145412 -166959 145468 -166915
rect 145512 -166959 145568 -166915
rect 145612 -166959 145668 -166915
rect 145712 -166959 145768 -166915
rect 145812 -166959 145868 -166915
rect 145912 -166959 145968 -166915
rect 146012 -166959 146068 -166915
rect 146112 -166959 146168 -166915
rect 146212 -166959 146268 -166915
rect 146312 -166959 146368 -166915
rect 146412 -166959 146468 -166915
rect 146512 -166959 146568 -166915
rect 146612 -166959 146668 -166915
rect 146712 -166959 146768 -166915
rect 146812 -166959 147268 -166915
rect 147312 -166959 147368 -166915
rect 147412 -166959 147468 -166915
rect 147512 -166959 147568 -166915
rect 147612 -166959 147668 -166915
rect 147712 -166959 147768 -166915
rect 147812 -166959 147868 -166915
rect 147912 -166959 147968 -166915
rect 148012 -166959 148068 -166915
rect 148112 -166959 148168 -166915
rect 148212 -166959 148268 -166915
rect 148312 -166959 148368 -166915
rect 148412 -166959 148468 -166915
rect 148512 -166959 148568 -166915
rect 148612 -166959 148668 -166915
rect 148712 -166959 148768 -166915
rect 148812 -166959 149268 -166915
rect 149312 -166959 149368 -166915
rect 149412 -166959 149468 -166915
rect 149512 -166959 149568 -166915
rect 149612 -166959 149668 -166915
rect 149712 -166959 149768 -166915
rect 149812 -166959 149868 -166915
rect 149912 -166959 149968 -166915
rect 150012 -166959 150068 -166915
rect 150112 -166959 150168 -166915
rect 150212 -166959 150268 -166915
rect 150312 -166959 150368 -166915
rect 150412 -166959 150468 -166915
rect 150512 -166959 150568 -166915
rect 150612 -166959 150668 -166915
rect 150712 -166959 150768 -166915
rect 150812 -166959 151268 -166915
rect 151312 -166959 151368 -166915
rect 151412 -166959 151468 -166915
rect 151512 -166959 151568 -166915
rect 151612 -166959 151668 -166915
rect 151712 -166959 151768 -166915
rect 151812 -166959 151868 -166915
rect 151912 -166959 151968 -166915
rect 152012 -166959 152068 -166915
rect 152112 -166959 152168 -166915
rect 152212 -166959 152268 -166915
rect 152312 -166959 152368 -166915
rect 152412 -166959 152468 -166915
rect 152512 -166959 152568 -166915
rect 152612 -166959 152668 -166915
rect 152712 -166959 152768 -166915
rect 152812 -166959 154949 -166915
rect 142660 -167015 154949 -166959
rect 142660 -167059 145268 -167015
rect 145312 -167059 145368 -167015
rect 145412 -167059 145468 -167015
rect 145512 -167059 145568 -167015
rect 145612 -167059 145668 -167015
rect 145712 -167059 145768 -167015
rect 145812 -167059 145868 -167015
rect 145912 -167059 145968 -167015
rect 146012 -167059 146068 -167015
rect 146112 -167059 146168 -167015
rect 146212 -167059 146268 -167015
rect 146312 -167059 146368 -167015
rect 146412 -167059 146468 -167015
rect 146512 -167059 146568 -167015
rect 146612 -167059 146668 -167015
rect 146712 -167059 146768 -167015
rect 146812 -167059 147268 -167015
rect 147312 -167059 147368 -167015
rect 147412 -167059 147468 -167015
rect 147512 -167059 147568 -167015
rect 147612 -167059 147668 -167015
rect 147712 -167059 147768 -167015
rect 147812 -167059 147868 -167015
rect 147912 -167059 147968 -167015
rect 148012 -167059 148068 -167015
rect 148112 -167059 148168 -167015
rect 148212 -167059 148268 -167015
rect 148312 -167059 148368 -167015
rect 148412 -167059 148468 -167015
rect 148512 -167059 148568 -167015
rect 148612 -167059 148668 -167015
rect 148712 -167059 148768 -167015
rect 148812 -167059 149268 -167015
rect 149312 -167059 149368 -167015
rect 149412 -167059 149468 -167015
rect 149512 -167059 149568 -167015
rect 149612 -167059 149668 -167015
rect 149712 -167059 149768 -167015
rect 149812 -167059 149868 -167015
rect 149912 -167059 149968 -167015
rect 150012 -167059 150068 -167015
rect 150112 -167059 150168 -167015
rect 150212 -167059 150268 -167015
rect 150312 -167059 150368 -167015
rect 150412 -167059 150468 -167015
rect 150512 -167059 150568 -167015
rect 150612 -167059 150668 -167015
rect 150712 -167059 150768 -167015
rect 150812 -167059 151268 -167015
rect 151312 -167059 151368 -167015
rect 151412 -167059 151468 -167015
rect 151512 -167059 151568 -167015
rect 151612 -167059 151668 -167015
rect 151712 -167059 151768 -167015
rect 151812 -167059 151868 -167015
rect 151912 -167059 151968 -167015
rect 152012 -167059 152068 -167015
rect 152112 -167059 152168 -167015
rect 152212 -167059 152268 -167015
rect 152312 -167059 152368 -167015
rect 152412 -167059 152468 -167015
rect 152512 -167059 152568 -167015
rect 152612 -167059 152668 -167015
rect 152712 -167059 152768 -167015
rect 152812 -167059 154949 -167015
rect 142660 -167115 154949 -167059
rect 142660 -167159 145268 -167115
rect 145312 -167159 145368 -167115
rect 145412 -167159 145468 -167115
rect 145512 -167159 145568 -167115
rect 145612 -167159 145668 -167115
rect 145712 -167159 145768 -167115
rect 145812 -167159 145868 -167115
rect 145912 -167159 145968 -167115
rect 146012 -167159 146068 -167115
rect 146112 -167159 146168 -167115
rect 146212 -167159 146268 -167115
rect 146312 -167159 146368 -167115
rect 146412 -167159 146468 -167115
rect 146512 -167159 146568 -167115
rect 146612 -167159 146668 -167115
rect 146712 -167159 146768 -167115
rect 146812 -167159 147268 -167115
rect 147312 -167159 147368 -167115
rect 147412 -167159 147468 -167115
rect 147512 -167159 147568 -167115
rect 147612 -167159 147668 -167115
rect 147712 -167159 147768 -167115
rect 147812 -167159 147868 -167115
rect 147912 -167159 147968 -167115
rect 148012 -167159 148068 -167115
rect 148112 -167159 148168 -167115
rect 148212 -167159 148268 -167115
rect 148312 -167159 148368 -167115
rect 148412 -167159 148468 -167115
rect 148512 -167159 148568 -167115
rect 148612 -167159 148668 -167115
rect 148712 -167159 148768 -167115
rect 148812 -167159 149268 -167115
rect 149312 -167159 149368 -167115
rect 149412 -167159 149468 -167115
rect 149512 -167159 149568 -167115
rect 149612 -167159 149668 -167115
rect 149712 -167159 149768 -167115
rect 149812 -167159 149868 -167115
rect 149912 -167159 149968 -167115
rect 150012 -167159 150068 -167115
rect 150112 -167159 150168 -167115
rect 150212 -167159 150268 -167115
rect 150312 -167159 150368 -167115
rect 150412 -167159 150468 -167115
rect 150512 -167159 150568 -167115
rect 150612 -167159 150668 -167115
rect 150712 -167159 150768 -167115
rect 150812 -167159 151268 -167115
rect 151312 -167159 151368 -167115
rect 151412 -167159 151468 -167115
rect 151512 -167159 151568 -167115
rect 151612 -167159 151668 -167115
rect 151712 -167159 151768 -167115
rect 151812 -167159 151868 -167115
rect 151912 -167159 151968 -167115
rect 152012 -167159 152068 -167115
rect 152112 -167159 152168 -167115
rect 152212 -167159 152268 -167115
rect 152312 -167159 152368 -167115
rect 152412 -167159 152468 -167115
rect 152512 -167159 152568 -167115
rect 152612 -167159 152668 -167115
rect 152712 -167159 152768 -167115
rect 152812 -167159 154949 -167115
rect 142660 -168667 154949 -167159
rect 188605 -172064 192404 6200
rect 81061 -173093 81627 -173049
rect 81671 -173093 81727 -173049
rect 81771 -173093 81827 -173049
rect 81871 -173093 81927 -173049
rect 81971 -173093 82027 -173049
rect 82071 -173093 82127 -173049
rect 82171 -173093 82227 -173049
rect 82271 -173093 82327 -173049
rect 82371 -173093 82427 -173049
rect 82471 -173093 82527 -173049
rect 82571 -173093 82627 -173049
rect 82671 -173093 82727 -173049
rect 82771 -173093 82827 -173049
rect 82871 -173093 82927 -173049
rect 82971 -173093 83027 -173049
rect 83071 -173093 83127 -173049
rect 83171 -173093 83627 -173049
rect 83671 -173093 83727 -173049
rect 83771 -173093 83827 -173049
rect 83871 -173093 83927 -173049
rect 83971 -173093 84027 -173049
rect 84071 -173093 84127 -173049
rect 84171 -173093 84227 -173049
rect 84271 -173093 84327 -173049
rect 84371 -173093 84427 -173049
rect 84471 -173093 84527 -173049
rect 84571 -173093 84627 -173049
rect 84671 -173093 84727 -173049
rect 84771 -173093 84827 -173049
rect 84871 -173093 84927 -173049
rect 84971 -173093 85027 -173049
rect 85071 -173093 85127 -173049
rect 85171 -173093 85627 -173049
rect 85671 -173093 85727 -173049
rect 85771 -173093 85827 -173049
rect 85871 -173093 85927 -173049
rect 85971 -173093 86027 -173049
rect 86071 -173093 86127 -173049
rect 86171 -173093 86227 -173049
rect 86271 -173093 86327 -173049
rect 86371 -173093 86427 -173049
rect 86471 -173093 86527 -173049
rect 86571 -173093 86627 -173049
rect 86671 -173093 86727 -173049
rect 86771 -173093 86827 -173049
rect 86871 -173093 86927 -173049
rect 86971 -173093 87027 -173049
rect 87071 -173093 87127 -173049
rect 87171 -173093 87627 -173049
rect 87671 -173093 87727 -173049
rect 87771 -173093 87827 -173049
rect 87871 -173093 87927 -173049
rect 87971 -173093 88027 -173049
rect 88071 -173093 88127 -173049
rect 88171 -173093 88227 -173049
rect 88271 -173093 88327 -173049
rect 88371 -173093 88427 -173049
rect 88471 -173093 88527 -173049
rect 88571 -173093 88627 -173049
rect 88671 -173093 88727 -173049
rect 88771 -173093 88827 -173049
rect 88871 -173093 88927 -173049
rect 88971 -173093 89027 -173049
rect 89071 -173093 89127 -173049
rect 89171 -173093 89740 -173049
rect 81061 -173149 89740 -173093
rect 81061 -173193 81627 -173149
rect 81671 -173193 81727 -173149
rect 81771 -173193 81827 -173149
rect 81871 -173193 81927 -173149
rect 81971 -173193 82027 -173149
rect 82071 -173193 82127 -173149
rect 82171 -173193 82227 -173149
rect 82271 -173193 82327 -173149
rect 82371 -173193 82427 -173149
rect 82471 -173193 82527 -173149
rect 82571 -173193 82627 -173149
rect 82671 -173193 82727 -173149
rect 82771 -173193 82827 -173149
rect 82871 -173193 82927 -173149
rect 82971 -173193 83027 -173149
rect 83071 -173193 83127 -173149
rect 83171 -173193 83627 -173149
rect 83671 -173193 83727 -173149
rect 83771 -173193 83827 -173149
rect 83871 -173193 83927 -173149
rect 83971 -173193 84027 -173149
rect 84071 -173193 84127 -173149
rect 84171 -173193 84227 -173149
rect 84271 -173193 84327 -173149
rect 84371 -173193 84427 -173149
rect 84471 -173193 84527 -173149
rect 84571 -173193 84627 -173149
rect 84671 -173193 84727 -173149
rect 84771 -173193 84827 -173149
rect 84871 -173193 84927 -173149
rect 84971 -173193 85027 -173149
rect 85071 -173193 85127 -173149
rect 85171 -173193 85627 -173149
rect 85671 -173193 85727 -173149
rect 85771 -173193 85827 -173149
rect 85871 -173193 85927 -173149
rect 85971 -173193 86027 -173149
rect 86071 -173193 86127 -173149
rect 86171 -173193 86227 -173149
rect 86271 -173193 86327 -173149
rect 86371 -173193 86427 -173149
rect 86471 -173193 86527 -173149
rect 86571 -173193 86627 -173149
rect 86671 -173193 86727 -173149
rect 86771 -173193 86827 -173149
rect 86871 -173193 86927 -173149
rect 86971 -173193 87027 -173149
rect 87071 -173193 87127 -173149
rect 87171 -173193 87627 -173149
rect 87671 -173193 87727 -173149
rect 87771 -173193 87827 -173149
rect 87871 -173193 87927 -173149
rect 87971 -173193 88027 -173149
rect 88071 -173193 88127 -173149
rect 88171 -173193 88227 -173149
rect 88271 -173193 88327 -173149
rect 88371 -173193 88427 -173149
rect 88471 -173193 88527 -173149
rect 88571 -173193 88627 -173149
rect 88671 -173193 88727 -173149
rect 88771 -173193 88827 -173149
rect 88871 -173193 88927 -173149
rect 88971 -173193 89027 -173149
rect 89071 -173193 89127 -173149
rect 89171 -173193 89740 -173149
rect 81061 -173249 89740 -173193
rect 81061 -173293 81627 -173249
rect 81671 -173293 81727 -173249
rect 81771 -173293 81827 -173249
rect 81871 -173293 81927 -173249
rect 81971 -173293 82027 -173249
rect 82071 -173293 82127 -173249
rect 82171 -173293 82227 -173249
rect 82271 -173293 82327 -173249
rect 82371 -173293 82427 -173249
rect 82471 -173293 82527 -173249
rect 82571 -173293 82627 -173249
rect 82671 -173293 82727 -173249
rect 82771 -173293 82827 -173249
rect 82871 -173293 82927 -173249
rect 82971 -173293 83027 -173249
rect 83071 -173293 83127 -173249
rect 83171 -173293 83627 -173249
rect 83671 -173293 83727 -173249
rect 83771 -173293 83827 -173249
rect 83871 -173293 83927 -173249
rect 83971 -173293 84027 -173249
rect 84071 -173293 84127 -173249
rect 84171 -173293 84227 -173249
rect 84271 -173293 84327 -173249
rect 84371 -173293 84427 -173249
rect 84471 -173293 84527 -173249
rect 84571 -173293 84627 -173249
rect 84671 -173293 84727 -173249
rect 84771 -173293 84827 -173249
rect 84871 -173293 84927 -173249
rect 84971 -173293 85027 -173249
rect 85071 -173293 85127 -173249
rect 85171 -173293 85627 -173249
rect 85671 -173293 85727 -173249
rect 85771 -173293 85827 -173249
rect 85871 -173293 85927 -173249
rect 85971 -173293 86027 -173249
rect 86071 -173293 86127 -173249
rect 86171 -173293 86227 -173249
rect 86271 -173293 86327 -173249
rect 86371 -173293 86427 -173249
rect 86471 -173293 86527 -173249
rect 86571 -173293 86627 -173249
rect 86671 -173293 86727 -173249
rect 86771 -173293 86827 -173249
rect 86871 -173293 86927 -173249
rect 86971 -173293 87027 -173249
rect 87071 -173293 87127 -173249
rect 87171 -173293 87627 -173249
rect 87671 -173293 87727 -173249
rect 87771 -173293 87827 -173249
rect 87871 -173293 87927 -173249
rect 87971 -173293 88027 -173249
rect 88071 -173293 88127 -173249
rect 88171 -173293 88227 -173249
rect 88271 -173293 88327 -173249
rect 88371 -173293 88427 -173249
rect 88471 -173293 88527 -173249
rect 88571 -173293 88627 -173249
rect 88671 -173293 88727 -173249
rect 88771 -173293 88827 -173249
rect 88871 -173293 88927 -173249
rect 88971 -173293 89027 -173249
rect 89071 -173293 89127 -173249
rect 89171 -173293 89740 -173249
rect 81061 -173349 89740 -173293
rect 81061 -173393 81627 -173349
rect 81671 -173393 81727 -173349
rect 81771 -173393 81827 -173349
rect 81871 -173393 81927 -173349
rect 81971 -173393 82027 -173349
rect 82071 -173393 82127 -173349
rect 82171 -173393 82227 -173349
rect 82271 -173393 82327 -173349
rect 82371 -173393 82427 -173349
rect 82471 -173393 82527 -173349
rect 82571 -173393 82627 -173349
rect 82671 -173393 82727 -173349
rect 82771 -173393 82827 -173349
rect 82871 -173393 82927 -173349
rect 82971 -173393 83027 -173349
rect 83071 -173393 83127 -173349
rect 83171 -173393 83627 -173349
rect 83671 -173393 83727 -173349
rect 83771 -173393 83827 -173349
rect 83871 -173393 83927 -173349
rect 83971 -173393 84027 -173349
rect 84071 -173393 84127 -173349
rect 84171 -173393 84227 -173349
rect 84271 -173393 84327 -173349
rect 84371 -173393 84427 -173349
rect 84471 -173393 84527 -173349
rect 84571 -173393 84627 -173349
rect 84671 -173393 84727 -173349
rect 84771 -173393 84827 -173349
rect 84871 -173393 84927 -173349
rect 84971 -173393 85027 -173349
rect 85071 -173393 85127 -173349
rect 85171 -173393 85627 -173349
rect 85671 -173393 85727 -173349
rect 85771 -173393 85827 -173349
rect 85871 -173393 85927 -173349
rect 85971 -173393 86027 -173349
rect 86071 -173393 86127 -173349
rect 86171 -173393 86227 -173349
rect 86271 -173393 86327 -173349
rect 86371 -173393 86427 -173349
rect 86471 -173393 86527 -173349
rect 86571 -173393 86627 -173349
rect 86671 -173393 86727 -173349
rect 86771 -173393 86827 -173349
rect 86871 -173393 86927 -173349
rect 86971 -173393 87027 -173349
rect 87071 -173393 87127 -173349
rect 87171 -173393 87627 -173349
rect 87671 -173393 87727 -173349
rect 87771 -173393 87827 -173349
rect 87871 -173393 87927 -173349
rect 87971 -173393 88027 -173349
rect 88071 -173393 88127 -173349
rect 88171 -173393 88227 -173349
rect 88271 -173393 88327 -173349
rect 88371 -173393 88427 -173349
rect 88471 -173393 88527 -173349
rect 88571 -173393 88627 -173349
rect 88671 -173393 88727 -173349
rect 88771 -173393 88827 -173349
rect 88871 -173393 88927 -173349
rect 88971 -173393 89027 -173349
rect 89071 -173393 89127 -173349
rect 89171 -173393 89740 -173349
rect 81061 -173449 89740 -173393
rect 81061 -173493 81627 -173449
rect 81671 -173493 81727 -173449
rect 81771 -173493 81827 -173449
rect 81871 -173493 81927 -173449
rect 81971 -173493 82027 -173449
rect 82071 -173493 82127 -173449
rect 82171 -173493 82227 -173449
rect 82271 -173493 82327 -173449
rect 82371 -173493 82427 -173449
rect 82471 -173493 82527 -173449
rect 82571 -173493 82627 -173449
rect 82671 -173493 82727 -173449
rect 82771 -173493 82827 -173449
rect 82871 -173493 82927 -173449
rect 82971 -173493 83027 -173449
rect 83071 -173493 83127 -173449
rect 83171 -173493 83627 -173449
rect 83671 -173493 83727 -173449
rect 83771 -173493 83827 -173449
rect 83871 -173493 83927 -173449
rect 83971 -173493 84027 -173449
rect 84071 -173493 84127 -173449
rect 84171 -173493 84227 -173449
rect 84271 -173493 84327 -173449
rect 84371 -173493 84427 -173449
rect 84471 -173493 84527 -173449
rect 84571 -173493 84627 -173449
rect 84671 -173493 84727 -173449
rect 84771 -173493 84827 -173449
rect 84871 -173493 84927 -173449
rect 84971 -173493 85027 -173449
rect 85071 -173493 85127 -173449
rect 85171 -173493 85627 -173449
rect 85671 -173493 85727 -173449
rect 85771 -173493 85827 -173449
rect 85871 -173493 85927 -173449
rect 85971 -173493 86027 -173449
rect 86071 -173493 86127 -173449
rect 86171 -173493 86227 -173449
rect 86271 -173493 86327 -173449
rect 86371 -173493 86427 -173449
rect 86471 -173493 86527 -173449
rect 86571 -173493 86627 -173449
rect 86671 -173493 86727 -173449
rect 86771 -173493 86827 -173449
rect 86871 -173493 86927 -173449
rect 86971 -173493 87027 -173449
rect 87071 -173493 87127 -173449
rect 87171 -173493 87627 -173449
rect 87671 -173493 87727 -173449
rect 87771 -173493 87827 -173449
rect 87871 -173493 87927 -173449
rect 87971 -173493 88027 -173449
rect 88071 -173493 88127 -173449
rect 88171 -173493 88227 -173449
rect 88271 -173493 88327 -173449
rect 88371 -173493 88427 -173449
rect 88471 -173493 88527 -173449
rect 88571 -173493 88627 -173449
rect 88671 -173493 88727 -173449
rect 88771 -173493 88827 -173449
rect 88871 -173493 88927 -173449
rect 88971 -173493 89027 -173449
rect 89071 -173493 89127 -173449
rect 89171 -173493 89740 -173449
rect 81061 -173549 89740 -173493
rect 81061 -173593 81627 -173549
rect 81671 -173593 81727 -173549
rect 81771 -173593 81827 -173549
rect 81871 -173593 81927 -173549
rect 81971 -173593 82027 -173549
rect 82071 -173593 82127 -173549
rect 82171 -173593 82227 -173549
rect 82271 -173593 82327 -173549
rect 82371 -173593 82427 -173549
rect 82471 -173593 82527 -173549
rect 82571 -173593 82627 -173549
rect 82671 -173593 82727 -173549
rect 82771 -173593 82827 -173549
rect 82871 -173593 82927 -173549
rect 82971 -173593 83027 -173549
rect 83071 -173593 83127 -173549
rect 83171 -173593 83627 -173549
rect 83671 -173593 83727 -173549
rect 83771 -173593 83827 -173549
rect 83871 -173593 83927 -173549
rect 83971 -173593 84027 -173549
rect 84071 -173593 84127 -173549
rect 84171 -173593 84227 -173549
rect 84271 -173593 84327 -173549
rect 84371 -173593 84427 -173549
rect 84471 -173593 84527 -173549
rect 84571 -173593 84627 -173549
rect 84671 -173593 84727 -173549
rect 84771 -173593 84827 -173549
rect 84871 -173593 84927 -173549
rect 84971 -173593 85027 -173549
rect 85071 -173593 85127 -173549
rect 85171 -173593 85627 -173549
rect 85671 -173593 85727 -173549
rect 85771 -173593 85827 -173549
rect 85871 -173593 85927 -173549
rect 85971 -173593 86027 -173549
rect 86071 -173593 86127 -173549
rect 86171 -173593 86227 -173549
rect 86271 -173593 86327 -173549
rect 86371 -173593 86427 -173549
rect 86471 -173593 86527 -173549
rect 86571 -173593 86627 -173549
rect 86671 -173593 86727 -173549
rect 86771 -173593 86827 -173549
rect 86871 -173593 86927 -173549
rect 86971 -173593 87027 -173549
rect 87071 -173593 87127 -173549
rect 87171 -173593 87627 -173549
rect 87671 -173593 87727 -173549
rect 87771 -173593 87827 -173549
rect 87871 -173593 87927 -173549
rect 87971 -173593 88027 -173549
rect 88071 -173593 88127 -173549
rect 88171 -173593 88227 -173549
rect 88271 -173593 88327 -173549
rect 88371 -173593 88427 -173549
rect 88471 -173593 88527 -173549
rect 88571 -173593 88627 -173549
rect 88671 -173593 88727 -173549
rect 88771 -173593 88827 -173549
rect 88871 -173593 88927 -173549
rect 88971 -173593 89027 -173549
rect 89071 -173593 89127 -173549
rect 89171 -173593 89740 -173549
rect 81061 -173649 89740 -173593
rect 81061 -173693 81627 -173649
rect 81671 -173693 81727 -173649
rect 81771 -173693 81827 -173649
rect 81871 -173693 81927 -173649
rect 81971 -173693 82027 -173649
rect 82071 -173693 82127 -173649
rect 82171 -173693 82227 -173649
rect 82271 -173693 82327 -173649
rect 82371 -173693 82427 -173649
rect 82471 -173693 82527 -173649
rect 82571 -173693 82627 -173649
rect 82671 -173693 82727 -173649
rect 82771 -173693 82827 -173649
rect 82871 -173693 82927 -173649
rect 82971 -173693 83027 -173649
rect 83071 -173693 83127 -173649
rect 83171 -173693 83627 -173649
rect 83671 -173693 83727 -173649
rect 83771 -173693 83827 -173649
rect 83871 -173693 83927 -173649
rect 83971 -173693 84027 -173649
rect 84071 -173693 84127 -173649
rect 84171 -173693 84227 -173649
rect 84271 -173693 84327 -173649
rect 84371 -173693 84427 -173649
rect 84471 -173693 84527 -173649
rect 84571 -173693 84627 -173649
rect 84671 -173693 84727 -173649
rect 84771 -173693 84827 -173649
rect 84871 -173693 84927 -173649
rect 84971 -173693 85027 -173649
rect 85071 -173693 85127 -173649
rect 85171 -173693 85627 -173649
rect 85671 -173693 85727 -173649
rect 85771 -173693 85827 -173649
rect 85871 -173693 85927 -173649
rect 85971 -173693 86027 -173649
rect 86071 -173693 86127 -173649
rect 86171 -173693 86227 -173649
rect 86271 -173693 86327 -173649
rect 86371 -173693 86427 -173649
rect 86471 -173693 86527 -173649
rect 86571 -173693 86627 -173649
rect 86671 -173693 86727 -173649
rect 86771 -173693 86827 -173649
rect 86871 -173693 86927 -173649
rect 86971 -173693 87027 -173649
rect 87071 -173693 87127 -173649
rect 87171 -173693 87627 -173649
rect 87671 -173693 87727 -173649
rect 87771 -173693 87827 -173649
rect 87871 -173693 87927 -173649
rect 87971 -173693 88027 -173649
rect 88071 -173693 88127 -173649
rect 88171 -173693 88227 -173649
rect 88271 -173693 88327 -173649
rect 88371 -173693 88427 -173649
rect 88471 -173693 88527 -173649
rect 88571 -173693 88627 -173649
rect 88671 -173693 88727 -173649
rect 88771 -173693 88827 -173649
rect 88871 -173693 88927 -173649
rect 88971 -173693 89027 -173649
rect 89071 -173693 89127 -173649
rect 89171 -173693 89740 -173649
rect 81061 -173749 89740 -173693
rect 81061 -173793 81627 -173749
rect 81671 -173793 81727 -173749
rect 81771 -173793 81827 -173749
rect 81871 -173793 81927 -173749
rect 81971 -173793 82027 -173749
rect 82071 -173793 82127 -173749
rect 82171 -173793 82227 -173749
rect 82271 -173793 82327 -173749
rect 82371 -173793 82427 -173749
rect 82471 -173793 82527 -173749
rect 82571 -173793 82627 -173749
rect 82671 -173793 82727 -173749
rect 82771 -173793 82827 -173749
rect 82871 -173793 82927 -173749
rect 82971 -173793 83027 -173749
rect 83071 -173793 83127 -173749
rect 83171 -173793 83627 -173749
rect 83671 -173793 83727 -173749
rect 83771 -173793 83827 -173749
rect 83871 -173793 83927 -173749
rect 83971 -173793 84027 -173749
rect 84071 -173793 84127 -173749
rect 84171 -173793 84227 -173749
rect 84271 -173793 84327 -173749
rect 84371 -173793 84427 -173749
rect 84471 -173793 84527 -173749
rect 84571 -173793 84627 -173749
rect 84671 -173793 84727 -173749
rect 84771 -173793 84827 -173749
rect 84871 -173793 84927 -173749
rect 84971 -173793 85027 -173749
rect 85071 -173793 85127 -173749
rect 85171 -173793 85627 -173749
rect 85671 -173793 85727 -173749
rect 85771 -173793 85827 -173749
rect 85871 -173793 85927 -173749
rect 85971 -173793 86027 -173749
rect 86071 -173793 86127 -173749
rect 86171 -173793 86227 -173749
rect 86271 -173793 86327 -173749
rect 86371 -173793 86427 -173749
rect 86471 -173793 86527 -173749
rect 86571 -173793 86627 -173749
rect 86671 -173793 86727 -173749
rect 86771 -173793 86827 -173749
rect 86871 -173793 86927 -173749
rect 86971 -173793 87027 -173749
rect 87071 -173793 87127 -173749
rect 87171 -173793 87627 -173749
rect 87671 -173793 87727 -173749
rect 87771 -173793 87827 -173749
rect 87871 -173793 87927 -173749
rect 87971 -173793 88027 -173749
rect 88071 -173793 88127 -173749
rect 88171 -173793 88227 -173749
rect 88271 -173793 88327 -173749
rect 88371 -173793 88427 -173749
rect 88471 -173793 88527 -173749
rect 88571 -173793 88627 -173749
rect 88671 -173793 88727 -173749
rect 88771 -173793 88827 -173749
rect 88871 -173793 88927 -173749
rect 88971 -173793 89027 -173749
rect 89071 -173793 89127 -173749
rect 89171 -173793 89740 -173749
rect 81061 -173849 89740 -173793
rect 81061 -173893 81627 -173849
rect 81671 -173893 81727 -173849
rect 81771 -173893 81827 -173849
rect 81871 -173893 81927 -173849
rect 81971 -173893 82027 -173849
rect 82071 -173893 82127 -173849
rect 82171 -173893 82227 -173849
rect 82271 -173893 82327 -173849
rect 82371 -173893 82427 -173849
rect 82471 -173893 82527 -173849
rect 82571 -173893 82627 -173849
rect 82671 -173893 82727 -173849
rect 82771 -173893 82827 -173849
rect 82871 -173893 82927 -173849
rect 82971 -173893 83027 -173849
rect 83071 -173893 83127 -173849
rect 83171 -173893 83627 -173849
rect 83671 -173893 83727 -173849
rect 83771 -173893 83827 -173849
rect 83871 -173893 83927 -173849
rect 83971 -173893 84027 -173849
rect 84071 -173893 84127 -173849
rect 84171 -173893 84227 -173849
rect 84271 -173893 84327 -173849
rect 84371 -173893 84427 -173849
rect 84471 -173893 84527 -173849
rect 84571 -173893 84627 -173849
rect 84671 -173893 84727 -173849
rect 84771 -173893 84827 -173849
rect 84871 -173893 84927 -173849
rect 84971 -173893 85027 -173849
rect 85071 -173893 85127 -173849
rect 85171 -173893 85627 -173849
rect 85671 -173893 85727 -173849
rect 85771 -173893 85827 -173849
rect 85871 -173893 85927 -173849
rect 85971 -173893 86027 -173849
rect 86071 -173893 86127 -173849
rect 86171 -173893 86227 -173849
rect 86271 -173893 86327 -173849
rect 86371 -173893 86427 -173849
rect 86471 -173893 86527 -173849
rect 86571 -173893 86627 -173849
rect 86671 -173893 86727 -173849
rect 86771 -173893 86827 -173849
rect 86871 -173893 86927 -173849
rect 86971 -173893 87027 -173849
rect 87071 -173893 87127 -173849
rect 87171 -173893 87627 -173849
rect 87671 -173893 87727 -173849
rect 87771 -173893 87827 -173849
rect 87871 -173893 87927 -173849
rect 87971 -173893 88027 -173849
rect 88071 -173893 88127 -173849
rect 88171 -173893 88227 -173849
rect 88271 -173893 88327 -173849
rect 88371 -173893 88427 -173849
rect 88471 -173893 88527 -173849
rect 88571 -173893 88627 -173849
rect 88671 -173893 88727 -173849
rect 88771 -173893 88827 -173849
rect 88871 -173893 88927 -173849
rect 88971 -173893 89027 -173849
rect 89071 -173893 89127 -173849
rect 89171 -173893 89740 -173849
rect 81061 -173949 89740 -173893
rect 81061 -173993 81627 -173949
rect 81671 -173993 81727 -173949
rect 81771 -173993 81827 -173949
rect 81871 -173993 81927 -173949
rect 81971 -173993 82027 -173949
rect 82071 -173993 82127 -173949
rect 82171 -173993 82227 -173949
rect 82271 -173993 82327 -173949
rect 82371 -173993 82427 -173949
rect 82471 -173993 82527 -173949
rect 82571 -173993 82627 -173949
rect 82671 -173993 82727 -173949
rect 82771 -173993 82827 -173949
rect 82871 -173993 82927 -173949
rect 82971 -173993 83027 -173949
rect 83071 -173993 83127 -173949
rect 83171 -173993 83627 -173949
rect 83671 -173993 83727 -173949
rect 83771 -173993 83827 -173949
rect 83871 -173993 83927 -173949
rect 83971 -173993 84027 -173949
rect 84071 -173993 84127 -173949
rect 84171 -173993 84227 -173949
rect 84271 -173993 84327 -173949
rect 84371 -173993 84427 -173949
rect 84471 -173993 84527 -173949
rect 84571 -173993 84627 -173949
rect 84671 -173993 84727 -173949
rect 84771 -173993 84827 -173949
rect 84871 -173993 84927 -173949
rect 84971 -173993 85027 -173949
rect 85071 -173993 85127 -173949
rect 85171 -173993 85627 -173949
rect 85671 -173993 85727 -173949
rect 85771 -173993 85827 -173949
rect 85871 -173993 85927 -173949
rect 85971 -173993 86027 -173949
rect 86071 -173993 86127 -173949
rect 86171 -173993 86227 -173949
rect 86271 -173993 86327 -173949
rect 86371 -173993 86427 -173949
rect 86471 -173993 86527 -173949
rect 86571 -173993 86627 -173949
rect 86671 -173993 86727 -173949
rect 86771 -173993 86827 -173949
rect 86871 -173993 86927 -173949
rect 86971 -173993 87027 -173949
rect 87071 -173993 87127 -173949
rect 87171 -173993 87627 -173949
rect 87671 -173993 87727 -173949
rect 87771 -173993 87827 -173949
rect 87871 -173993 87927 -173949
rect 87971 -173993 88027 -173949
rect 88071 -173993 88127 -173949
rect 88171 -173993 88227 -173949
rect 88271 -173993 88327 -173949
rect 88371 -173993 88427 -173949
rect 88471 -173993 88527 -173949
rect 88571 -173993 88627 -173949
rect 88671 -173993 88727 -173949
rect 88771 -173993 88827 -173949
rect 88871 -173993 88927 -173949
rect 88971 -173993 89027 -173949
rect 89071 -173993 89127 -173949
rect 89171 -173993 89740 -173949
rect 81061 -174049 89740 -173993
rect 81061 -174093 81627 -174049
rect 81671 -174093 81727 -174049
rect 81771 -174093 81827 -174049
rect 81871 -174093 81927 -174049
rect 81971 -174093 82027 -174049
rect 82071 -174093 82127 -174049
rect 82171 -174093 82227 -174049
rect 82271 -174093 82327 -174049
rect 82371 -174093 82427 -174049
rect 82471 -174093 82527 -174049
rect 82571 -174093 82627 -174049
rect 82671 -174093 82727 -174049
rect 82771 -174093 82827 -174049
rect 82871 -174093 82927 -174049
rect 82971 -174093 83027 -174049
rect 83071 -174093 83127 -174049
rect 83171 -174093 83627 -174049
rect 83671 -174093 83727 -174049
rect 83771 -174093 83827 -174049
rect 83871 -174093 83927 -174049
rect 83971 -174093 84027 -174049
rect 84071 -174093 84127 -174049
rect 84171 -174093 84227 -174049
rect 84271 -174093 84327 -174049
rect 84371 -174093 84427 -174049
rect 84471 -174093 84527 -174049
rect 84571 -174093 84627 -174049
rect 84671 -174093 84727 -174049
rect 84771 -174093 84827 -174049
rect 84871 -174093 84927 -174049
rect 84971 -174093 85027 -174049
rect 85071 -174093 85127 -174049
rect 85171 -174093 85627 -174049
rect 85671 -174093 85727 -174049
rect 85771 -174093 85827 -174049
rect 85871 -174093 85927 -174049
rect 85971 -174093 86027 -174049
rect 86071 -174093 86127 -174049
rect 86171 -174093 86227 -174049
rect 86271 -174093 86327 -174049
rect 86371 -174093 86427 -174049
rect 86471 -174093 86527 -174049
rect 86571 -174093 86627 -174049
rect 86671 -174093 86727 -174049
rect 86771 -174093 86827 -174049
rect 86871 -174093 86927 -174049
rect 86971 -174093 87027 -174049
rect 87071 -174093 87127 -174049
rect 87171 -174093 87627 -174049
rect 87671 -174093 87727 -174049
rect 87771 -174093 87827 -174049
rect 87871 -174093 87927 -174049
rect 87971 -174093 88027 -174049
rect 88071 -174093 88127 -174049
rect 88171 -174093 88227 -174049
rect 88271 -174093 88327 -174049
rect 88371 -174093 88427 -174049
rect 88471 -174093 88527 -174049
rect 88571 -174093 88627 -174049
rect 88671 -174093 88727 -174049
rect 88771 -174093 88827 -174049
rect 88871 -174093 88927 -174049
rect 88971 -174093 89027 -174049
rect 89071 -174093 89127 -174049
rect 89171 -174093 89740 -174049
rect 81061 -174149 89740 -174093
rect 81061 -174193 81627 -174149
rect 81671 -174193 81727 -174149
rect 81771 -174193 81827 -174149
rect 81871 -174193 81927 -174149
rect 81971 -174193 82027 -174149
rect 82071 -174193 82127 -174149
rect 82171 -174193 82227 -174149
rect 82271 -174193 82327 -174149
rect 82371 -174193 82427 -174149
rect 82471 -174193 82527 -174149
rect 82571 -174193 82627 -174149
rect 82671 -174193 82727 -174149
rect 82771 -174193 82827 -174149
rect 82871 -174193 82927 -174149
rect 82971 -174193 83027 -174149
rect 83071 -174193 83127 -174149
rect 83171 -174193 83627 -174149
rect 83671 -174193 83727 -174149
rect 83771 -174193 83827 -174149
rect 83871 -174193 83927 -174149
rect 83971 -174193 84027 -174149
rect 84071 -174193 84127 -174149
rect 84171 -174193 84227 -174149
rect 84271 -174193 84327 -174149
rect 84371 -174193 84427 -174149
rect 84471 -174193 84527 -174149
rect 84571 -174193 84627 -174149
rect 84671 -174193 84727 -174149
rect 84771 -174193 84827 -174149
rect 84871 -174193 84927 -174149
rect 84971 -174193 85027 -174149
rect 85071 -174193 85127 -174149
rect 85171 -174193 85627 -174149
rect 85671 -174193 85727 -174149
rect 85771 -174193 85827 -174149
rect 85871 -174193 85927 -174149
rect 85971 -174193 86027 -174149
rect 86071 -174193 86127 -174149
rect 86171 -174193 86227 -174149
rect 86271 -174193 86327 -174149
rect 86371 -174193 86427 -174149
rect 86471 -174193 86527 -174149
rect 86571 -174193 86627 -174149
rect 86671 -174193 86727 -174149
rect 86771 -174193 86827 -174149
rect 86871 -174193 86927 -174149
rect 86971 -174193 87027 -174149
rect 87071 -174193 87127 -174149
rect 87171 -174193 87627 -174149
rect 87671 -174193 87727 -174149
rect 87771 -174193 87827 -174149
rect 87871 -174193 87927 -174149
rect 87971 -174193 88027 -174149
rect 88071 -174193 88127 -174149
rect 88171 -174193 88227 -174149
rect 88271 -174193 88327 -174149
rect 88371 -174193 88427 -174149
rect 88471 -174193 88527 -174149
rect 88571 -174193 88627 -174149
rect 88671 -174193 88727 -174149
rect 88771 -174193 88827 -174149
rect 88871 -174193 88927 -174149
rect 88971 -174193 89027 -174149
rect 89071 -174193 89127 -174149
rect 89171 -174193 89740 -174149
rect 81061 -174249 89740 -174193
rect 81061 -174293 81627 -174249
rect 81671 -174293 81727 -174249
rect 81771 -174293 81827 -174249
rect 81871 -174293 81927 -174249
rect 81971 -174293 82027 -174249
rect 82071 -174293 82127 -174249
rect 82171 -174293 82227 -174249
rect 82271 -174293 82327 -174249
rect 82371 -174293 82427 -174249
rect 82471 -174293 82527 -174249
rect 82571 -174293 82627 -174249
rect 82671 -174293 82727 -174249
rect 82771 -174293 82827 -174249
rect 82871 -174293 82927 -174249
rect 82971 -174293 83027 -174249
rect 83071 -174293 83127 -174249
rect 83171 -174293 83627 -174249
rect 83671 -174293 83727 -174249
rect 83771 -174293 83827 -174249
rect 83871 -174293 83927 -174249
rect 83971 -174293 84027 -174249
rect 84071 -174293 84127 -174249
rect 84171 -174293 84227 -174249
rect 84271 -174293 84327 -174249
rect 84371 -174293 84427 -174249
rect 84471 -174293 84527 -174249
rect 84571 -174293 84627 -174249
rect 84671 -174293 84727 -174249
rect 84771 -174293 84827 -174249
rect 84871 -174293 84927 -174249
rect 84971 -174293 85027 -174249
rect 85071 -174293 85127 -174249
rect 85171 -174293 85627 -174249
rect 85671 -174293 85727 -174249
rect 85771 -174293 85827 -174249
rect 85871 -174293 85927 -174249
rect 85971 -174293 86027 -174249
rect 86071 -174293 86127 -174249
rect 86171 -174293 86227 -174249
rect 86271 -174293 86327 -174249
rect 86371 -174293 86427 -174249
rect 86471 -174293 86527 -174249
rect 86571 -174293 86627 -174249
rect 86671 -174293 86727 -174249
rect 86771 -174293 86827 -174249
rect 86871 -174293 86927 -174249
rect 86971 -174293 87027 -174249
rect 87071 -174293 87127 -174249
rect 87171 -174293 87627 -174249
rect 87671 -174293 87727 -174249
rect 87771 -174293 87827 -174249
rect 87871 -174293 87927 -174249
rect 87971 -174293 88027 -174249
rect 88071 -174293 88127 -174249
rect 88171 -174293 88227 -174249
rect 88271 -174293 88327 -174249
rect 88371 -174293 88427 -174249
rect 88471 -174293 88527 -174249
rect 88571 -174293 88627 -174249
rect 88671 -174293 88727 -174249
rect 88771 -174293 88827 -174249
rect 88871 -174293 88927 -174249
rect 88971 -174293 89027 -174249
rect 89071 -174293 89127 -174249
rect 89171 -174293 89740 -174249
rect 81061 -174349 89740 -174293
rect 81061 -174393 81627 -174349
rect 81671 -174393 81727 -174349
rect 81771 -174393 81827 -174349
rect 81871 -174393 81927 -174349
rect 81971 -174393 82027 -174349
rect 82071 -174393 82127 -174349
rect 82171 -174393 82227 -174349
rect 82271 -174393 82327 -174349
rect 82371 -174393 82427 -174349
rect 82471 -174393 82527 -174349
rect 82571 -174393 82627 -174349
rect 82671 -174393 82727 -174349
rect 82771 -174393 82827 -174349
rect 82871 -174393 82927 -174349
rect 82971 -174393 83027 -174349
rect 83071 -174393 83127 -174349
rect 83171 -174393 83627 -174349
rect 83671 -174393 83727 -174349
rect 83771 -174393 83827 -174349
rect 83871 -174393 83927 -174349
rect 83971 -174393 84027 -174349
rect 84071 -174393 84127 -174349
rect 84171 -174393 84227 -174349
rect 84271 -174393 84327 -174349
rect 84371 -174393 84427 -174349
rect 84471 -174393 84527 -174349
rect 84571 -174393 84627 -174349
rect 84671 -174393 84727 -174349
rect 84771 -174393 84827 -174349
rect 84871 -174393 84927 -174349
rect 84971 -174393 85027 -174349
rect 85071 -174393 85127 -174349
rect 85171 -174393 85627 -174349
rect 85671 -174393 85727 -174349
rect 85771 -174393 85827 -174349
rect 85871 -174393 85927 -174349
rect 85971 -174393 86027 -174349
rect 86071 -174393 86127 -174349
rect 86171 -174393 86227 -174349
rect 86271 -174393 86327 -174349
rect 86371 -174393 86427 -174349
rect 86471 -174393 86527 -174349
rect 86571 -174393 86627 -174349
rect 86671 -174393 86727 -174349
rect 86771 -174393 86827 -174349
rect 86871 -174393 86927 -174349
rect 86971 -174393 87027 -174349
rect 87071 -174393 87127 -174349
rect 87171 -174393 87627 -174349
rect 87671 -174393 87727 -174349
rect 87771 -174393 87827 -174349
rect 87871 -174393 87927 -174349
rect 87971 -174393 88027 -174349
rect 88071 -174393 88127 -174349
rect 88171 -174393 88227 -174349
rect 88271 -174393 88327 -174349
rect 88371 -174393 88427 -174349
rect 88471 -174393 88527 -174349
rect 88571 -174393 88627 -174349
rect 88671 -174393 88727 -174349
rect 88771 -174393 88827 -174349
rect 88871 -174393 88927 -174349
rect 88971 -174393 89027 -174349
rect 89071 -174393 89127 -174349
rect 89171 -174393 89740 -174349
rect 81061 -174449 89740 -174393
rect 81061 -174493 81627 -174449
rect 81671 -174493 81727 -174449
rect 81771 -174493 81827 -174449
rect 81871 -174493 81927 -174449
rect 81971 -174493 82027 -174449
rect 82071 -174493 82127 -174449
rect 82171 -174493 82227 -174449
rect 82271 -174493 82327 -174449
rect 82371 -174493 82427 -174449
rect 82471 -174493 82527 -174449
rect 82571 -174493 82627 -174449
rect 82671 -174493 82727 -174449
rect 82771 -174493 82827 -174449
rect 82871 -174493 82927 -174449
rect 82971 -174493 83027 -174449
rect 83071 -174493 83127 -174449
rect 83171 -174493 83627 -174449
rect 83671 -174493 83727 -174449
rect 83771 -174493 83827 -174449
rect 83871 -174493 83927 -174449
rect 83971 -174493 84027 -174449
rect 84071 -174493 84127 -174449
rect 84171 -174493 84227 -174449
rect 84271 -174493 84327 -174449
rect 84371 -174493 84427 -174449
rect 84471 -174493 84527 -174449
rect 84571 -174493 84627 -174449
rect 84671 -174493 84727 -174449
rect 84771 -174493 84827 -174449
rect 84871 -174493 84927 -174449
rect 84971 -174493 85027 -174449
rect 85071 -174493 85127 -174449
rect 85171 -174493 85627 -174449
rect 85671 -174493 85727 -174449
rect 85771 -174493 85827 -174449
rect 85871 -174493 85927 -174449
rect 85971 -174493 86027 -174449
rect 86071 -174493 86127 -174449
rect 86171 -174493 86227 -174449
rect 86271 -174493 86327 -174449
rect 86371 -174493 86427 -174449
rect 86471 -174493 86527 -174449
rect 86571 -174493 86627 -174449
rect 86671 -174493 86727 -174449
rect 86771 -174493 86827 -174449
rect 86871 -174493 86927 -174449
rect 86971 -174493 87027 -174449
rect 87071 -174493 87127 -174449
rect 87171 -174493 87627 -174449
rect 87671 -174493 87727 -174449
rect 87771 -174493 87827 -174449
rect 87871 -174493 87927 -174449
rect 87971 -174493 88027 -174449
rect 88071 -174493 88127 -174449
rect 88171 -174493 88227 -174449
rect 88271 -174493 88327 -174449
rect 88371 -174493 88427 -174449
rect 88471 -174493 88527 -174449
rect 88571 -174493 88627 -174449
rect 88671 -174493 88727 -174449
rect 88771 -174493 88827 -174449
rect 88871 -174493 88927 -174449
rect 88971 -174493 89027 -174449
rect 89071 -174493 89127 -174449
rect 89171 -174493 89740 -174449
rect 81061 -174549 89740 -174493
rect 81061 -174593 81627 -174549
rect 81671 -174593 81727 -174549
rect 81771 -174593 81827 -174549
rect 81871 -174593 81927 -174549
rect 81971 -174593 82027 -174549
rect 82071 -174593 82127 -174549
rect 82171 -174593 82227 -174549
rect 82271 -174593 82327 -174549
rect 82371 -174593 82427 -174549
rect 82471 -174593 82527 -174549
rect 82571 -174593 82627 -174549
rect 82671 -174593 82727 -174549
rect 82771 -174593 82827 -174549
rect 82871 -174593 82927 -174549
rect 82971 -174593 83027 -174549
rect 83071 -174593 83127 -174549
rect 83171 -174593 83627 -174549
rect 83671 -174593 83727 -174549
rect 83771 -174593 83827 -174549
rect 83871 -174593 83927 -174549
rect 83971 -174593 84027 -174549
rect 84071 -174593 84127 -174549
rect 84171 -174593 84227 -174549
rect 84271 -174593 84327 -174549
rect 84371 -174593 84427 -174549
rect 84471 -174593 84527 -174549
rect 84571 -174593 84627 -174549
rect 84671 -174593 84727 -174549
rect 84771 -174593 84827 -174549
rect 84871 -174593 84927 -174549
rect 84971 -174593 85027 -174549
rect 85071 -174593 85127 -174549
rect 85171 -174593 85627 -174549
rect 85671 -174593 85727 -174549
rect 85771 -174593 85827 -174549
rect 85871 -174593 85927 -174549
rect 85971 -174593 86027 -174549
rect 86071 -174593 86127 -174549
rect 86171 -174593 86227 -174549
rect 86271 -174593 86327 -174549
rect 86371 -174593 86427 -174549
rect 86471 -174593 86527 -174549
rect 86571 -174593 86627 -174549
rect 86671 -174593 86727 -174549
rect 86771 -174593 86827 -174549
rect 86871 -174593 86927 -174549
rect 86971 -174593 87027 -174549
rect 87071 -174593 87127 -174549
rect 87171 -174593 87627 -174549
rect 87671 -174593 87727 -174549
rect 87771 -174593 87827 -174549
rect 87871 -174593 87927 -174549
rect 87971 -174593 88027 -174549
rect 88071 -174593 88127 -174549
rect 88171 -174593 88227 -174549
rect 88271 -174593 88327 -174549
rect 88371 -174593 88427 -174549
rect 88471 -174593 88527 -174549
rect 88571 -174593 88627 -174549
rect 88671 -174593 88727 -174549
rect 88771 -174593 88827 -174549
rect 88871 -174593 88927 -174549
rect 88971 -174593 89027 -174549
rect 89071 -174593 89127 -174549
rect 89171 -174593 89740 -174549
rect 81061 -175655 89740 -174593
rect 162407 -172989 192404 -172064
rect 162407 -173033 165525 -172989
rect 165569 -173033 165625 -172989
rect 165669 -173033 165725 -172989
rect 165769 -173033 165825 -172989
rect 165869 -173033 165925 -172989
rect 165969 -173033 166025 -172989
rect 166069 -173033 166125 -172989
rect 166169 -173033 166225 -172989
rect 166269 -173033 166325 -172989
rect 166369 -173033 166425 -172989
rect 166469 -173033 166525 -172989
rect 166569 -173033 166625 -172989
rect 166669 -173033 166725 -172989
rect 166769 -173033 166825 -172989
rect 166869 -173033 166925 -172989
rect 166969 -173033 167025 -172989
rect 167069 -173033 167525 -172989
rect 167569 -173033 167625 -172989
rect 167669 -173033 167725 -172989
rect 167769 -173033 167825 -172989
rect 167869 -173033 167925 -172989
rect 167969 -173033 168025 -172989
rect 168069 -173033 168125 -172989
rect 168169 -173033 168225 -172989
rect 168269 -173033 168325 -172989
rect 168369 -173033 168425 -172989
rect 168469 -173033 168525 -172989
rect 168569 -173033 168625 -172989
rect 168669 -173033 168725 -172989
rect 168769 -173033 168825 -172989
rect 168869 -173033 168925 -172989
rect 168969 -173033 169025 -172989
rect 169069 -173033 169525 -172989
rect 169569 -173033 169625 -172989
rect 169669 -173033 169725 -172989
rect 169769 -173033 169825 -172989
rect 169869 -173033 169925 -172989
rect 169969 -173033 170025 -172989
rect 170069 -173033 170125 -172989
rect 170169 -173033 170225 -172989
rect 170269 -173033 170325 -172989
rect 170369 -173033 170425 -172989
rect 170469 -173033 170525 -172989
rect 170569 -173033 170625 -172989
rect 170669 -173033 170725 -172989
rect 170769 -173033 170825 -172989
rect 170869 -173033 170925 -172989
rect 170969 -173033 171025 -172989
rect 171069 -173033 171525 -172989
rect 171569 -173033 171625 -172989
rect 171669 -173033 171725 -172989
rect 171769 -173033 171825 -172989
rect 171869 -173033 171925 -172989
rect 171969 -173033 172025 -172989
rect 172069 -173033 172125 -172989
rect 172169 -173033 172225 -172989
rect 172269 -173033 172325 -172989
rect 172369 -173033 172425 -172989
rect 172469 -173033 172525 -172989
rect 172569 -173033 172625 -172989
rect 172669 -173033 172725 -172989
rect 172769 -173033 172825 -172989
rect 172869 -173033 172925 -172989
rect 172969 -173033 173025 -172989
rect 173069 -173033 192404 -172989
rect 162407 -173089 192404 -173033
rect 162407 -173133 165525 -173089
rect 165569 -173133 165625 -173089
rect 165669 -173133 165725 -173089
rect 165769 -173133 165825 -173089
rect 165869 -173133 165925 -173089
rect 165969 -173133 166025 -173089
rect 166069 -173133 166125 -173089
rect 166169 -173133 166225 -173089
rect 166269 -173133 166325 -173089
rect 166369 -173133 166425 -173089
rect 166469 -173133 166525 -173089
rect 166569 -173133 166625 -173089
rect 166669 -173133 166725 -173089
rect 166769 -173133 166825 -173089
rect 166869 -173133 166925 -173089
rect 166969 -173133 167025 -173089
rect 167069 -173133 167525 -173089
rect 167569 -173133 167625 -173089
rect 167669 -173133 167725 -173089
rect 167769 -173133 167825 -173089
rect 167869 -173133 167925 -173089
rect 167969 -173133 168025 -173089
rect 168069 -173133 168125 -173089
rect 168169 -173133 168225 -173089
rect 168269 -173133 168325 -173089
rect 168369 -173133 168425 -173089
rect 168469 -173133 168525 -173089
rect 168569 -173133 168625 -173089
rect 168669 -173133 168725 -173089
rect 168769 -173133 168825 -173089
rect 168869 -173133 168925 -173089
rect 168969 -173133 169025 -173089
rect 169069 -173133 169525 -173089
rect 169569 -173133 169625 -173089
rect 169669 -173133 169725 -173089
rect 169769 -173133 169825 -173089
rect 169869 -173133 169925 -173089
rect 169969 -173133 170025 -173089
rect 170069 -173133 170125 -173089
rect 170169 -173133 170225 -173089
rect 170269 -173133 170325 -173089
rect 170369 -173133 170425 -173089
rect 170469 -173133 170525 -173089
rect 170569 -173133 170625 -173089
rect 170669 -173133 170725 -173089
rect 170769 -173133 170825 -173089
rect 170869 -173133 170925 -173089
rect 170969 -173133 171025 -173089
rect 171069 -173133 171525 -173089
rect 171569 -173133 171625 -173089
rect 171669 -173133 171725 -173089
rect 171769 -173133 171825 -173089
rect 171869 -173133 171925 -173089
rect 171969 -173133 172025 -173089
rect 172069 -173133 172125 -173089
rect 172169 -173133 172225 -173089
rect 172269 -173133 172325 -173089
rect 172369 -173133 172425 -173089
rect 172469 -173133 172525 -173089
rect 172569 -173133 172625 -173089
rect 172669 -173133 172725 -173089
rect 172769 -173133 172825 -173089
rect 172869 -173133 172925 -173089
rect 172969 -173133 173025 -173089
rect 173069 -173133 192404 -173089
rect 162407 -173189 192404 -173133
rect 162407 -173233 165525 -173189
rect 165569 -173233 165625 -173189
rect 165669 -173233 165725 -173189
rect 165769 -173233 165825 -173189
rect 165869 -173233 165925 -173189
rect 165969 -173233 166025 -173189
rect 166069 -173233 166125 -173189
rect 166169 -173233 166225 -173189
rect 166269 -173233 166325 -173189
rect 166369 -173233 166425 -173189
rect 166469 -173233 166525 -173189
rect 166569 -173233 166625 -173189
rect 166669 -173233 166725 -173189
rect 166769 -173233 166825 -173189
rect 166869 -173233 166925 -173189
rect 166969 -173233 167025 -173189
rect 167069 -173233 167525 -173189
rect 167569 -173233 167625 -173189
rect 167669 -173233 167725 -173189
rect 167769 -173233 167825 -173189
rect 167869 -173233 167925 -173189
rect 167969 -173233 168025 -173189
rect 168069 -173233 168125 -173189
rect 168169 -173233 168225 -173189
rect 168269 -173233 168325 -173189
rect 168369 -173233 168425 -173189
rect 168469 -173233 168525 -173189
rect 168569 -173233 168625 -173189
rect 168669 -173233 168725 -173189
rect 168769 -173233 168825 -173189
rect 168869 -173233 168925 -173189
rect 168969 -173233 169025 -173189
rect 169069 -173233 169525 -173189
rect 169569 -173233 169625 -173189
rect 169669 -173233 169725 -173189
rect 169769 -173233 169825 -173189
rect 169869 -173233 169925 -173189
rect 169969 -173233 170025 -173189
rect 170069 -173233 170125 -173189
rect 170169 -173233 170225 -173189
rect 170269 -173233 170325 -173189
rect 170369 -173233 170425 -173189
rect 170469 -173233 170525 -173189
rect 170569 -173233 170625 -173189
rect 170669 -173233 170725 -173189
rect 170769 -173233 170825 -173189
rect 170869 -173233 170925 -173189
rect 170969 -173233 171025 -173189
rect 171069 -173233 171525 -173189
rect 171569 -173233 171625 -173189
rect 171669 -173233 171725 -173189
rect 171769 -173233 171825 -173189
rect 171869 -173233 171925 -173189
rect 171969 -173233 172025 -173189
rect 172069 -173233 172125 -173189
rect 172169 -173233 172225 -173189
rect 172269 -173233 172325 -173189
rect 172369 -173233 172425 -173189
rect 172469 -173233 172525 -173189
rect 172569 -173233 172625 -173189
rect 172669 -173233 172725 -173189
rect 172769 -173233 172825 -173189
rect 172869 -173233 172925 -173189
rect 172969 -173233 173025 -173189
rect 173069 -173233 192404 -173189
rect 162407 -173289 192404 -173233
rect 162407 -173333 165525 -173289
rect 165569 -173333 165625 -173289
rect 165669 -173333 165725 -173289
rect 165769 -173333 165825 -173289
rect 165869 -173333 165925 -173289
rect 165969 -173333 166025 -173289
rect 166069 -173333 166125 -173289
rect 166169 -173333 166225 -173289
rect 166269 -173333 166325 -173289
rect 166369 -173333 166425 -173289
rect 166469 -173333 166525 -173289
rect 166569 -173333 166625 -173289
rect 166669 -173333 166725 -173289
rect 166769 -173333 166825 -173289
rect 166869 -173333 166925 -173289
rect 166969 -173333 167025 -173289
rect 167069 -173333 167525 -173289
rect 167569 -173333 167625 -173289
rect 167669 -173333 167725 -173289
rect 167769 -173333 167825 -173289
rect 167869 -173333 167925 -173289
rect 167969 -173333 168025 -173289
rect 168069 -173333 168125 -173289
rect 168169 -173333 168225 -173289
rect 168269 -173333 168325 -173289
rect 168369 -173333 168425 -173289
rect 168469 -173333 168525 -173289
rect 168569 -173333 168625 -173289
rect 168669 -173333 168725 -173289
rect 168769 -173333 168825 -173289
rect 168869 -173333 168925 -173289
rect 168969 -173333 169025 -173289
rect 169069 -173333 169525 -173289
rect 169569 -173333 169625 -173289
rect 169669 -173333 169725 -173289
rect 169769 -173333 169825 -173289
rect 169869 -173333 169925 -173289
rect 169969 -173333 170025 -173289
rect 170069 -173333 170125 -173289
rect 170169 -173333 170225 -173289
rect 170269 -173333 170325 -173289
rect 170369 -173333 170425 -173289
rect 170469 -173333 170525 -173289
rect 170569 -173333 170625 -173289
rect 170669 -173333 170725 -173289
rect 170769 -173333 170825 -173289
rect 170869 -173333 170925 -173289
rect 170969 -173333 171025 -173289
rect 171069 -173333 171525 -173289
rect 171569 -173333 171625 -173289
rect 171669 -173333 171725 -173289
rect 171769 -173333 171825 -173289
rect 171869 -173333 171925 -173289
rect 171969 -173333 172025 -173289
rect 172069 -173333 172125 -173289
rect 172169 -173333 172225 -173289
rect 172269 -173333 172325 -173289
rect 172369 -173333 172425 -173289
rect 172469 -173333 172525 -173289
rect 172569 -173333 172625 -173289
rect 172669 -173333 172725 -173289
rect 172769 -173333 172825 -173289
rect 172869 -173333 172925 -173289
rect 172969 -173333 173025 -173289
rect 173069 -173333 192404 -173289
rect 162407 -173389 192404 -173333
rect 162407 -173433 165525 -173389
rect 165569 -173433 165625 -173389
rect 165669 -173433 165725 -173389
rect 165769 -173433 165825 -173389
rect 165869 -173433 165925 -173389
rect 165969 -173433 166025 -173389
rect 166069 -173433 166125 -173389
rect 166169 -173433 166225 -173389
rect 166269 -173433 166325 -173389
rect 166369 -173433 166425 -173389
rect 166469 -173433 166525 -173389
rect 166569 -173433 166625 -173389
rect 166669 -173433 166725 -173389
rect 166769 -173433 166825 -173389
rect 166869 -173433 166925 -173389
rect 166969 -173433 167025 -173389
rect 167069 -173433 167525 -173389
rect 167569 -173433 167625 -173389
rect 167669 -173433 167725 -173389
rect 167769 -173433 167825 -173389
rect 167869 -173433 167925 -173389
rect 167969 -173433 168025 -173389
rect 168069 -173433 168125 -173389
rect 168169 -173433 168225 -173389
rect 168269 -173433 168325 -173389
rect 168369 -173433 168425 -173389
rect 168469 -173433 168525 -173389
rect 168569 -173433 168625 -173389
rect 168669 -173433 168725 -173389
rect 168769 -173433 168825 -173389
rect 168869 -173433 168925 -173389
rect 168969 -173433 169025 -173389
rect 169069 -173433 169525 -173389
rect 169569 -173433 169625 -173389
rect 169669 -173433 169725 -173389
rect 169769 -173433 169825 -173389
rect 169869 -173433 169925 -173389
rect 169969 -173433 170025 -173389
rect 170069 -173433 170125 -173389
rect 170169 -173433 170225 -173389
rect 170269 -173433 170325 -173389
rect 170369 -173433 170425 -173389
rect 170469 -173433 170525 -173389
rect 170569 -173433 170625 -173389
rect 170669 -173433 170725 -173389
rect 170769 -173433 170825 -173389
rect 170869 -173433 170925 -173389
rect 170969 -173433 171025 -173389
rect 171069 -173433 171525 -173389
rect 171569 -173433 171625 -173389
rect 171669 -173433 171725 -173389
rect 171769 -173433 171825 -173389
rect 171869 -173433 171925 -173389
rect 171969 -173433 172025 -173389
rect 172069 -173433 172125 -173389
rect 172169 -173433 172225 -173389
rect 172269 -173433 172325 -173389
rect 172369 -173433 172425 -173389
rect 172469 -173433 172525 -173389
rect 172569 -173433 172625 -173389
rect 172669 -173433 172725 -173389
rect 172769 -173433 172825 -173389
rect 172869 -173433 172925 -173389
rect 172969 -173433 173025 -173389
rect 173069 -173433 192404 -173389
rect 162407 -173489 192404 -173433
rect 162407 -173533 165525 -173489
rect 165569 -173533 165625 -173489
rect 165669 -173533 165725 -173489
rect 165769 -173533 165825 -173489
rect 165869 -173533 165925 -173489
rect 165969 -173533 166025 -173489
rect 166069 -173533 166125 -173489
rect 166169 -173533 166225 -173489
rect 166269 -173533 166325 -173489
rect 166369 -173533 166425 -173489
rect 166469 -173533 166525 -173489
rect 166569 -173533 166625 -173489
rect 166669 -173533 166725 -173489
rect 166769 -173533 166825 -173489
rect 166869 -173533 166925 -173489
rect 166969 -173533 167025 -173489
rect 167069 -173533 167525 -173489
rect 167569 -173533 167625 -173489
rect 167669 -173533 167725 -173489
rect 167769 -173533 167825 -173489
rect 167869 -173533 167925 -173489
rect 167969 -173533 168025 -173489
rect 168069 -173533 168125 -173489
rect 168169 -173533 168225 -173489
rect 168269 -173533 168325 -173489
rect 168369 -173533 168425 -173489
rect 168469 -173533 168525 -173489
rect 168569 -173533 168625 -173489
rect 168669 -173533 168725 -173489
rect 168769 -173533 168825 -173489
rect 168869 -173533 168925 -173489
rect 168969 -173533 169025 -173489
rect 169069 -173533 169525 -173489
rect 169569 -173533 169625 -173489
rect 169669 -173533 169725 -173489
rect 169769 -173533 169825 -173489
rect 169869 -173533 169925 -173489
rect 169969 -173533 170025 -173489
rect 170069 -173533 170125 -173489
rect 170169 -173533 170225 -173489
rect 170269 -173533 170325 -173489
rect 170369 -173533 170425 -173489
rect 170469 -173533 170525 -173489
rect 170569 -173533 170625 -173489
rect 170669 -173533 170725 -173489
rect 170769 -173533 170825 -173489
rect 170869 -173533 170925 -173489
rect 170969 -173533 171025 -173489
rect 171069 -173533 171525 -173489
rect 171569 -173533 171625 -173489
rect 171669 -173533 171725 -173489
rect 171769 -173533 171825 -173489
rect 171869 -173533 171925 -173489
rect 171969 -173533 172025 -173489
rect 172069 -173533 172125 -173489
rect 172169 -173533 172225 -173489
rect 172269 -173533 172325 -173489
rect 172369 -173533 172425 -173489
rect 172469 -173533 172525 -173489
rect 172569 -173533 172625 -173489
rect 172669 -173533 172725 -173489
rect 172769 -173533 172825 -173489
rect 172869 -173533 172925 -173489
rect 172969 -173533 173025 -173489
rect 173069 -173533 192404 -173489
rect 162407 -173589 192404 -173533
rect 162407 -173633 165525 -173589
rect 165569 -173633 165625 -173589
rect 165669 -173633 165725 -173589
rect 165769 -173633 165825 -173589
rect 165869 -173633 165925 -173589
rect 165969 -173633 166025 -173589
rect 166069 -173633 166125 -173589
rect 166169 -173633 166225 -173589
rect 166269 -173633 166325 -173589
rect 166369 -173633 166425 -173589
rect 166469 -173633 166525 -173589
rect 166569 -173633 166625 -173589
rect 166669 -173633 166725 -173589
rect 166769 -173633 166825 -173589
rect 166869 -173633 166925 -173589
rect 166969 -173633 167025 -173589
rect 167069 -173633 167525 -173589
rect 167569 -173633 167625 -173589
rect 167669 -173633 167725 -173589
rect 167769 -173633 167825 -173589
rect 167869 -173633 167925 -173589
rect 167969 -173633 168025 -173589
rect 168069 -173633 168125 -173589
rect 168169 -173633 168225 -173589
rect 168269 -173633 168325 -173589
rect 168369 -173633 168425 -173589
rect 168469 -173633 168525 -173589
rect 168569 -173633 168625 -173589
rect 168669 -173633 168725 -173589
rect 168769 -173633 168825 -173589
rect 168869 -173633 168925 -173589
rect 168969 -173633 169025 -173589
rect 169069 -173633 169525 -173589
rect 169569 -173633 169625 -173589
rect 169669 -173633 169725 -173589
rect 169769 -173633 169825 -173589
rect 169869 -173633 169925 -173589
rect 169969 -173633 170025 -173589
rect 170069 -173633 170125 -173589
rect 170169 -173633 170225 -173589
rect 170269 -173633 170325 -173589
rect 170369 -173633 170425 -173589
rect 170469 -173633 170525 -173589
rect 170569 -173633 170625 -173589
rect 170669 -173633 170725 -173589
rect 170769 -173633 170825 -173589
rect 170869 -173633 170925 -173589
rect 170969 -173633 171025 -173589
rect 171069 -173633 171525 -173589
rect 171569 -173633 171625 -173589
rect 171669 -173633 171725 -173589
rect 171769 -173633 171825 -173589
rect 171869 -173633 171925 -173589
rect 171969 -173633 172025 -173589
rect 172069 -173633 172125 -173589
rect 172169 -173633 172225 -173589
rect 172269 -173633 172325 -173589
rect 172369 -173633 172425 -173589
rect 172469 -173633 172525 -173589
rect 172569 -173633 172625 -173589
rect 172669 -173633 172725 -173589
rect 172769 -173633 172825 -173589
rect 172869 -173633 172925 -173589
rect 172969 -173633 173025 -173589
rect 173069 -173633 192404 -173589
rect 162407 -173689 192404 -173633
rect 162407 -173733 165525 -173689
rect 165569 -173733 165625 -173689
rect 165669 -173733 165725 -173689
rect 165769 -173733 165825 -173689
rect 165869 -173733 165925 -173689
rect 165969 -173733 166025 -173689
rect 166069 -173733 166125 -173689
rect 166169 -173733 166225 -173689
rect 166269 -173733 166325 -173689
rect 166369 -173733 166425 -173689
rect 166469 -173733 166525 -173689
rect 166569 -173733 166625 -173689
rect 166669 -173733 166725 -173689
rect 166769 -173733 166825 -173689
rect 166869 -173733 166925 -173689
rect 166969 -173733 167025 -173689
rect 167069 -173733 167525 -173689
rect 167569 -173733 167625 -173689
rect 167669 -173733 167725 -173689
rect 167769 -173733 167825 -173689
rect 167869 -173733 167925 -173689
rect 167969 -173733 168025 -173689
rect 168069 -173733 168125 -173689
rect 168169 -173733 168225 -173689
rect 168269 -173733 168325 -173689
rect 168369 -173733 168425 -173689
rect 168469 -173733 168525 -173689
rect 168569 -173733 168625 -173689
rect 168669 -173733 168725 -173689
rect 168769 -173733 168825 -173689
rect 168869 -173733 168925 -173689
rect 168969 -173733 169025 -173689
rect 169069 -173733 169525 -173689
rect 169569 -173733 169625 -173689
rect 169669 -173733 169725 -173689
rect 169769 -173733 169825 -173689
rect 169869 -173733 169925 -173689
rect 169969 -173733 170025 -173689
rect 170069 -173733 170125 -173689
rect 170169 -173733 170225 -173689
rect 170269 -173733 170325 -173689
rect 170369 -173733 170425 -173689
rect 170469 -173733 170525 -173689
rect 170569 -173733 170625 -173689
rect 170669 -173733 170725 -173689
rect 170769 -173733 170825 -173689
rect 170869 -173733 170925 -173689
rect 170969 -173733 171025 -173689
rect 171069 -173733 171525 -173689
rect 171569 -173733 171625 -173689
rect 171669 -173733 171725 -173689
rect 171769 -173733 171825 -173689
rect 171869 -173733 171925 -173689
rect 171969 -173733 172025 -173689
rect 172069 -173733 172125 -173689
rect 172169 -173733 172225 -173689
rect 172269 -173733 172325 -173689
rect 172369 -173733 172425 -173689
rect 172469 -173733 172525 -173689
rect 172569 -173733 172625 -173689
rect 172669 -173733 172725 -173689
rect 172769 -173733 172825 -173689
rect 172869 -173733 172925 -173689
rect 172969 -173733 173025 -173689
rect 173069 -173733 192404 -173689
rect 162407 -173789 192404 -173733
rect 162407 -173833 165525 -173789
rect 165569 -173833 165625 -173789
rect 165669 -173833 165725 -173789
rect 165769 -173833 165825 -173789
rect 165869 -173833 165925 -173789
rect 165969 -173833 166025 -173789
rect 166069 -173833 166125 -173789
rect 166169 -173833 166225 -173789
rect 166269 -173833 166325 -173789
rect 166369 -173833 166425 -173789
rect 166469 -173833 166525 -173789
rect 166569 -173833 166625 -173789
rect 166669 -173833 166725 -173789
rect 166769 -173833 166825 -173789
rect 166869 -173833 166925 -173789
rect 166969 -173833 167025 -173789
rect 167069 -173833 167525 -173789
rect 167569 -173833 167625 -173789
rect 167669 -173833 167725 -173789
rect 167769 -173833 167825 -173789
rect 167869 -173833 167925 -173789
rect 167969 -173833 168025 -173789
rect 168069 -173833 168125 -173789
rect 168169 -173833 168225 -173789
rect 168269 -173833 168325 -173789
rect 168369 -173833 168425 -173789
rect 168469 -173833 168525 -173789
rect 168569 -173833 168625 -173789
rect 168669 -173833 168725 -173789
rect 168769 -173833 168825 -173789
rect 168869 -173833 168925 -173789
rect 168969 -173833 169025 -173789
rect 169069 -173833 169525 -173789
rect 169569 -173833 169625 -173789
rect 169669 -173833 169725 -173789
rect 169769 -173833 169825 -173789
rect 169869 -173833 169925 -173789
rect 169969 -173833 170025 -173789
rect 170069 -173833 170125 -173789
rect 170169 -173833 170225 -173789
rect 170269 -173833 170325 -173789
rect 170369 -173833 170425 -173789
rect 170469 -173833 170525 -173789
rect 170569 -173833 170625 -173789
rect 170669 -173833 170725 -173789
rect 170769 -173833 170825 -173789
rect 170869 -173833 170925 -173789
rect 170969 -173833 171025 -173789
rect 171069 -173833 171525 -173789
rect 171569 -173833 171625 -173789
rect 171669 -173833 171725 -173789
rect 171769 -173833 171825 -173789
rect 171869 -173833 171925 -173789
rect 171969 -173833 172025 -173789
rect 172069 -173833 172125 -173789
rect 172169 -173833 172225 -173789
rect 172269 -173833 172325 -173789
rect 172369 -173833 172425 -173789
rect 172469 -173833 172525 -173789
rect 172569 -173833 172625 -173789
rect 172669 -173833 172725 -173789
rect 172769 -173833 172825 -173789
rect 172869 -173833 172925 -173789
rect 172969 -173833 173025 -173789
rect 173069 -173833 192404 -173789
rect 162407 -173889 192404 -173833
rect 162407 -173933 165525 -173889
rect 165569 -173933 165625 -173889
rect 165669 -173933 165725 -173889
rect 165769 -173933 165825 -173889
rect 165869 -173933 165925 -173889
rect 165969 -173933 166025 -173889
rect 166069 -173933 166125 -173889
rect 166169 -173933 166225 -173889
rect 166269 -173933 166325 -173889
rect 166369 -173933 166425 -173889
rect 166469 -173933 166525 -173889
rect 166569 -173933 166625 -173889
rect 166669 -173933 166725 -173889
rect 166769 -173933 166825 -173889
rect 166869 -173933 166925 -173889
rect 166969 -173933 167025 -173889
rect 167069 -173933 167525 -173889
rect 167569 -173933 167625 -173889
rect 167669 -173933 167725 -173889
rect 167769 -173933 167825 -173889
rect 167869 -173933 167925 -173889
rect 167969 -173933 168025 -173889
rect 168069 -173933 168125 -173889
rect 168169 -173933 168225 -173889
rect 168269 -173933 168325 -173889
rect 168369 -173933 168425 -173889
rect 168469 -173933 168525 -173889
rect 168569 -173933 168625 -173889
rect 168669 -173933 168725 -173889
rect 168769 -173933 168825 -173889
rect 168869 -173933 168925 -173889
rect 168969 -173933 169025 -173889
rect 169069 -173933 169525 -173889
rect 169569 -173933 169625 -173889
rect 169669 -173933 169725 -173889
rect 169769 -173933 169825 -173889
rect 169869 -173933 169925 -173889
rect 169969 -173933 170025 -173889
rect 170069 -173933 170125 -173889
rect 170169 -173933 170225 -173889
rect 170269 -173933 170325 -173889
rect 170369 -173933 170425 -173889
rect 170469 -173933 170525 -173889
rect 170569 -173933 170625 -173889
rect 170669 -173933 170725 -173889
rect 170769 -173933 170825 -173889
rect 170869 -173933 170925 -173889
rect 170969 -173933 171025 -173889
rect 171069 -173933 171525 -173889
rect 171569 -173933 171625 -173889
rect 171669 -173933 171725 -173889
rect 171769 -173933 171825 -173889
rect 171869 -173933 171925 -173889
rect 171969 -173933 172025 -173889
rect 172069 -173933 172125 -173889
rect 172169 -173933 172225 -173889
rect 172269 -173933 172325 -173889
rect 172369 -173933 172425 -173889
rect 172469 -173933 172525 -173889
rect 172569 -173933 172625 -173889
rect 172669 -173933 172725 -173889
rect 172769 -173933 172825 -173889
rect 172869 -173933 172925 -173889
rect 172969 -173933 173025 -173889
rect 173069 -173933 192404 -173889
rect 162407 -173989 192404 -173933
rect 162407 -174033 165525 -173989
rect 165569 -174033 165625 -173989
rect 165669 -174033 165725 -173989
rect 165769 -174033 165825 -173989
rect 165869 -174033 165925 -173989
rect 165969 -174033 166025 -173989
rect 166069 -174033 166125 -173989
rect 166169 -174033 166225 -173989
rect 166269 -174033 166325 -173989
rect 166369 -174033 166425 -173989
rect 166469 -174033 166525 -173989
rect 166569 -174033 166625 -173989
rect 166669 -174033 166725 -173989
rect 166769 -174033 166825 -173989
rect 166869 -174033 166925 -173989
rect 166969 -174033 167025 -173989
rect 167069 -174033 167525 -173989
rect 167569 -174033 167625 -173989
rect 167669 -174033 167725 -173989
rect 167769 -174033 167825 -173989
rect 167869 -174033 167925 -173989
rect 167969 -174033 168025 -173989
rect 168069 -174033 168125 -173989
rect 168169 -174033 168225 -173989
rect 168269 -174033 168325 -173989
rect 168369 -174033 168425 -173989
rect 168469 -174033 168525 -173989
rect 168569 -174033 168625 -173989
rect 168669 -174033 168725 -173989
rect 168769 -174033 168825 -173989
rect 168869 -174033 168925 -173989
rect 168969 -174033 169025 -173989
rect 169069 -174033 169525 -173989
rect 169569 -174033 169625 -173989
rect 169669 -174033 169725 -173989
rect 169769 -174033 169825 -173989
rect 169869 -174033 169925 -173989
rect 169969 -174033 170025 -173989
rect 170069 -174033 170125 -173989
rect 170169 -174033 170225 -173989
rect 170269 -174033 170325 -173989
rect 170369 -174033 170425 -173989
rect 170469 -174033 170525 -173989
rect 170569 -174033 170625 -173989
rect 170669 -174033 170725 -173989
rect 170769 -174033 170825 -173989
rect 170869 -174033 170925 -173989
rect 170969 -174033 171025 -173989
rect 171069 -174033 171525 -173989
rect 171569 -174033 171625 -173989
rect 171669 -174033 171725 -173989
rect 171769 -174033 171825 -173989
rect 171869 -174033 171925 -173989
rect 171969 -174033 172025 -173989
rect 172069 -174033 172125 -173989
rect 172169 -174033 172225 -173989
rect 172269 -174033 172325 -173989
rect 172369 -174033 172425 -173989
rect 172469 -174033 172525 -173989
rect 172569 -174033 172625 -173989
rect 172669 -174033 172725 -173989
rect 172769 -174033 172825 -173989
rect 172869 -174033 172925 -173989
rect 172969 -174033 173025 -173989
rect 173069 -174033 192404 -173989
rect 162407 -174089 192404 -174033
rect 162407 -174133 165525 -174089
rect 165569 -174133 165625 -174089
rect 165669 -174133 165725 -174089
rect 165769 -174133 165825 -174089
rect 165869 -174133 165925 -174089
rect 165969 -174133 166025 -174089
rect 166069 -174133 166125 -174089
rect 166169 -174133 166225 -174089
rect 166269 -174133 166325 -174089
rect 166369 -174133 166425 -174089
rect 166469 -174133 166525 -174089
rect 166569 -174133 166625 -174089
rect 166669 -174133 166725 -174089
rect 166769 -174133 166825 -174089
rect 166869 -174133 166925 -174089
rect 166969 -174133 167025 -174089
rect 167069 -174133 167525 -174089
rect 167569 -174133 167625 -174089
rect 167669 -174133 167725 -174089
rect 167769 -174133 167825 -174089
rect 167869 -174133 167925 -174089
rect 167969 -174133 168025 -174089
rect 168069 -174133 168125 -174089
rect 168169 -174133 168225 -174089
rect 168269 -174133 168325 -174089
rect 168369 -174133 168425 -174089
rect 168469 -174133 168525 -174089
rect 168569 -174133 168625 -174089
rect 168669 -174133 168725 -174089
rect 168769 -174133 168825 -174089
rect 168869 -174133 168925 -174089
rect 168969 -174133 169025 -174089
rect 169069 -174133 169525 -174089
rect 169569 -174133 169625 -174089
rect 169669 -174133 169725 -174089
rect 169769 -174133 169825 -174089
rect 169869 -174133 169925 -174089
rect 169969 -174133 170025 -174089
rect 170069 -174133 170125 -174089
rect 170169 -174133 170225 -174089
rect 170269 -174133 170325 -174089
rect 170369 -174133 170425 -174089
rect 170469 -174133 170525 -174089
rect 170569 -174133 170625 -174089
rect 170669 -174133 170725 -174089
rect 170769 -174133 170825 -174089
rect 170869 -174133 170925 -174089
rect 170969 -174133 171025 -174089
rect 171069 -174133 171525 -174089
rect 171569 -174133 171625 -174089
rect 171669 -174133 171725 -174089
rect 171769 -174133 171825 -174089
rect 171869 -174133 171925 -174089
rect 171969 -174133 172025 -174089
rect 172069 -174133 172125 -174089
rect 172169 -174133 172225 -174089
rect 172269 -174133 172325 -174089
rect 172369 -174133 172425 -174089
rect 172469 -174133 172525 -174089
rect 172569 -174133 172625 -174089
rect 172669 -174133 172725 -174089
rect 172769 -174133 172825 -174089
rect 172869 -174133 172925 -174089
rect 172969 -174133 173025 -174089
rect 173069 -174133 192404 -174089
rect 162407 -174189 192404 -174133
rect 162407 -174233 165525 -174189
rect 165569 -174233 165625 -174189
rect 165669 -174233 165725 -174189
rect 165769 -174233 165825 -174189
rect 165869 -174233 165925 -174189
rect 165969 -174233 166025 -174189
rect 166069 -174233 166125 -174189
rect 166169 -174233 166225 -174189
rect 166269 -174233 166325 -174189
rect 166369 -174233 166425 -174189
rect 166469 -174233 166525 -174189
rect 166569 -174233 166625 -174189
rect 166669 -174233 166725 -174189
rect 166769 -174233 166825 -174189
rect 166869 -174233 166925 -174189
rect 166969 -174233 167025 -174189
rect 167069 -174233 167525 -174189
rect 167569 -174233 167625 -174189
rect 167669 -174233 167725 -174189
rect 167769 -174233 167825 -174189
rect 167869 -174233 167925 -174189
rect 167969 -174233 168025 -174189
rect 168069 -174233 168125 -174189
rect 168169 -174233 168225 -174189
rect 168269 -174233 168325 -174189
rect 168369 -174233 168425 -174189
rect 168469 -174233 168525 -174189
rect 168569 -174233 168625 -174189
rect 168669 -174233 168725 -174189
rect 168769 -174233 168825 -174189
rect 168869 -174233 168925 -174189
rect 168969 -174233 169025 -174189
rect 169069 -174233 169525 -174189
rect 169569 -174233 169625 -174189
rect 169669 -174233 169725 -174189
rect 169769 -174233 169825 -174189
rect 169869 -174233 169925 -174189
rect 169969 -174233 170025 -174189
rect 170069 -174233 170125 -174189
rect 170169 -174233 170225 -174189
rect 170269 -174233 170325 -174189
rect 170369 -174233 170425 -174189
rect 170469 -174233 170525 -174189
rect 170569 -174233 170625 -174189
rect 170669 -174233 170725 -174189
rect 170769 -174233 170825 -174189
rect 170869 -174233 170925 -174189
rect 170969 -174233 171025 -174189
rect 171069 -174233 171525 -174189
rect 171569 -174233 171625 -174189
rect 171669 -174233 171725 -174189
rect 171769 -174233 171825 -174189
rect 171869 -174233 171925 -174189
rect 171969 -174233 172025 -174189
rect 172069 -174233 172125 -174189
rect 172169 -174233 172225 -174189
rect 172269 -174233 172325 -174189
rect 172369 -174233 172425 -174189
rect 172469 -174233 172525 -174189
rect 172569 -174233 172625 -174189
rect 172669 -174233 172725 -174189
rect 172769 -174233 172825 -174189
rect 172869 -174233 172925 -174189
rect 172969 -174233 173025 -174189
rect 173069 -174233 192404 -174189
rect 162407 -174289 192404 -174233
rect 162407 -174333 165525 -174289
rect 165569 -174333 165625 -174289
rect 165669 -174333 165725 -174289
rect 165769 -174333 165825 -174289
rect 165869 -174333 165925 -174289
rect 165969 -174333 166025 -174289
rect 166069 -174333 166125 -174289
rect 166169 -174333 166225 -174289
rect 166269 -174333 166325 -174289
rect 166369 -174333 166425 -174289
rect 166469 -174333 166525 -174289
rect 166569 -174333 166625 -174289
rect 166669 -174333 166725 -174289
rect 166769 -174333 166825 -174289
rect 166869 -174333 166925 -174289
rect 166969 -174333 167025 -174289
rect 167069 -174333 167525 -174289
rect 167569 -174333 167625 -174289
rect 167669 -174333 167725 -174289
rect 167769 -174333 167825 -174289
rect 167869 -174333 167925 -174289
rect 167969 -174333 168025 -174289
rect 168069 -174333 168125 -174289
rect 168169 -174333 168225 -174289
rect 168269 -174333 168325 -174289
rect 168369 -174333 168425 -174289
rect 168469 -174333 168525 -174289
rect 168569 -174333 168625 -174289
rect 168669 -174333 168725 -174289
rect 168769 -174333 168825 -174289
rect 168869 -174333 168925 -174289
rect 168969 -174333 169025 -174289
rect 169069 -174333 169525 -174289
rect 169569 -174333 169625 -174289
rect 169669 -174333 169725 -174289
rect 169769 -174333 169825 -174289
rect 169869 -174333 169925 -174289
rect 169969 -174333 170025 -174289
rect 170069 -174333 170125 -174289
rect 170169 -174333 170225 -174289
rect 170269 -174333 170325 -174289
rect 170369 -174333 170425 -174289
rect 170469 -174333 170525 -174289
rect 170569 -174333 170625 -174289
rect 170669 -174333 170725 -174289
rect 170769 -174333 170825 -174289
rect 170869 -174333 170925 -174289
rect 170969 -174333 171025 -174289
rect 171069 -174333 171525 -174289
rect 171569 -174333 171625 -174289
rect 171669 -174333 171725 -174289
rect 171769 -174333 171825 -174289
rect 171869 -174333 171925 -174289
rect 171969 -174333 172025 -174289
rect 172069 -174333 172125 -174289
rect 172169 -174333 172225 -174289
rect 172269 -174333 172325 -174289
rect 172369 -174333 172425 -174289
rect 172469 -174333 172525 -174289
rect 172569 -174333 172625 -174289
rect 172669 -174333 172725 -174289
rect 172769 -174333 172825 -174289
rect 172869 -174333 172925 -174289
rect 172969 -174333 173025 -174289
rect 173069 -174333 192404 -174289
rect 162407 -174389 192404 -174333
rect 162407 -174433 165525 -174389
rect 165569 -174433 165625 -174389
rect 165669 -174433 165725 -174389
rect 165769 -174433 165825 -174389
rect 165869 -174433 165925 -174389
rect 165969 -174433 166025 -174389
rect 166069 -174433 166125 -174389
rect 166169 -174433 166225 -174389
rect 166269 -174433 166325 -174389
rect 166369 -174433 166425 -174389
rect 166469 -174433 166525 -174389
rect 166569 -174433 166625 -174389
rect 166669 -174433 166725 -174389
rect 166769 -174433 166825 -174389
rect 166869 -174433 166925 -174389
rect 166969 -174433 167025 -174389
rect 167069 -174433 167525 -174389
rect 167569 -174433 167625 -174389
rect 167669 -174433 167725 -174389
rect 167769 -174433 167825 -174389
rect 167869 -174433 167925 -174389
rect 167969 -174433 168025 -174389
rect 168069 -174433 168125 -174389
rect 168169 -174433 168225 -174389
rect 168269 -174433 168325 -174389
rect 168369 -174433 168425 -174389
rect 168469 -174433 168525 -174389
rect 168569 -174433 168625 -174389
rect 168669 -174433 168725 -174389
rect 168769 -174433 168825 -174389
rect 168869 -174433 168925 -174389
rect 168969 -174433 169025 -174389
rect 169069 -174433 169525 -174389
rect 169569 -174433 169625 -174389
rect 169669 -174433 169725 -174389
rect 169769 -174433 169825 -174389
rect 169869 -174433 169925 -174389
rect 169969 -174433 170025 -174389
rect 170069 -174433 170125 -174389
rect 170169 -174433 170225 -174389
rect 170269 -174433 170325 -174389
rect 170369 -174433 170425 -174389
rect 170469 -174433 170525 -174389
rect 170569 -174433 170625 -174389
rect 170669 -174433 170725 -174389
rect 170769 -174433 170825 -174389
rect 170869 -174433 170925 -174389
rect 170969 -174433 171025 -174389
rect 171069 -174433 171525 -174389
rect 171569 -174433 171625 -174389
rect 171669 -174433 171725 -174389
rect 171769 -174433 171825 -174389
rect 171869 -174433 171925 -174389
rect 171969 -174433 172025 -174389
rect 172069 -174433 172125 -174389
rect 172169 -174433 172225 -174389
rect 172269 -174433 172325 -174389
rect 172369 -174433 172425 -174389
rect 172469 -174433 172525 -174389
rect 172569 -174433 172625 -174389
rect 172669 -174433 172725 -174389
rect 172769 -174433 172825 -174389
rect 172869 -174433 172925 -174389
rect 172969 -174433 173025 -174389
rect 173069 -174433 192404 -174389
rect 162407 -174489 192404 -174433
rect 162407 -174533 165525 -174489
rect 165569 -174533 165625 -174489
rect 165669 -174533 165725 -174489
rect 165769 -174533 165825 -174489
rect 165869 -174533 165925 -174489
rect 165969 -174533 166025 -174489
rect 166069 -174533 166125 -174489
rect 166169 -174533 166225 -174489
rect 166269 -174533 166325 -174489
rect 166369 -174533 166425 -174489
rect 166469 -174533 166525 -174489
rect 166569 -174533 166625 -174489
rect 166669 -174533 166725 -174489
rect 166769 -174533 166825 -174489
rect 166869 -174533 166925 -174489
rect 166969 -174533 167025 -174489
rect 167069 -174533 167525 -174489
rect 167569 -174533 167625 -174489
rect 167669 -174533 167725 -174489
rect 167769 -174533 167825 -174489
rect 167869 -174533 167925 -174489
rect 167969 -174533 168025 -174489
rect 168069 -174533 168125 -174489
rect 168169 -174533 168225 -174489
rect 168269 -174533 168325 -174489
rect 168369 -174533 168425 -174489
rect 168469 -174533 168525 -174489
rect 168569 -174533 168625 -174489
rect 168669 -174533 168725 -174489
rect 168769 -174533 168825 -174489
rect 168869 -174533 168925 -174489
rect 168969 -174533 169025 -174489
rect 169069 -174533 169525 -174489
rect 169569 -174533 169625 -174489
rect 169669 -174533 169725 -174489
rect 169769 -174533 169825 -174489
rect 169869 -174533 169925 -174489
rect 169969 -174533 170025 -174489
rect 170069 -174533 170125 -174489
rect 170169 -174533 170225 -174489
rect 170269 -174533 170325 -174489
rect 170369 -174533 170425 -174489
rect 170469 -174533 170525 -174489
rect 170569 -174533 170625 -174489
rect 170669 -174533 170725 -174489
rect 170769 -174533 170825 -174489
rect 170869 -174533 170925 -174489
rect 170969 -174533 171025 -174489
rect 171069 -174533 171525 -174489
rect 171569 -174533 171625 -174489
rect 171669 -174533 171725 -174489
rect 171769 -174533 171825 -174489
rect 171869 -174533 171925 -174489
rect 171969 -174533 172025 -174489
rect 172069 -174533 172125 -174489
rect 172169 -174533 172225 -174489
rect 172269 -174533 172325 -174489
rect 172369 -174533 172425 -174489
rect 172469 -174533 172525 -174489
rect 172569 -174533 172625 -174489
rect 172669 -174533 172725 -174489
rect 172769 -174533 172825 -174489
rect 172869 -174533 172925 -174489
rect 172969 -174533 173025 -174489
rect 173069 -174533 192404 -174489
rect 162407 -175575 192404 -174533
rect 188605 -176154 192404 -175575
<< via2 >>
rect 179458 9144 180057 9674
rect 122315 2353 123454 3016
rect 190005 6200 191144 6863
<< mimcap >>
rect 113625 31171 133625 31743
rect 113625 30875 114357 31171
rect 114653 30875 115117 31171
rect 115413 30875 115877 31171
rect 116173 30875 116637 31171
rect 116933 30875 117397 31171
rect 117693 30875 118157 31171
rect 118453 30875 118917 31171
rect 119213 30875 119677 31171
rect 119973 30875 120437 31171
rect 120733 30875 121197 31171
rect 121493 30875 121957 31171
rect 122253 30875 122717 31171
rect 123013 30875 123477 31171
rect 123773 30875 124237 31171
rect 124533 30875 124997 31171
rect 125293 30875 125757 31171
rect 126053 30875 126517 31171
rect 126813 30875 127277 31171
rect 127573 30875 128037 31171
rect 128333 30875 128797 31171
rect 129093 30875 129557 31171
rect 129853 30875 130317 31171
rect 130613 30875 131077 31171
rect 131373 30875 131837 31171
rect 132133 30875 132597 31171
rect 132893 30875 133625 31171
rect 113625 30411 133625 30875
rect 113625 30115 114357 30411
rect 114653 30115 115117 30411
rect 115413 30115 115877 30411
rect 116173 30115 116637 30411
rect 116933 30115 117397 30411
rect 117693 30115 118157 30411
rect 118453 30115 118917 30411
rect 119213 30115 119677 30411
rect 119973 30115 120437 30411
rect 120733 30115 121197 30411
rect 121493 30115 121957 30411
rect 122253 30115 122717 30411
rect 123013 30115 123477 30411
rect 123773 30115 124237 30411
rect 124533 30115 124997 30411
rect 125293 30115 125757 30411
rect 126053 30115 126517 30411
rect 126813 30115 127277 30411
rect 127573 30115 128037 30411
rect 128333 30115 128797 30411
rect 129093 30115 129557 30411
rect 129853 30115 130317 30411
rect 130613 30115 131077 30411
rect 131373 30115 131837 30411
rect 132133 30115 132597 30411
rect 132893 30115 133625 30411
rect 113625 29651 133625 30115
rect 113625 29355 114357 29651
rect 114653 29355 115117 29651
rect 115413 29355 115877 29651
rect 116173 29355 116637 29651
rect 116933 29355 117397 29651
rect 117693 29355 118157 29651
rect 118453 29355 118917 29651
rect 119213 29355 119677 29651
rect 119973 29355 120437 29651
rect 120733 29355 121197 29651
rect 121493 29355 121957 29651
rect 122253 29355 122717 29651
rect 123013 29355 123477 29651
rect 123773 29355 124237 29651
rect 124533 29355 124997 29651
rect 125293 29355 125757 29651
rect 126053 29355 126517 29651
rect 126813 29355 127277 29651
rect 127573 29355 128037 29651
rect 128333 29355 128797 29651
rect 129093 29355 129557 29651
rect 129853 29355 130317 29651
rect 130613 29355 131077 29651
rect 131373 29355 131837 29651
rect 132133 29355 132597 29651
rect 132893 29355 133625 29651
rect 113625 28891 133625 29355
rect 113625 28595 114357 28891
rect 114653 28595 115117 28891
rect 115413 28595 115877 28891
rect 116173 28595 116637 28891
rect 116933 28595 117397 28891
rect 117693 28595 118157 28891
rect 118453 28595 118917 28891
rect 119213 28595 119677 28891
rect 119973 28595 120437 28891
rect 120733 28595 121197 28891
rect 121493 28595 121957 28891
rect 122253 28595 122717 28891
rect 123013 28595 123477 28891
rect 123773 28595 124237 28891
rect 124533 28595 124997 28891
rect 125293 28595 125757 28891
rect 126053 28595 126517 28891
rect 126813 28595 127277 28891
rect 127573 28595 128037 28891
rect 128333 28595 128797 28891
rect 129093 28595 129557 28891
rect 129853 28595 130317 28891
rect 130613 28595 131077 28891
rect 131373 28595 131837 28891
rect 132133 28595 132597 28891
rect 132893 28595 133625 28891
rect 113625 28131 133625 28595
rect 113625 27835 114357 28131
rect 114653 27835 115117 28131
rect 115413 27835 115877 28131
rect 116173 27835 116637 28131
rect 116933 27835 117397 28131
rect 117693 27835 118157 28131
rect 118453 27835 118917 28131
rect 119213 27835 119677 28131
rect 119973 27835 120437 28131
rect 120733 27835 121197 28131
rect 121493 27835 121957 28131
rect 122253 27835 122717 28131
rect 123013 27835 123477 28131
rect 123773 27835 124237 28131
rect 124533 27835 124997 28131
rect 125293 27835 125757 28131
rect 126053 27835 126517 28131
rect 126813 27835 127277 28131
rect 127573 27835 128037 28131
rect 128333 27835 128797 28131
rect 129093 27835 129557 28131
rect 129853 27835 130317 28131
rect 130613 27835 131077 28131
rect 131373 27835 131837 28131
rect 132133 27835 132597 28131
rect 132893 27835 133625 28131
rect 113625 27371 133625 27835
rect 113625 27075 114357 27371
rect 114653 27075 115117 27371
rect 115413 27075 115877 27371
rect 116173 27075 116637 27371
rect 116933 27075 117397 27371
rect 117693 27075 118157 27371
rect 118453 27075 118917 27371
rect 119213 27075 119677 27371
rect 119973 27075 120437 27371
rect 120733 27075 121197 27371
rect 121493 27075 121957 27371
rect 122253 27075 122717 27371
rect 123013 27075 123477 27371
rect 123773 27075 124237 27371
rect 124533 27075 124997 27371
rect 125293 27075 125757 27371
rect 126053 27075 126517 27371
rect 126813 27075 127277 27371
rect 127573 27075 128037 27371
rect 128333 27075 128797 27371
rect 129093 27075 129557 27371
rect 129853 27075 130317 27371
rect 130613 27075 131077 27371
rect 131373 27075 131837 27371
rect 132133 27075 132597 27371
rect 132893 27075 133625 27371
rect 113625 26611 133625 27075
rect 113625 26315 114357 26611
rect 114653 26315 115117 26611
rect 115413 26315 115877 26611
rect 116173 26315 116637 26611
rect 116933 26315 117397 26611
rect 117693 26315 118157 26611
rect 118453 26315 118917 26611
rect 119213 26315 119677 26611
rect 119973 26315 120437 26611
rect 120733 26315 121197 26611
rect 121493 26315 121957 26611
rect 122253 26315 122717 26611
rect 123013 26315 123477 26611
rect 123773 26315 124237 26611
rect 124533 26315 124997 26611
rect 125293 26315 125757 26611
rect 126053 26315 126517 26611
rect 126813 26315 127277 26611
rect 127573 26315 128037 26611
rect 128333 26315 128797 26611
rect 129093 26315 129557 26611
rect 129853 26315 130317 26611
rect 130613 26315 131077 26611
rect 131373 26315 131837 26611
rect 132133 26315 132597 26611
rect 132893 26315 133625 26611
rect 113625 25851 133625 26315
rect 113625 25555 114357 25851
rect 114653 25555 115117 25851
rect 115413 25555 115877 25851
rect 116173 25555 116637 25851
rect 116933 25555 117397 25851
rect 117693 25555 118157 25851
rect 118453 25555 118917 25851
rect 119213 25555 119677 25851
rect 119973 25555 120437 25851
rect 120733 25555 121197 25851
rect 121493 25555 121957 25851
rect 122253 25555 122717 25851
rect 123013 25555 123477 25851
rect 123773 25555 124237 25851
rect 124533 25555 124997 25851
rect 125293 25555 125757 25851
rect 126053 25555 126517 25851
rect 126813 25555 127277 25851
rect 127573 25555 128037 25851
rect 128333 25555 128797 25851
rect 129093 25555 129557 25851
rect 129853 25555 130317 25851
rect 130613 25555 131077 25851
rect 131373 25555 131837 25851
rect 132133 25555 132597 25851
rect 132893 25555 133625 25851
rect 113625 25091 133625 25555
rect 113625 24795 114357 25091
rect 114653 24795 115117 25091
rect 115413 24795 115877 25091
rect 116173 24795 116637 25091
rect 116933 24795 117397 25091
rect 117693 24795 118157 25091
rect 118453 24795 118917 25091
rect 119213 24795 119677 25091
rect 119973 24795 120437 25091
rect 120733 24795 121197 25091
rect 121493 24795 121957 25091
rect 122253 24795 122717 25091
rect 123013 24795 123477 25091
rect 123773 24795 124237 25091
rect 124533 24795 124997 25091
rect 125293 24795 125757 25091
rect 126053 24795 126517 25091
rect 126813 24795 127277 25091
rect 127573 24795 128037 25091
rect 128333 24795 128797 25091
rect 129093 24795 129557 25091
rect 129853 24795 130317 25091
rect 130613 24795 131077 25091
rect 131373 24795 131837 25091
rect 132133 24795 132597 25091
rect 132893 24795 133625 25091
rect 113625 24331 133625 24795
rect 113625 24035 114357 24331
rect 114653 24035 115117 24331
rect 115413 24035 115877 24331
rect 116173 24035 116637 24331
rect 116933 24035 117397 24331
rect 117693 24035 118157 24331
rect 118453 24035 118917 24331
rect 119213 24035 119677 24331
rect 119973 24035 120437 24331
rect 120733 24035 121197 24331
rect 121493 24035 121957 24331
rect 122253 24035 122717 24331
rect 123013 24035 123477 24331
rect 123773 24035 124237 24331
rect 124533 24035 124997 24331
rect 125293 24035 125757 24331
rect 126053 24035 126517 24331
rect 126813 24035 127277 24331
rect 127573 24035 128037 24331
rect 128333 24035 128797 24331
rect 129093 24035 129557 24331
rect 129853 24035 130317 24331
rect 130613 24035 131077 24331
rect 131373 24035 131837 24331
rect 132133 24035 132597 24331
rect 132893 24035 133625 24331
rect 113625 23571 133625 24035
rect 113625 23275 114357 23571
rect 114653 23275 115117 23571
rect 115413 23275 115877 23571
rect 116173 23275 116637 23571
rect 116933 23275 117397 23571
rect 117693 23275 118157 23571
rect 118453 23275 118917 23571
rect 119213 23275 119677 23571
rect 119973 23275 120437 23571
rect 120733 23275 121197 23571
rect 121493 23275 121957 23571
rect 122253 23275 122717 23571
rect 123013 23275 123477 23571
rect 123773 23275 124237 23571
rect 124533 23275 124997 23571
rect 125293 23275 125757 23571
rect 126053 23275 126517 23571
rect 126813 23275 127277 23571
rect 127573 23275 128037 23571
rect 128333 23275 128797 23571
rect 129093 23275 129557 23571
rect 129853 23275 130317 23571
rect 130613 23275 131077 23571
rect 131373 23275 131837 23571
rect 132133 23275 132597 23571
rect 132893 23275 133625 23571
rect 113625 22811 133625 23275
rect 113625 22515 114357 22811
rect 114653 22515 115117 22811
rect 115413 22515 115877 22811
rect 116173 22515 116637 22811
rect 116933 22515 117397 22811
rect 117693 22515 118157 22811
rect 118453 22515 118917 22811
rect 119213 22515 119677 22811
rect 119973 22515 120437 22811
rect 120733 22515 121197 22811
rect 121493 22515 121957 22811
rect 122253 22515 122717 22811
rect 123013 22515 123477 22811
rect 123773 22515 124237 22811
rect 124533 22515 124997 22811
rect 125293 22515 125757 22811
rect 126053 22515 126517 22811
rect 126813 22515 127277 22811
rect 127573 22515 128037 22811
rect 128333 22515 128797 22811
rect 129093 22515 129557 22811
rect 129853 22515 130317 22811
rect 130613 22515 131077 22811
rect 131373 22515 131837 22811
rect 132133 22515 132597 22811
rect 132893 22515 133625 22811
rect 113625 22051 133625 22515
rect 113625 21755 114357 22051
rect 114653 21755 115117 22051
rect 115413 21755 115877 22051
rect 116173 21755 116637 22051
rect 116933 21755 117397 22051
rect 117693 21755 118157 22051
rect 118453 21755 118917 22051
rect 119213 21755 119677 22051
rect 119973 21755 120437 22051
rect 120733 21755 121197 22051
rect 121493 21755 121957 22051
rect 122253 21755 122717 22051
rect 123013 21755 123477 22051
rect 123773 21755 124237 22051
rect 124533 21755 124997 22051
rect 125293 21755 125757 22051
rect 126053 21755 126517 22051
rect 126813 21755 127277 22051
rect 127573 21755 128037 22051
rect 128333 21755 128797 22051
rect 129093 21755 129557 22051
rect 129853 21755 130317 22051
rect 130613 21755 131077 22051
rect 131373 21755 131837 22051
rect 132133 21755 132597 22051
rect 132893 21755 133625 22051
rect 113625 21291 133625 21755
rect 113625 20995 114357 21291
rect 114653 20995 115117 21291
rect 115413 20995 115877 21291
rect 116173 20995 116637 21291
rect 116933 20995 117397 21291
rect 117693 20995 118157 21291
rect 118453 20995 118917 21291
rect 119213 20995 119677 21291
rect 119973 20995 120437 21291
rect 120733 20995 121197 21291
rect 121493 20995 121957 21291
rect 122253 20995 122717 21291
rect 123013 20995 123477 21291
rect 123773 20995 124237 21291
rect 124533 20995 124997 21291
rect 125293 20995 125757 21291
rect 126053 20995 126517 21291
rect 126813 20995 127277 21291
rect 127573 20995 128037 21291
rect 128333 20995 128797 21291
rect 129093 20995 129557 21291
rect 129853 20995 130317 21291
rect 130613 20995 131077 21291
rect 131373 20995 131837 21291
rect 132133 20995 132597 21291
rect 132893 20995 133625 21291
rect 113625 20531 133625 20995
rect 113625 20235 114357 20531
rect 114653 20235 115117 20531
rect 115413 20235 115877 20531
rect 116173 20235 116637 20531
rect 116933 20235 117397 20531
rect 117693 20235 118157 20531
rect 118453 20235 118917 20531
rect 119213 20235 119677 20531
rect 119973 20235 120437 20531
rect 120733 20235 121197 20531
rect 121493 20235 121957 20531
rect 122253 20235 122717 20531
rect 123013 20235 123477 20531
rect 123773 20235 124237 20531
rect 124533 20235 124997 20531
rect 125293 20235 125757 20531
rect 126053 20235 126517 20531
rect 126813 20235 127277 20531
rect 127573 20235 128037 20531
rect 128333 20235 128797 20531
rect 129093 20235 129557 20531
rect 129853 20235 130317 20531
rect 130613 20235 131077 20531
rect 131373 20235 131837 20531
rect 132133 20235 132597 20531
rect 132893 20235 133625 20531
rect 113625 19771 133625 20235
rect 113625 19475 114357 19771
rect 114653 19475 115117 19771
rect 115413 19475 115877 19771
rect 116173 19475 116637 19771
rect 116933 19475 117397 19771
rect 117693 19475 118157 19771
rect 118453 19475 118917 19771
rect 119213 19475 119677 19771
rect 119973 19475 120437 19771
rect 120733 19475 121197 19771
rect 121493 19475 121957 19771
rect 122253 19475 122717 19771
rect 123013 19475 123477 19771
rect 123773 19475 124237 19771
rect 124533 19475 124997 19771
rect 125293 19475 125757 19771
rect 126053 19475 126517 19771
rect 126813 19475 127277 19771
rect 127573 19475 128037 19771
rect 128333 19475 128797 19771
rect 129093 19475 129557 19771
rect 129853 19475 130317 19771
rect 130613 19475 131077 19771
rect 131373 19475 131837 19771
rect 132133 19475 132597 19771
rect 132893 19475 133625 19771
rect 113625 19011 133625 19475
rect 113625 18715 114357 19011
rect 114653 18715 115117 19011
rect 115413 18715 115877 19011
rect 116173 18715 116637 19011
rect 116933 18715 117397 19011
rect 117693 18715 118157 19011
rect 118453 18715 118917 19011
rect 119213 18715 119677 19011
rect 119973 18715 120437 19011
rect 120733 18715 121197 19011
rect 121493 18715 121957 19011
rect 122253 18715 122717 19011
rect 123013 18715 123477 19011
rect 123773 18715 124237 19011
rect 124533 18715 124997 19011
rect 125293 18715 125757 19011
rect 126053 18715 126517 19011
rect 126813 18715 127277 19011
rect 127573 18715 128037 19011
rect 128333 18715 128797 19011
rect 129093 18715 129557 19011
rect 129853 18715 130317 19011
rect 130613 18715 131077 19011
rect 131373 18715 131837 19011
rect 132133 18715 132597 19011
rect 132893 18715 133625 19011
rect 113625 18251 133625 18715
rect 113625 17955 114357 18251
rect 114653 17955 115117 18251
rect 115413 17955 115877 18251
rect 116173 17955 116637 18251
rect 116933 17955 117397 18251
rect 117693 17955 118157 18251
rect 118453 17955 118917 18251
rect 119213 17955 119677 18251
rect 119973 17955 120437 18251
rect 120733 17955 121197 18251
rect 121493 17955 121957 18251
rect 122253 17955 122717 18251
rect 123013 17955 123477 18251
rect 123773 17955 124237 18251
rect 124533 17955 124997 18251
rect 125293 17955 125757 18251
rect 126053 17955 126517 18251
rect 126813 17955 127277 18251
rect 127573 17955 128037 18251
rect 128333 17955 128797 18251
rect 129093 17955 129557 18251
rect 129853 17955 130317 18251
rect 130613 17955 131077 18251
rect 131373 17955 131837 18251
rect 132133 17955 132597 18251
rect 132893 17955 133625 18251
rect 113625 17491 133625 17955
rect 113625 17195 114357 17491
rect 114653 17195 115117 17491
rect 115413 17195 115877 17491
rect 116173 17195 116637 17491
rect 116933 17195 117397 17491
rect 117693 17195 118157 17491
rect 118453 17195 118917 17491
rect 119213 17195 119677 17491
rect 119973 17195 120437 17491
rect 120733 17195 121197 17491
rect 121493 17195 121957 17491
rect 122253 17195 122717 17491
rect 123013 17195 123477 17491
rect 123773 17195 124237 17491
rect 124533 17195 124997 17491
rect 125293 17195 125757 17491
rect 126053 17195 126517 17491
rect 126813 17195 127277 17491
rect 127573 17195 128037 17491
rect 128333 17195 128797 17491
rect 129093 17195 129557 17491
rect 129853 17195 130317 17491
rect 130613 17195 131077 17491
rect 131373 17195 131837 17491
rect 132133 17195 132597 17491
rect 132893 17195 133625 17491
rect 113625 16731 133625 17195
rect 113625 16435 114357 16731
rect 114653 16435 115117 16731
rect 115413 16435 115877 16731
rect 116173 16435 116637 16731
rect 116933 16435 117397 16731
rect 117693 16435 118157 16731
rect 118453 16435 118917 16731
rect 119213 16435 119677 16731
rect 119973 16435 120437 16731
rect 120733 16435 121197 16731
rect 121493 16435 121957 16731
rect 122253 16435 122717 16731
rect 123013 16435 123477 16731
rect 123773 16435 124237 16731
rect 124533 16435 124997 16731
rect 125293 16435 125757 16731
rect 126053 16435 126517 16731
rect 126813 16435 127277 16731
rect 127573 16435 128037 16731
rect 128333 16435 128797 16731
rect 129093 16435 129557 16731
rect 129853 16435 130317 16731
rect 130613 16435 131077 16731
rect 131373 16435 131837 16731
rect 132133 16435 132597 16731
rect 132893 16435 133625 16731
rect 113625 15971 133625 16435
rect 113625 15675 114357 15971
rect 114653 15675 115117 15971
rect 115413 15675 115877 15971
rect 116173 15675 116637 15971
rect 116933 15675 117397 15971
rect 117693 15675 118157 15971
rect 118453 15675 118917 15971
rect 119213 15675 119677 15971
rect 119973 15675 120437 15971
rect 120733 15675 121197 15971
rect 121493 15675 121957 15971
rect 122253 15675 122717 15971
rect 123013 15675 123477 15971
rect 123773 15675 124237 15971
rect 124533 15675 124997 15971
rect 125293 15675 125757 15971
rect 126053 15675 126517 15971
rect 126813 15675 127277 15971
rect 127573 15675 128037 15971
rect 128333 15675 128797 15971
rect 129093 15675 129557 15971
rect 129853 15675 130317 15971
rect 130613 15675 131077 15971
rect 131373 15675 131837 15971
rect 132133 15675 132597 15971
rect 132893 15675 133625 15971
rect 113625 15211 133625 15675
rect 113625 14915 114357 15211
rect 114653 14915 115117 15211
rect 115413 14915 115877 15211
rect 116173 14915 116637 15211
rect 116933 14915 117397 15211
rect 117693 14915 118157 15211
rect 118453 14915 118917 15211
rect 119213 14915 119677 15211
rect 119973 14915 120437 15211
rect 120733 14915 121197 15211
rect 121493 14915 121957 15211
rect 122253 14915 122717 15211
rect 123013 14915 123477 15211
rect 123773 14915 124237 15211
rect 124533 14915 124997 15211
rect 125293 14915 125757 15211
rect 126053 14915 126517 15211
rect 126813 14915 127277 15211
rect 127573 14915 128037 15211
rect 128333 14915 128797 15211
rect 129093 14915 129557 15211
rect 129853 14915 130317 15211
rect 130613 14915 131077 15211
rect 131373 14915 131837 15211
rect 132133 14915 132597 15211
rect 132893 14915 133625 15211
rect 113625 14451 133625 14915
rect 113625 14155 114357 14451
rect 114653 14155 115117 14451
rect 115413 14155 115877 14451
rect 116173 14155 116637 14451
rect 116933 14155 117397 14451
rect 117693 14155 118157 14451
rect 118453 14155 118917 14451
rect 119213 14155 119677 14451
rect 119973 14155 120437 14451
rect 120733 14155 121197 14451
rect 121493 14155 121957 14451
rect 122253 14155 122717 14451
rect 123013 14155 123477 14451
rect 123773 14155 124237 14451
rect 124533 14155 124997 14451
rect 125293 14155 125757 14451
rect 126053 14155 126517 14451
rect 126813 14155 127277 14451
rect 127573 14155 128037 14451
rect 128333 14155 128797 14451
rect 129093 14155 129557 14451
rect 129853 14155 130317 14451
rect 130613 14155 131077 14451
rect 131373 14155 131837 14451
rect 132133 14155 132597 14451
rect 132893 14155 133625 14451
rect 113625 13691 133625 14155
rect 113625 13395 114357 13691
rect 114653 13395 115117 13691
rect 115413 13395 115877 13691
rect 116173 13395 116637 13691
rect 116933 13395 117397 13691
rect 117693 13395 118157 13691
rect 118453 13395 118917 13691
rect 119213 13395 119677 13691
rect 119973 13395 120437 13691
rect 120733 13395 121197 13691
rect 121493 13395 121957 13691
rect 122253 13395 122717 13691
rect 123013 13395 123477 13691
rect 123773 13395 124237 13691
rect 124533 13395 124997 13691
rect 125293 13395 125757 13691
rect 126053 13395 126517 13691
rect 126813 13395 127277 13691
rect 127573 13395 128037 13691
rect 128333 13395 128797 13691
rect 129093 13395 129557 13691
rect 129853 13395 130317 13691
rect 130613 13395 131077 13691
rect 131373 13395 131837 13691
rect 132133 13395 132597 13691
rect 132893 13395 133625 13691
rect 113625 12931 133625 13395
rect 113625 12635 114357 12931
rect 114653 12635 115117 12931
rect 115413 12635 115877 12931
rect 116173 12635 116637 12931
rect 116933 12635 117397 12931
rect 117693 12635 118157 12931
rect 118453 12635 118917 12931
rect 119213 12635 119677 12931
rect 119973 12635 120437 12931
rect 120733 12635 121197 12931
rect 121493 12635 121957 12931
rect 122253 12635 122717 12931
rect 123013 12635 123477 12931
rect 123773 12635 124237 12931
rect 124533 12635 124997 12931
rect 125293 12635 125757 12931
rect 126053 12635 126517 12931
rect 126813 12635 127277 12931
rect 127573 12635 128037 12931
rect 128333 12635 128797 12931
rect 129093 12635 129557 12931
rect 129853 12635 130317 12931
rect 130613 12635 131077 12931
rect 131373 12635 131837 12931
rect 132133 12635 132597 12931
rect 132893 12635 133625 12931
rect 113625 12171 133625 12635
rect 113625 11875 114357 12171
rect 114653 11875 115117 12171
rect 115413 11875 115877 12171
rect 116173 11875 116637 12171
rect 116933 11875 117397 12171
rect 117693 11875 118157 12171
rect 118453 11875 118917 12171
rect 119213 11875 119677 12171
rect 119973 11875 120437 12171
rect 120733 11875 121197 12171
rect 121493 11875 121957 12171
rect 122253 11875 122717 12171
rect 123013 11875 123477 12171
rect 123773 11875 124237 12171
rect 124533 11875 124997 12171
rect 125293 11875 125757 12171
rect 126053 11875 126517 12171
rect 126813 11875 127277 12171
rect 127573 11875 128037 12171
rect 128333 11875 128797 12171
rect 129093 11875 129557 12171
rect 129853 11875 130317 12171
rect 130613 11875 131077 12171
rect 131373 11875 131837 12171
rect 132133 11875 132597 12171
rect 132893 11875 133625 12171
rect 113625 11411 133625 11875
rect 113625 11115 114357 11411
rect 114653 11115 115117 11411
rect 115413 11115 115877 11411
rect 116173 11115 116637 11411
rect 116933 11115 117397 11411
rect 117693 11115 118157 11411
rect 118453 11115 118917 11411
rect 119213 11115 119677 11411
rect 119973 11115 120437 11411
rect 120733 11115 121197 11411
rect 121493 11115 121957 11411
rect 122253 11115 122717 11411
rect 123013 11115 123477 11411
rect 123773 11115 124237 11411
rect 124533 11115 124997 11411
rect 125293 11115 125757 11411
rect 126053 11115 126517 11411
rect 126813 11115 127277 11411
rect 127573 11115 128037 11411
rect 128333 11115 128797 11411
rect 129093 11115 129557 11411
rect 129853 11115 130317 11411
rect 130613 11115 131077 11411
rect 131373 11115 131837 11411
rect 132133 11115 132597 11411
rect 132893 11115 133625 11411
rect 113625 10651 133625 11115
rect 113625 10355 114357 10651
rect 114653 10355 115117 10651
rect 115413 10355 115877 10651
rect 116173 10355 116637 10651
rect 116933 10355 117397 10651
rect 117693 10355 118157 10651
rect 118453 10355 118917 10651
rect 119213 10355 119677 10651
rect 119973 10355 120437 10651
rect 120733 10355 121197 10651
rect 121493 10355 121957 10651
rect 122253 10355 122717 10651
rect 123013 10355 123477 10651
rect 123773 10355 124237 10651
rect 124533 10355 124997 10651
rect 125293 10355 125757 10651
rect 126053 10355 126517 10651
rect 126813 10355 127277 10651
rect 127573 10355 128037 10651
rect 128333 10355 128797 10651
rect 129093 10355 129557 10651
rect 129853 10355 130317 10651
rect 130613 10355 131077 10651
rect 131373 10355 131837 10651
rect 132133 10355 132597 10651
rect 132893 10355 133625 10651
rect 113625 9891 133625 10355
rect 113625 9595 114357 9891
rect 114653 9595 115117 9891
rect 115413 9595 115877 9891
rect 116173 9595 116637 9891
rect 116933 9595 117397 9891
rect 117693 9595 118157 9891
rect 118453 9595 118917 9891
rect 119213 9595 119677 9891
rect 119973 9595 120437 9891
rect 120733 9595 121197 9891
rect 121493 9595 121957 9891
rect 122253 9595 122717 9891
rect 123013 9595 123477 9891
rect 123773 9595 124237 9891
rect 124533 9595 124997 9891
rect 125293 9595 125757 9891
rect 126053 9595 126517 9891
rect 126813 9595 127277 9891
rect 127573 9595 128037 9891
rect 128333 9595 128797 9891
rect 129093 9595 129557 9891
rect 129853 9595 130317 9891
rect 130613 9595 131077 9891
rect 131373 9595 131837 9891
rect 132133 9595 132597 9891
rect 132893 9595 133625 9891
rect 113625 9131 133625 9595
rect 113625 8835 114357 9131
rect 114653 8835 115117 9131
rect 115413 8835 115877 9131
rect 116173 8835 116637 9131
rect 116933 8835 117397 9131
rect 117693 8835 118157 9131
rect 118453 8835 118917 9131
rect 119213 8835 119677 9131
rect 119973 8835 120437 9131
rect 120733 8835 121197 9131
rect 121493 8835 121957 9131
rect 122253 8835 122717 9131
rect 123013 8835 123477 9131
rect 123773 8835 124237 9131
rect 124533 8835 124997 9131
rect 125293 8835 125757 9131
rect 126053 8835 126517 9131
rect 126813 8835 127277 9131
rect 127573 8835 128037 9131
rect 128333 8835 128797 9131
rect 129093 8835 129557 9131
rect 129853 8835 130317 9131
rect 130613 8835 131077 9131
rect 131373 8835 131837 9131
rect 132133 8835 132597 9131
rect 132893 8835 133625 9131
rect 113625 8371 133625 8835
rect 113625 8075 114357 8371
rect 114653 8075 115117 8371
rect 115413 8075 115877 8371
rect 116173 8075 116637 8371
rect 116933 8075 117397 8371
rect 117693 8075 118157 8371
rect 118453 8075 118917 8371
rect 119213 8075 119677 8371
rect 119973 8075 120437 8371
rect 120733 8075 121197 8371
rect 121493 8075 121957 8371
rect 122253 8075 122717 8371
rect 123013 8075 123477 8371
rect 123773 8075 124237 8371
rect 124533 8075 124997 8371
rect 125293 8075 125757 8371
rect 126053 8075 126517 8371
rect 126813 8075 127277 8371
rect 127573 8075 128037 8371
rect 128333 8075 128797 8371
rect 129093 8075 129557 8371
rect 129853 8075 130317 8371
rect 130613 8075 131077 8371
rect 131373 8075 131837 8371
rect 132133 8075 132597 8371
rect 132893 8075 133625 8371
rect 113625 7611 133625 8075
rect 113625 7315 114357 7611
rect 114653 7315 115117 7611
rect 115413 7315 115877 7611
rect 116173 7315 116637 7611
rect 116933 7315 117397 7611
rect 117693 7315 118157 7611
rect 118453 7315 118917 7611
rect 119213 7315 119677 7611
rect 119973 7315 120437 7611
rect 120733 7315 121197 7611
rect 121493 7315 121957 7611
rect 122253 7315 122717 7611
rect 123013 7315 123477 7611
rect 123773 7315 124237 7611
rect 124533 7315 124997 7611
rect 125293 7315 125757 7611
rect 126053 7315 126517 7611
rect 126813 7315 127277 7611
rect 127573 7315 128037 7611
rect 128333 7315 128797 7611
rect 129093 7315 129557 7611
rect 129853 7315 130317 7611
rect 130613 7315 131077 7611
rect 131373 7315 131837 7611
rect 132133 7315 132597 7611
rect 132893 7315 133625 7611
rect 113625 6743 133625 7315
rect 135425 31171 155425 31743
rect 135425 30875 136157 31171
rect 136453 30875 136917 31171
rect 137213 30875 137677 31171
rect 137973 30875 138437 31171
rect 138733 30875 139197 31171
rect 139493 30875 139957 31171
rect 140253 30875 140717 31171
rect 141013 30875 141477 31171
rect 141773 30875 142237 31171
rect 142533 30875 142997 31171
rect 143293 30875 143757 31171
rect 144053 30875 144517 31171
rect 144813 30875 145277 31171
rect 145573 30875 146037 31171
rect 146333 30875 146797 31171
rect 147093 30875 147557 31171
rect 147853 30875 148317 31171
rect 148613 30875 149077 31171
rect 149373 30875 149837 31171
rect 150133 30875 150597 31171
rect 150893 30875 151357 31171
rect 151653 30875 152117 31171
rect 152413 30875 152877 31171
rect 153173 30875 153637 31171
rect 153933 30875 154397 31171
rect 154693 30875 155425 31171
rect 135425 30411 155425 30875
rect 135425 30115 136157 30411
rect 136453 30115 136917 30411
rect 137213 30115 137677 30411
rect 137973 30115 138437 30411
rect 138733 30115 139197 30411
rect 139493 30115 139957 30411
rect 140253 30115 140717 30411
rect 141013 30115 141477 30411
rect 141773 30115 142237 30411
rect 142533 30115 142997 30411
rect 143293 30115 143757 30411
rect 144053 30115 144517 30411
rect 144813 30115 145277 30411
rect 145573 30115 146037 30411
rect 146333 30115 146797 30411
rect 147093 30115 147557 30411
rect 147853 30115 148317 30411
rect 148613 30115 149077 30411
rect 149373 30115 149837 30411
rect 150133 30115 150597 30411
rect 150893 30115 151357 30411
rect 151653 30115 152117 30411
rect 152413 30115 152877 30411
rect 153173 30115 153637 30411
rect 153933 30115 154397 30411
rect 154693 30115 155425 30411
rect 135425 29651 155425 30115
rect 135425 29355 136157 29651
rect 136453 29355 136917 29651
rect 137213 29355 137677 29651
rect 137973 29355 138437 29651
rect 138733 29355 139197 29651
rect 139493 29355 139957 29651
rect 140253 29355 140717 29651
rect 141013 29355 141477 29651
rect 141773 29355 142237 29651
rect 142533 29355 142997 29651
rect 143293 29355 143757 29651
rect 144053 29355 144517 29651
rect 144813 29355 145277 29651
rect 145573 29355 146037 29651
rect 146333 29355 146797 29651
rect 147093 29355 147557 29651
rect 147853 29355 148317 29651
rect 148613 29355 149077 29651
rect 149373 29355 149837 29651
rect 150133 29355 150597 29651
rect 150893 29355 151357 29651
rect 151653 29355 152117 29651
rect 152413 29355 152877 29651
rect 153173 29355 153637 29651
rect 153933 29355 154397 29651
rect 154693 29355 155425 29651
rect 135425 28891 155425 29355
rect 135425 28595 136157 28891
rect 136453 28595 136917 28891
rect 137213 28595 137677 28891
rect 137973 28595 138437 28891
rect 138733 28595 139197 28891
rect 139493 28595 139957 28891
rect 140253 28595 140717 28891
rect 141013 28595 141477 28891
rect 141773 28595 142237 28891
rect 142533 28595 142997 28891
rect 143293 28595 143757 28891
rect 144053 28595 144517 28891
rect 144813 28595 145277 28891
rect 145573 28595 146037 28891
rect 146333 28595 146797 28891
rect 147093 28595 147557 28891
rect 147853 28595 148317 28891
rect 148613 28595 149077 28891
rect 149373 28595 149837 28891
rect 150133 28595 150597 28891
rect 150893 28595 151357 28891
rect 151653 28595 152117 28891
rect 152413 28595 152877 28891
rect 153173 28595 153637 28891
rect 153933 28595 154397 28891
rect 154693 28595 155425 28891
rect 135425 28131 155425 28595
rect 135425 27835 136157 28131
rect 136453 27835 136917 28131
rect 137213 27835 137677 28131
rect 137973 27835 138437 28131
rect 138733 27835 139197 28131
rect 139493 27835 139957 28131
rect 140253 27835 140717 28131
rect 141013 27835 141477 28131
rect 141773 27835 142237 28131
rect 142533 27835 142997 28131
rect 143293 27835 143757 28131
rect 144053 27835 144517 28131
rect 144813 27835 145277 28131
rect 145573 27835 146037 28131
rect 146333 27835 146797 28131
rect 147093 27835 147557 28131
rect 147853 27835 148317 28131
rect 148613 27835 149077 28131
rect 149373 27835 149837 28131
rect 150133 27835 150597 28131
rect 150893 27835 151357 28131
rect 151653 27835 152117 28131
rect 152413 27835 152877 28131
rect 153173 27835 153637 28131
rect 153933 27835 154397 28131
rect 154693 27835 155425 28131
rect 135425 27371 155425 27835
rect 135425 27075 136157 27371
rect 136453 27075 136917 27371
rect 137213 27075 137677 27371
rect 137973 27075 138437 27371
rect 138733 27075 139197 27371
rect 139493 27075 139957 27371
rect 140253 27075 140717 27371
rect 141013 27075 141477 27371
rect 141773 27075 142237 27371
rect 142533 27075 142997 27371
rect 143293 27075 143757 27371
rect 144053 27075 144517 27371
rect 144813 27075 145277 27371
rect 145573 27075 146037 27371
rect 146333 27075 146797 27371
rect 147093 27075 147557 27371
rect 147853 27075 148317 27371
rect 148613 27075 149077 27371
rect 149373 27075 149837 27371
rect 150133 27075 150597 27371
rect 150893 27075 151357 27371
rect 151653 27075 152117 27371
rect 152413 27075 152877 27371
rect 153173 27075 153637 27371
rect 153933 27075 154397 27371
rect 154693 27075 155425 27371
rect 135425 26611 155425 27075
rect 135425 26315 136157 26611
rect 136453 26315 136917 26611
rect 137213 26315 137677 26611
rect 137973 26315 138437 26611
rect 138733 26315 139197 26611
rect 139493 26315 139957 26611
rect 140253 26315 140717 26611
rect 141013 26315 141477 26611
rect 141773 26315 142237 26611
rect 142533 26315 142997 26611
rect 143293 26315 143757 26611
rect 144053 26315 144517 26611
rect 144813 26315 145277 26611
rect 145573 26315 146037 26611
rect 146333 26315 146797 26611
rect 147093 26315 147557 26611
rect 147853 26315 148317 26611
rect 148613 26315 149077 26611
rect 149373 26315 149837 26611
rect 150133 26315 150597 26611
rect 150893 26315 151357 26611
rect 151653 26315 152117 26611
rect 152413 26315 152877 26611
rect 153173 26315 153637 26611
rect 153933 26315 154397 26611
rect 154693 26315 155425 26611
rect 135425 25851 155425 26315
rect 135425 25555 136157 25851
rect 136453 25555 136917 25851
rect 137213 25555 137677 25851
rect 137973 25555 138437 25851
rect 138733 25555 139197 25851
rect 139493 25555 139957 25851
rect 140253 25555 140717 25851
rect 141013 25555 141477 25851
rect 141773 25555 142237 25851
rect 142533 25555 142997 25851
rect 143293 25555 143757 25851
rect 144053 25555 144517 25851
rect 144813 25555 145277 25851
rect 145573 25555 146037 25851
rect 146333 25555 146797 25851
rect 147093 25555 147557 25851
rect 147853 25555 148317 25851
rect 148613 25555 149077 25851
rect 149373 25555 149837 25851
rect 150133 25555 150597 25851
rect 150893 25555 151357 25851
rect 151653 25555 152117 25851
rect 152413 25555 152877 25851
rect 153173 25555 153637 25851
rect 153933 25555 154397 25851
rect 154693 25555 155425 25851
rect 135425 25091 155425 25555
rect 135425 24795 136157 25091
rect 136453 24795 136917 25091
rect 137213 24795 137677 25091
rect 137973 24795 138437 25091
rect 138733 24795 139197 25091
rect 139493 24795 139957 25091
rect 140253 24795 140717 25091
rect 141013 24795 141477 25091
rect 141773 24795 142237 25091
rect 142533 24795 142997 25091
rect 143293 24795 143757 25091
rect 144053 24795 144517 25091
rect 144813 24795 145277 25091
rect 145573 24795 146037 25091
rect 146333 24795 146797 25091
rect 147093 24795 147557 25091
rect 147853 24795 148317 25091
rect 148613 24795 149077 25091
rect 149373 24795 149837 25091
rect 150133 24795 150597 25091
rect 150893 24795 151357 25091
rect 151653 24795 152117 25091
rect 152413 24795 152877 25091
rect 153173 24795 153637 25091
rect 153933 24795 154397 25091
rect 154693 24795 155425 25091
rect 135425 24331 155425 24795
rect 135425 24035 136157 24331
rect 136453 24035 136917 24331
rect 137213 24035 137677 24331
rect 137973 24035 138437 24331
rect 138733 24035 139197 24331
rect 139493 24035 139957 24331
rect 140253 24035 140717 24331
rect 141013 24035 141477 24331
rect 141773 24035 142237 24331
rect 142533 24035 142997 24331
rect 143293 24035 143757 24331
rect 144053 24035 144517 24331
rect 144813 24035 145277 24331
rect 145573 24035 146037 24331
rect 146333 24035 146797 24331
rect 147093 24035 147557 24331
rect 147853 24035 148317 24331
rect 148613 24035 149077 24331
rect 149373 24035 149837 24331
rect 150133 24035 150597 24331
rect 150893 24035 151357 24331
rect 151653 24035 152117 24331
rect 152413 24035 152877 24331
rect 153173 24035 153637 24331
rect 153933 24035 154397 24331
rect 154693 24035 155425 24331
rect 135425 23571 155425 24035
rect 135425 23275 136157 23571
rect 136453 23275 136917 23571
rect 137213 23275 137677 23571
rect 137973 23275 138437 23571
rect 138733 23275 139197 23571
rect 139493 23275 139957 23571
rect 140253 23275 140717 23571
rect 141013 23275 141477 23571
rect 141773 23275 142237 23571
rect 142533 23275 142997 23571
rect 143293 23275 143757 23571
rect 144053 23275 144517 23571
rect 144813 23275 145277 23571
rect 145573 23275 146037 23571
rect 146333 23275 146797 23571
rect 147093 23275 147557 23571
rect 147853 23275 148317 23571
rect 148613 23275 149077 23571
rect 149373 23275 149837 23571
rect 150133 23275 150597 23571
rect 150893 23275 151357 23571
rect 151653 23275 152117 23571
rect 152413 23275 152877 23571
rect 153173 23275 153637 23571
rect 153933 23275 154397 23571
rect 154693 23275 155425 23571
rect 135425 22811 155425 23275
rect 135425 22515 136157 22811
rect 136453 22515 136917 22811
rect 137213 22515 137677 22811
rect 137973 22515 138437 22811
rect 138733 22515 139197 22811
rect 139493 22515 139957 22811
rect 140253 22515 140717 22811
rect 141013 22515 141477 22811
rect 141773 22515 142237 22811
rect 142533 22515 142997 22811
rect 143293 22515 143757 22811
rect 144053 22515 144517 22811
rect 144813 22515 145277 22811
rect 145573 22515 146037 22811
rect 146333 22515 146797 22811
rect 147093 22515 147557 22811
rect 147853 22515 148317 22811
rect 148613 22515 149077 22811
rect 149373 22515 149837 22811
rect 150133 22515 150597 22811
rect 150893 22515 151357 22811
rect 151653 22515 152117 22811
rect 152413 22515 152877 22811
rect 153173 22515 153637 22811
rect 153933 22515 154397 22811
rect 154693 22515 155425 22811
rect 135425 22051 155425 22515
rect 135425 21755 136157 22051
rect 136453 21755 136917 22051
rect 137213 21755 137677 22051
rect 137973 21755 138437 22051
rect 138733 21755 139197 22051
rect 139493 21755 139957 22051
rect 140253 21755 140717 22051
rect 141013 21755 141477 22051
rect 141773 21755 142237 22051
rect 142533 21755 142997 22051
rect 143293 21755 143757 22051
rect 144053 21755 144517 22051
rect 144813 21755 145277 22051
rect 145573 21755 146037 22051
rect 146333 21755 146797 22051
rect 147093 21755 147557 22051
rect 147853 21755 148317 22051
rect 148613 21755 149077 22051
rect 149373 21755 149837 22051
rect 150133 21755 150597 22051
rect 150893 21755 151357 22051
rect 151653 21755 152117 22051
rect 152413 21755 152877 22051
rect 153173 21755 153637 22051
rect 153933 21755 154397 22051
rect 154693 21755 155425 22051
rect 135425 21291 155425 21755
rect 135425 20995 136157 21291
rect 136453 20995 136917 21291
rect 137213 20995 137677 21291
rect 137973 20995 138437 21291
rect 138733 20995 139197 21291
rect 139493 20995 139957 21291
rect 140253 20995 140717 21291
rect 141013 20995 141477 21291
rect 141773 20995 142237 21291
rect 142533 20995 142997 21291
rect 143293 20995 143757 21291
rect 144053 20995 144517 21291
rect 144813 20995 145277 21291
rect 145573 20995 146037 21291
rect 146333 20995 146797 21291
rect 147093 20995 147557 21291
rect 147853 20995 148317 21291
rect 148613 20995 149077 21291
rect 149373 20995 149837 21291
rect 150133 20995 150597 21291
rect 150893 20995 151357 21291
rect 151653 20995 152117 21291
rect 152413 20995 152877 21291
rect 153173 20995 153637 21291
rect 153933 20995 154397 21291
rect 154693 20995 155425 21291
rect 135425 20531 155425 20995
rect 135425 20235 136157 20531
rect 136453 20235 136917 20531
rect 137213 20235 137677 20531
rect 137973 20235 138437 20531
rect 138733 20235 139197 20531
rect 139493 20235 139957 20531
rect 140253 20235 140717 20531
rect 141013 20235 141477 20531
rect 141773 20235 142237 20531
rect 142533 20235 142997 20531
rect 143293 20235 143757 20531
rect 144053 20235 144517 20531
rect 144813 20235 145277 20531
rect 145573 20235 146037 20531
rect 146333 20235 146797 20531
rect 147093 20235 147557 20531
rect 147853 20235 148317 20531
rect 148613 20235 149077 20531
rect 149373 20235 149837 20531
rect 150133 20235 150597 20531
rect 150893 20235 151357 20531
rect 151653 20235 152117 20531
rect 152413 20235 152877 20531
rect 153173 20235 153637 20531
rect 153933 20235 154397 20531
rect 154693 20235 155425 20531
rect 135425 19771 155425 20235
rect 135425 19475 136157 19771
rect 136453 19475 136917 19771
rect 137213 19475 137677 19771
rect 137973 19475 138437 19771
rect 138733 19475 139197 19771
rect 139493 19475 139957 19771
rect 140253 19475 140717 19771
rect 141013 19475 141477 19771
rect 141773 19475 142237 19771
rect 142533 19475 142997 19771
rect 143293 19475 143757 19771
rect 144053 19475 144517 19771
rect 144813 19475 145277 19771
rect 145573 19475 146037 19771
rect 146333 19475 146797 19771
rect 147093 19475 147557 19771
rect 147853 19475 148317 19771
rect 148613 19475 149077 19771
rect 149373 19475 149837 19771
rect 150133 19475 150597 19771
rect 150893 19475 151357 19771
rect 151653 19475 152117 19771
rect 152413 19475 152877 19771
rect 153173 19475 153637 19771
rect 153933 19475 154397 19771
rect 154693 19475 155425 19771
rect 135425 19011 155425 19475
rect 135425 18715 136157 19011
rect 136453 18715 136917 19011
rect 137213 18715 137677 19011
rect 137973 18715 138437 19011
rect 138733 18715 139197 19011
rect 139493 18715 139957 19011
rect 140253 18715 140717 19011
rect 141013 18715 141477 19011
rect 141773 18715 142237 19011
rect 142533 18715 142997 19011
rect 143293 18715 143757 19011
rect 144053 18715 144517 19011
rect 144813 18715 145277 19011
rect 145573 18715 146037 19011
rect 146333 18715 146797 19011
rect 147093 18715 147557 19011
rect 147853 18715 148317 19011
rect 148613 18715 149077 19011
rect 149373 18715 149837 19011
rect 150133 18715 150597 19011
rect 150893 18715 151357 19011
rect 151653 18715 152117 19011
rect 152413 18715 152877 19011
rect 153173 18715 153637 19011
rect 153933 18715 154397 19011
rect 154693 18715 155425 19011
rect 135425 18251 155425 18715
rect 135425 17955 136157 18251
rect 136453 17955 136917 18251
rect 137213 17955 137677 18251
rect 137973 17955 138437 18251
rect 138733 17955 139197 18251
rect 139493 17955 139957 18251
rect 140253 17955 140717 18251
rect 141013 17955 141477 18251
rect 141773 17955 142237 18251
rect 142533 17955 142997 18251
rect 143293 17955 143757 18251
rect 144053 17955 144517 18251
rect 144813 17955 145277 18251
rect 145573 17955 146037 18251
rect 146333 17955 146797 18251
rect 147093 17955 147557 18251
rect 147853 17955 148317 18251
rect 148613 17955 149077 18251
rect 149373 17955 149837 18251
rect 150133 17955 150597 18251
rect 150893 17955 151357 18251
rect 151653 17955 152117 18251
rect 152413 17955 152877 18251
rect 153173 17955 153637 18251
rect 153933 17955 154397 18251
rect 154693 17955 155425 18251
rect 135425 17491 155425 17955
rect 135425 17195 136157 17491
rect 136453 17195 136917 17491
rect 137213 17195 137677 17491
rect 137973 17195 138437 17491
rect 138733 17195 139197 17491
rect 139493 17195 139957 17491
rect 140253 17195 140717 17491
rect 141013 17195 141477 17491
rect 141773 17195 142237 17491
rect 142533 17195 142997 17491
rect 143293 17195 143757 17491
rect 144053 17195 144517 17491
rect 144813 17195 145277 17491
rect 145573 17195 146037 17491
rect 146333 17195 146797 17491
rect 147093 17195 147557 17491
rect 147853 17195 148317 17491
rect 148613 17195 149077 17491
rect 149373 17195 149837 17491
rect 150133 17195 150597 17491
rect 150893 17195 151357 17491
rect 151653 17195 152117 17491
rect 152413 17195 152877 17491
rect 153173 17195 153637 17491
rect 153933 17195 154397 17491
rect 154693 17195 155425 17491
rect 135425 16731 155425 17195
rect 135425 16435 136157 16731
rect 136453 16435 136917 16731
rect 137213 16435 137677 16731
rect 137973 16435 138437 16731
rect 138733 16435 139197 16731
rect 139493 16435 139957 16731
rect 140253 16435 140717 16731
rect 141013 16435 141477 16731
rect 141773 16435 142237 16731
rect 142533 16435 142997 16731
rect 143293 16435 143757 16731
rect 144053 16435 144517 16731
rect 144813 16435 145277 16731
rect 145573 16435 146037 16731
rect 146333 16435 146797 16731
rect 147093 16435 147557 16731
rect 147853 16435 148317 16731
rect 148613 16435 149077 16731
rect 149373 16435 149837 16731
rect 150133 16435 150597 16731
rect 150893 16435 151357 16731
rect 151653 16435 152117 16731
rect 152413 16435 152877 16731
rect 153173 16435 153637 16731
rect 153933 16435 154397 16731
rect 154693 16435 155425 16731
rect 135425 15971 155425 16435
rect 135425 15675 136157 15971
rect 136453 15675 136917 15971
rect 137213 15675 137677 15971
rect 137973 15675 138437 15971
rect 138733 15675 139197 15971
rect 139493 15675 139957 15971
rect 140253 15675 140717 15971
rect 141013 15675 141477 15971
rect 141773 15675 142237 15971
rect 142533 15675 142997 15971
rect 143293 15675 143757 15971
rect 144053 15675 144517 15971
rect 144813 15675 145277 15971
rect 145573 15675 146037 15971
rect 146333 15675 146797 15971
rect 147093 15675 147557 15971
rect 147853 15675 148317 15971
rect 148613 15675 149077 15971
rect 149373 15675 149837 15971
rect 150133 15675 150597 15971
rect 150893 15675 151357 15971
rect 151653 15675 152117 15971
rect 152413 15675 152877 15971
rect 153173 15675 153637 15971
rect 153933 15675 154397 15971
rect 154693 15675 155425 15971
rect 135425 15211 155425 15675
rect 135425 14915 136157 15211
rect 136453 14915 136917 15211
rect 137213 14915 137677 15211
rect 137973 14915 138437 15211
rect 138733 14915 139197 15211
rect 139493 14915 139957 15211
rect 140253 14915 140717 15211
rect 141013 14915 141477 15211
rect 141773 14915 142237 15211
rect 142533 14915 142997 15211
rect 143293 14915 143757 15211
rect 144053 14915 144517 15211
rect 144813 14915 145277 15211
rect 145573 14915 146037 15211
rect 146333 14915 146797 15211
rect 147093 14915 147557 15211
rect 147853 14915 148317 15211
rect 148613 14915 149077 15211
rect 149373 14915 149837 15211
rect 150133 14915 150597 15211
rect 150893 14915 151357 15211
rect 151653 14915 152117 15211
rect 152413 14915 152877 15211
rect 153173 14915 153637 15211
rect 153933 14915 154397 15211
rect 154693 14915 155425 15211
rect 135425 14451 155425 14915
rect 135425 14155 136157 14451
rect 136453 14155 136917 14451
rect 137213 14155 137677 14451
rect 137973 14155 138437 14451
rect 138733 14155 139197 14451
rect 139493 14155 139957 14451
rect 140253 14155 140717 14451
rect 141013 14155 141477 14451
rect 141773 14155 142237 14451
rect 142533 14155 142997 14451
rect 143293 14155 143757 14451
rect 144053 14155 144517 14451
rect 144813 14155 145277 14451
rect 145573 14155 146037 14451
rect 146333 14155 146797 14451
rect 147093 14155 147557 14451
rect 147853 14155 148317 14451
rect 148613 14155 149077 14451
rect 149373 14155 149837 14451
rect 150133 14155 150597 14451
rect 150893 14155 151357 14451
rect 151653 14155 152117 14451
rect 152413 14155 152877 14451
rect 153173 14155 153637 14451
rect 153933 14155 154397 14451
rect 154693 14155 155425 14451
rect 135425 13691 155425 14155
rect 135425 13395 136157 13691
rect 136453 13395 136917 13691
rect 137213 13395 137677 13691
rect 137973 13395 138437 13691
rect 138733 13395 139197 13691
rect 139493 13395 139957 13691
rect 140253 13395 140717 13691
rect 141013 13395 141477 13691
rect 141773 13395 142237 13691
rect 142533 13395 142997 13691
rect 143293 13395 143757 13691
rect 144053 13395 144517 13691
rect 144813 13395 145277 13691
rect 145573 13395 146037 13691
rect 146333 13395 146797 13691
rect 147093 13395 147557 13691
rect 147853 13395 148317 13691
rect 148613 13395 149077 13691
rect 149373 13395 149837 13691
rect 150133 13395 150597 13691
rect 150893 13395 151357 13691
rect 151653 13395 152117 13691
rect 152413 13395 152877 13691
rect 153173 13395 153637 13691
rect 153933 13395 154397 13691
rect 154693 13395 155425 13691
rect 135425 12931 155425 13395
rect 135425 12635 136157 12931
rect 136453 12635 136917 12931
rect 137213 12635 137677 12931
rect 137973 12635 138437 12931
rect 138733 12635 139197 12931
rect 139493 12635 139957 12931
rect 140253 12635 140717 12931
rect 141013 12635 141477 12931
rect 141773 12635 142237 12931
rect 142533 12635 142997 12931
rect 143293 12635 143757 12931
rect 144053 12635 144517 12931
rect 144813 12635 145277 12931
rect 145573 12635 146037 12931
rect 146333 12635 146797 12931
rect 147093 12635 147557 12931
rect 147853 12635 148317 12931
rect 148613 12635 149077 12931
rect 149373 12635 149837 12931
rect 150133 12635 150597 12931
rect 150893 12635 151357 12931
rect 151653 12635 152117 12931
rect 152413 12635 152877 12931
rect 153173 12635 153637 12931
rect 153933 12635 154397 12931
rect 154693 12635 155425 12931
rect 135425 12171 155425 12635
rect 135425 11875 136157 12171
rect 136453 11875 136917 12171
rect 137213 11875 137677 12171
rect 137973 11875 138437 12171
rect 138733 11875 139197 12171
rect 139493 11875 139957 12171
rect 140253 11875 140717 12171
rect 141013 11875 141477 12171
rect 141773 11875 142237 12171
rect 142533 11875 142997 12171
rect 143293 11875 143757 12171
rect 144053 11875 144517 12171
rect 144813 11875 145277 12171
rect 145573 11875 146037 12171
rect 146333 11875 146797 12171
rect 147093 11875 147557 12171
rect 147853 11875 148317 12171
rect 148613 11875 149077 12171
rect 149373 11875 149837 12171
rect 150133 11875 150597 12171
rect 150893 11875 151357 12171
rect 151653 11875 152117 12171
rect 152413 11875 152877 12171
rect 153173 11875 153637 12171
rect 153933 11875 154397 12171
rect 154693 11875 155425 12171
rect 135425 11411 155425 11875
rect 135425 11115 136157 11411
rect 136453 11115 136917 11411
rect 137213 11115 137677 11411
rect 137973 11115 138437 11411
rect 138733 11115 139197 11411
rect 139493 11115 139957 11411
rect 140253 11115 140717 11411
rect 141013 11115 141477 11411
rect 141773 11115 142237 11411
rect 142533 11115 142997 11411
rect 143293 11115 143757 11411
rect 144053 11115 144517 11411
rect 144813 11115 145277 11411
rect 145573 11115 146037 11411
rect 146333 11115 146797 11411
rect 147093 11115 147557 11411
rect 147853 11115 148317 11411
rect 148613 11115 149077 11411
rect 149373 11115 149837 11411
rect 150133 11115 150597 11411
rect 150893 11115 151357 11411
rect 151653 11115 152117 11411
rect 152413 11115 152877 11411
rect 153173 11115 153637 11411
rect 153933 11115 154397 11411
rect 154693 11115 155425 11411
rect 135425 10651 155425 11115
rect 135425 10355 136157 10651
rect 136453 10355 136917 10651
rect 137213 10355 137677 10651
rect 137973 10355 138437 10651
rect 138733 10355 139197 10651
rect 139493 10355 139957 10651
rect 140253 10355 140717 10651
rect 141013 10355 141477 10651
rect 141773 10355 142237 10651
rect 142533 10355 142997 10651
rect 143293 10355 143757 10651
rect 144053 10355 144517 10651
rect 144813 10355 145277 10651
rect 145573 10355 146037 10651
rect 146333 10355 146797 10651
rect 147093 10355 147557 10651
rect 147853 10355 148317 10651
rect 148613 10355 149077 10651
rect 149373 10355 149837 10651
rect 150133 10355 150597 10651
rect 150893 10355 151357 10651
rect 151653 10355 152117 10651
rect 152413 10355 152877 10651
rect 153173 10355 153637 10651
rect 153933 10355 154397 10651
rect 154693 10355 155425 10651
rect 135425 9891 155425 10355
rect 135425 9595 136157 9891
rect 136453 9595 136917 9891
rect 137213 9595 137677 9891
rect 137973 9595 138437 9891
rect 138733 9595 139197 9891
rect 139493 9595 139957 9891
rect 140253 9595 140717 9891
rect 141013 9595 141477 9891
rect 141773 9595 142237 9891
rect 142533 9595 142997 9891
rect 143293 9595 143757 9891
rect 144053 9595 144517 9891
rect 144813 9595 145277 9891
rect 145573 9595 146037 9891
rect 146333 9595 146797 9891
rect 147093 9595 147557 9891
rect 147853 9595 148317 9891
rect 148613 9595 149077 9891
rect 149373 9595 149837 9891
rect 150133 9595 150597 9891
rect 150893 9595 151357 9891
rect 151653 9595 152117 9891
rect 152413 9595 152877 9891
rect 153173 9595 153637 9891
rect 153933 9595 154397 9891
rect 154693 9595 155425 9891
rect 135425 9131 155425 9595
rect 135425 8835 136157 9131
rect 136453 8835 136917 9131
rect 137213 8835 137677 9131
rect 137973 8835 138437 9131
rect 138733 8835 139197 9131
rect 139493 8835 139957 9131
rect 140253 8835 140717 9131
rect 141013 8835 141477 9131
rect 141773 8835 142237 9131
rect 142533 8835 142997 9131
rect 143293 8835 143757 9131
rect 144053 8835 144517 9131
rect 144813 8835 145277 9131
rect 145573 8835 146037 9131
rect 146333 8835 146797 9131
rect 147093 8835 147557 9131
rect 147853 8835 148317 9131
rect 148613 8835 149077 9131
rect 149373 8835 149837 9131
rect 150133 8835 150597 9131
rect 150893 8835 151357 9131
rect 151653 8835 152117 9131
rect 152413 8835 152877 9131
rect 153173 8835 153637 9131
rect 153933 8835 154397 9131
rect 154693 8835 155425 9131
rect 135425 8371 155425 8835
rect 135425 8075 136157 8371
rect 136453 8075 136917 8371
rect 137213 8075 137677 8371
rect 137973 8075 138437 8371
rect 138733 8075 139197 8371
rect 139493 8075 139957 8371
rect 140253 8075 140717 8371
rect 141013 8075 141477 8371
rect 141773 8075 142237 8371
rect 142533 8075 142997 8371
rect 143293 8075 143757 8371
rect 144053 8075 144517 8371
rect 144813 8075 145277 8371
rect 145573 8075 146037 8371
rect 146333 8075 146797 8371
rect 147093 8075 147557 8371
rect 147853 8075 148317 8371
rect 148613 8075 149077 8371
rect 149373 8075 149837 8371
rect 150133 8075 150597 8371
rect 150893 8075 151357 8371
rect 151653 8075 152117 8371
rect 152413 8075 152877 8371
rect 153173 8075 153637 8371
rect 153933 8075 154397 8371
rect 154693 8075 155425 8371
rect 135425 7611 155425 8075
rect 135425 7315 136157 7611
rect 136453 7315 136917 7611
rect 137213 7315 137677 7611
rect 137973 7315 138437 7611
rect 138733 7315 139197 7611
rect 139493 7315 139957 7611
rect 140253 7315 140717 7611
rect 141013 7315 141477 7611
rect 141773 7315 142237 7611
rect 142533 7315 142997 7611
rect 143293 7315 143757 7611
rect 144053 7315 144517 7611
rect 144813 7315 145277 7611
rect 145573 7315 146037 7611
rect 146333 7315 146797 7611
rect 147093 7315 147557 7611
rect 147853 7315 148317 7611
rect 148613 7315 149077 7611
rect 149373 7315 149837 7611
rect 150133 7315 150597 7611
rect 150893 7315 151357 7611
rect 151653 7315 152117 7611
rect 152413 7315 152877 7611
rect 153173 7315 153637 7611
rect 153933 7315 154397 7611
rect 154693 7315 155425 7611
rect 135425 6743 155425 7315
rect 157225 31171 177225 31743
rect 157225 30875 157957 31171
rect 158253 30875 158717 31171
rect 159013 30875 159477 31171
rect 159773 30875 160237 31171
rect 160533 30875 160997 31171
rect 161293 30875 161757 31171
rect 162053 30875 162517 31171
rect 162813 30875 163277 31171
rect 163573 30875 164037 31171
rect 164333 30875 164797 31171
rect 165093 30875 165557 31171
rect 165853 30875 166317 31171
rect 166613 30875 167077 31171
rect 167373 30875 167837 31171
rect 168133 30875 168597 31171
rect 168893 30875 169357 31171
rect 169653 30875 170117 31171
rect 170413 30875 170877 31171
rect 171173 30875 171637 31171
rect 171933 30875 172397 31171
rect 172693 30875 173157 31171
rect 173453 30875 173917 31171
rect 174213 30875 174677 31171
rect 174973 30875 175437 31171
rect 175733 30875 176197 31171
rect 176493 30875 177225 31171
rect 157225 30411 177225 30875
rect 157225 30115 157957 30411
rect 158253 30115 158717 30411
rect 159013 30115 159477 30411
rect 159773 30115 160237 30411
rect 160533 30115 160997 30411
rect 161293 30115 161757 30411
rect 162053 30115 162517 30411
rect 162813 30115 163277 30411
rect 163573 30115 164037 30411
rect 164333 30115 164797 30411
rect 165093 30115 165557 30411
rect 165853 30115 166317 30411
rect 166613 30115 167077 30411
rect 167373 30115 167837 30411
rect 168133 30115 168597 30411
rect 168893 30115 169357 30411
rect 169653 30115 170117 30411
rect 170413 30115 170877 30411
rect 171173 30115 171637 30411
rect 171933 30115 172397 30411
rect 172693 30115 173157 30411
rect 173453 30115 173917 30411
rect 174213 30115 174677 30411
rect 174973 30115 175437 30411
rect 175733 30115 176197 30411
rect 176493 30115 177225 30411
rect 157225 29651 177225 30115
rect 157225 29355 157957 29651
rect 158253 29355 158717 29651
rect 159013 29355 159477 29651
rect 159773 29355 160237 29651
rect 160533 29355 160997 29651
rect 161293 29355 161757 29651
rect 162053 29355 162517 29651
rect 162813 29355 163277 29651
rect 163573 29355 164037 29651
rect 164333 29355 164797 29651
rect 165093 29355 165557 29651
rect 165853 29355 166317 29651
rect 166613 29355 167077 29651
rect 167373 29355 167837 29651
rect 168133 29355 168597 29651
rect 168893 29355 169357 29651
rect 169653 29355 170117 29651
rect 170413 29355 170877 29651
rect 171173 29355 171637 29651
rect 171933 29355 172397 29651
rect 172693 29355 173157 29651
rect 173453 29355 173917 29651
rect 174213 29355 174677 29651
rect 174973 29355 175437 29651
rect 175733 29355 176197 29651
rect 176493 29355 177225 29651
rect 157225 28891 177225 29355
rect 157225 28595 157957 28891
rect 158253 28595 158717 28891
rect 159013 28595 159477 28891
rect 159773 28595 160237 28891
rect 160533 28595 160997 28891
rect 161293 28595 161757 28891
rect 162053 28595 162517 28891
rect 162813 28595 163277 28891
rect 163573 28595 164037 28891
rect 164333 28595 164797 28891
rect 165093 28595 165557 28891
rect 165853 28595 166317 28891
rect 166613 28595 167077 28891
rect 167373 28595 167837 28891
rect 168133 28595 168597 28891
rect 168893 28595 169357 28891
rect 169653 28595 170117 28891
rect 170413 28595 170877 28891
rect 171173 28595 171637 28891
rect 171933 28595 172397 28891
rect 172693 28595 173157 28891
rect 173453 28595 173917 28891
rect 174213 28595 174677 28891
rect 174973 28595 175437 28891
rect 175733 28595 176197 28891
rect 176493 28595 177225 28891
rect 157225 28131 177225 28595
rect 157225 27835 157957 28131
rect 158253 27835 158717 28131
rect 159013 27835 159477 28131
rect 159773 27835 160237 28131
rect 160533 27835 160997 28131
rect 161293 27835 161757 28131
rect 162053 27835 162517 28131
rect 162813 27835 163277 28131
rect 163573 27835 164037 28131
rect 164333 27835 164797 28131
rect 165093 27835 165557 28131
rect 165853 27835 166317 28131
rect 166613 27835 167077 28131
rect 167373 27835 167837 28131
rect 168133 27835 168597 28131
rect 168893 27835 169357 28131
rect 169653 27835 170117 28131
rect 170413 27835 170877 28131
rect 171173 27835 171637 28131
rect 171933 27835 172397 28131
rect 172693 27835 173157 28131
rect 173453 27835 173917 28131
rect 174213 27835 174677 28131
rect 174973 27835 175437 28131
rect 175733 27835 176197 28131
rect 176493 27835 177225 28131
rect 157225 27371 177225 27835
rect 157225 27075 157957 27371
rect 158253 27075 158717 27371
rect 159013 27075 159477 27371
rect 159773 27075 160237 27371
rect 160533 27075 160997 27371
rect 161293 27075 161757 27371
rect 162053 27075 162517 27371
rect 162813 27075 163277 27371
rect 163573 27075 164037 27371
rect 164333 27075 164797 27371
rect 165093 27075 165557 27371
rect 165853 27075 166317 27371
rect 166613 27075 167077 27371
rect 167373 27075 167837 27371
rect 168133 27075 168597 27371
rect 168893 27075 169357 27371
rect 169653 27075 170117 27371
rect 170413 27075 170877 27371
rect 171173 27075 171637 27371
rect 171933 27075 172397 27371
rect 172693 27075 173157 27371
rect 173453 27075 173917 27371
rect 174213 27075 174677 27371
rect 174973 27075 175437 27371
rect 175733 27075 176197 27371
rect 176493 27075 177225 27371
rect 157225 26611 177225 27075
rect 157225 26315 157957 26611
rect 158253 26315 158717 26611
rect 159013 26315 159477 26611
rect 159773 26315 160237 26611
rect 160533 26315 160997 26611
rect 161293 26315 161757 26611
rect 162053 26315 162517 26611
rect 162813 26315 163277 26611
rect 163573 26315 164037 26611
rect 164333 26315 164797 26611
rect 165093 26315 165557 26611
rect 165853 26315 166317 26611
rect 166613 26315 167077 26611
rect 167373 26315 167837 26611
rect 168133 26315 168597 26611
rect 168893 26315 169357 26611
rect 169653 26315 170117 26611
rect 170413 26315 170877 26611
rect 171173 26315 171637 26611
rect 171933 26315 172397 26611
rect 172693 26315 173157 26611
rect 173453 26315 173917 26611
rect 174213 26315 174677 26611
rect 174973 26315 175437 26611
rect 175733 26315 176197 26611
rect 176493 26315 177225 26611
rect 157225 25851 177225 26315
rect 157225 25555 157957 25851
rect 158253 25555 158717 25851
rect 159013 25555 159477 25851
rect 159773 25555 160237 25851
rect 160533 25555 160997 25851
rect 161293 25555 161757 25851
rect 162053 25555 162517 25851
rect 162813 25555 163277 25851
rect 163573 25555 164037 25851
rect 164333 25555 164797 25851
rect 165093 25555 165557 25851
rect 165853 25555 166317 25851
rect 166613 25555 167077 25851
rect 167373 25555 167837 25851
rect 168133 25555 168597 25851
rect 168893 25555 169357 25851
rect 169653 25555 170117 25851
rect 170413 25555 170877 25851
rect 171173 25555 171637 25851
rect 171933 25555 172397 25851
rect 172693 25555 173157 25851
rect 173453 25555 173917 25851
rect 174213 25555 174677 25851
rect 174973 25555 175437 25851
rect 175733 25555 176197 25851
rect 176493 25555 177225 25851
rect 157225 25091 177225 25555
rect 157225 24795 157957 25091
rect 158253 24795 158717 25091
rect 159013 24795 159477 25091
rect 159773 24795 160237 25091
rect 160533 24795 160997 25091
rect 161293 24795 161757 25091
rect 162053 24795 162517 25091
rect 162813 24795 163277 25091
rect 163573 24795 164037 25091
rect 164333 24795 164797 25091
rect 165093 24795 165557 25091
rect 165853 24795 166317 25091
rect 166613 24795 167077 25091
rect 167373 24795 167837 25091
rect 168133 24795 168597 25091
rect 168893 24795 169357 25091
rect 169653 24795 170117 25091
rect 170413 24795 170877 25091
rect 171173 24795 171637 25091
rect 171933 24795 172397 25091
rect 172693 24795 173157 25091
rect 173453 24795 173917 25091
rect 174213 24795 174677 25091
rect 174973 24795 175437 25091
rect 175733 24795 176197 25091
rect 176493 24795 177225 25091
rect 157225 24331 177225 24795
rect 157225 24035 157957 24331
rect 158253 24035 158717 24331
rect 159013 24035 159477 24331
rect 159773 24035 160237 24331
rect 160533 24035 160997 24331
rect 161293 24035 161757 24331
rect 162053 24035 162517 24331
rect 162813 24035 163277 24331
rect 163573 24035 164037 24331
rect 164333 24035 164797 24331
rect 165093 24035 165557 24331
rect 165853 24035 166317 24331
rect 166613 24035 167077 24331
rect 167373 24035 167837 24331
rect 168133 24035 168597 24331
rect 168893 24035 169357 24331
rect 169653 24035 170117 24331
rect 170413 24035 170877 24331
rect 171173 24035 171637 24331
rect 171933 24035 172397 24331
rect 172693 24035 173157 24331
rect 173453 24035 173917 24331
rect 174213 24035 174677 24331
rect 174973 24035 175437 24331
rect 175733 24035 176197 24331
rect 176493 24035 177225 24331
rect 157225 23571 177225 24035
rect 157225 23275 157957 23571
rect 158253 23275 158717 23571
rect 159013 23275 159477 23571
rect 159773 23275 160237 23571
rect 160533 23275 160997 23571
rect 161293 23275 161757 23571
rect 162053 23275 162517 23571
rect 162813 23275 163277 23571
rect 163573 23275 164037 23571
rect 164333 23275 164797 23571
rect 165093 23275 165557 23571
rect 165853 23275 166317 23571
rect 166613 23275 167077 23571
rect 167373 23275 167837 23571
rect 168133 23275 168597 23571
rect 168893 23275 169357 23571
rect 169653 23275 170117 23571
rect 170413 23275 170877 23571
rect 171173 23275 171637 23571
rect 171933 23275 172397 23571
rect 172693 23275 173157 23571
rect 173453 23275 173917 23571
rect 174213 23275 174677 23571
rect 174973 23275 175437 23571
rect 175733 23275 176197 23571
rect 176493 23275 177225 23571
rect 157225 22811 177225 23275
rect 157225 22515 157957 22811
rect 158253 22515 158717 22811
rect 159013 22515 159477 22811
rect 159773 22515 160237 22811
rect 160533 22515 160997 22811
rect 161293 22515 161757 22811
rect 162053 22515 162517 22811
rect 162813 22515 163277 22811
rect 163573 22515 164037 22811
rect 164333 22515 164797 22811
rect 165093 22515 165557 22811
rect 165853 22515 166317 22811
rect 166613 22515 167077 22811
rect 167373 22515 167837 22811
rect 168133 22515 168597 22811
rect 168893 22515 169357 22811
rect 169653 22515 170117 22811
rect 170413 22515 170877 22811
rect 171173 22515 171637 22811
rect 171933 22515 172397 22811
rect 172693 22515 173157 22811
rect 173453 22515 173917 22811
rect 174213 22515 174677 22811
rect 174973 22515 175437 22811
rect 175733 22515 176197 22811
rect 176493 22515 177225 22811
rect 157225 22051 177225 22515
rect 157225 21755 157957 22051
rect 158253 21755 158717 22051
rect 159013 21755 159477 22051
rect 159773 21755 160237 22051
rect 160533 21755 160997 22051
rect 161293 21755 161757 22051
rect 162053 21755 162517 22051
rect 162813 21755 163277 22051
rect 163573 21755 164037 22051
rect 164333 21755 164797 22051
rect 165093 21755 165557 22051
rect 165853 21755 166317 22051
rect 166613 21755 167077 22051
rect 167373 21755 167837 22051
rect 168133 21755 168597 22051
rect 168893 21755 169357 22051
rect 169653 21755 170117 22051
rect 170413 21755 170877 22051
rect 171173 21755 171637 22051
rect 171933 21755 172397 22051
rect 172693 21755 173157 22051
rect 173453 21755 173917 22051
rect 174213 21755 174677 22051
rect 174973 21755 175437 22051
rect 175733 21755 176197 22051
rect 176493 21755 177225 22051
rect 157225 21291 177225 21755
rect 157225 20995 157957 21291
rect 158253 20995 158717 21291
rect 159013 20995 159477 21291
rect 159773 20995 160237 21291
rect 160533 20995 160997 21291
rect 161293 20995 161757 21291
rect 162053 20995 162517 21291
rect 162813 20995 163277 21291
rect 163573 20995 164037 21291
rect 164333 20995 164797 21291
rect 165093 20995 165557 21291
rect 165853 20995 166317 21291
rect 166613 20995 167077 21291
rect 167373 20995 167837 21291
rect 168133 20995 168597 21291
rect 168893 20995 169357 21291
rect 169653 20995 170117 21291
rect 170413 20995 170877 21291
rect 171173 20995 171637 21291
rect 171933 20995 172397 21291
rect 172693 20995 173157 21291
rect 173453 20995 173917 21291
rect 174213 20995 174677 21291
rect 174973 20995 175437 21291
rect 175733 20995 176197 21291
rect 176493 20995 177225 21291
rect 157225 20531 177225 20995
rect 157225 20235 157957 20531
rect 158253 20235 158717 20531
rect 159013 20235 159477 20531
rect 159773 20235 160237 20531
rect 160533 20235 160997 20531
rect 161293 20235 161757 20531
rect 162053 20235 162517 20531
rect 162813 20235 163277 20531
rect 163573 20235 164037 20531
rect 164333 20235 164797 20531
rect 165093 20235 165557 20531
rect 165853 20235 166317 20531
rect 166613 20235 167077 20531
rect 167373 20235 167837 20531
rect 168133 20235 168597 20531
rect 168893 20235 169357 20531
rect 169653 20235 170117 20531
rect 170413 20235 170877 20531
rect 171173 20235 171637 20531
rect 171933 20235 172397 20531
rect 172693 20235 173157 20531
rect 173453 20235 173917 20531
rect 174213 20235 174677 20531
rect 174973 20235 175437 20531
rect 175733 20235 176197 20531
rect 176493 20235 177225 20531
rect 157225 19771 177225 20235
rect 157225 19475 157957 19771
rect 158253 19475 158717 19771
rect 159013 19475 159477 19771
rect 159773 19475 160237 19771
rect 160533 19475 160997 19771
rect 161293 19475 161757 19771
rect 162053 19475 162517 19771
rect 162813 19475 163277 19771
rect 163573 19475 164037 19771
rect 164333 19475 164797 19771
rect 165093 19475 165557 19771
rect 165853 19475 166317 19771
rect 166613 19475 167077 19771
rect 167373 19475 167837 19771
rect 168133 19475 168597 19771
rect 168893 19475 169357 19771
rect 169653 19475 170117 19771
rect 170413 19475 170877 19771
rect 171173 19475 171637 19771
rect 171933 19475 172397 19771
rect 172693 19475 173157 19771
rect 173453 19475 173917 19771
rect 174213 19475 174677 19771
rect 174973 19475 175437 19771
rect 175733 19475 176197 19771
rect 176493 19475 177225 19771
rect 157225 19011 177225 19475
rect 157225 18715 157957 19011
rect 158253 18715 158717 19011
rect 159013 18715 159477 19011
rect 159773 18715 160237 19011
rect 160533 18715 160997 19011
rect 161293 18715 161757 19011
rect 162053 18715 162517 19011
rect 162813 18715 163277 19011
rect 163573 18715 164037 19011
rect 164333 18715 164797 19011
rect 165093 18715 165557 19011
rect 165853 18715 166317 19011
rect 166613 18715 167077 19011
rect 167373 18715 167837 19011
rect 168133 18715 168597 19011
rect 168893 18715 169357 19011
rect 169653 18715 170117 19011
rect 170413 18715 170877 19011
rect 171173 18715 171637 19011
rect 171933 18715 172397 19011
rect 172693 18715 173157 19011
rect 173453 18715 173917 19011
rect 174213 18715 174677 19011
rect 174973 18715 175437 19011
rect 175733 18715 176197 19011
rect 176493 18715 177225 19011
rect 157225 18251 177225 18715
rect 157225 17955 157957 18251
rect 158253 17955 158717 18251
rect 159013 17955 159477 18251
rect 159773 17955 160237 18251
rect 160533 17955 160997 18251
rect 161293 17955 161757 18251
rect 162053 17955 162517 18251
rect 162813 17955 163277 18251
rect 163573 17955 164037 18251
rect 164333 17955 164797 18251
rect 165093 17955 165557 18251
rect 165853 17955 166317 18251
rect 166613 17955 167077 18251
rect 167373 17955 167837 18251
rect 168133 17955 168597 18251
rect 168893 17955 169357 18251
rect 169653 17955 170117 18251
rect 170413 17955 170877 18251
rect 171173 17955 171637 18251
rect 171933 17955 172397 18251
rect 172693 17955 173157 18251
rect 173453 17955 173917 18251
rect 174213 17955 174677 18251
rect 174973 17955 175437 18251
rect 175733 17955 176197 18251
rect 176493 17955 177225 18251
rect 157225 17491 177225 17955
rect 157225 17195 157957 17491
rect 158253 17195 158717 17491
rect 159013 17195 159477 17491
rect 159773 17195 160237 17491
rect 160533 17195 160997 17491
rect 161293 17195 161757 17491
rect 162053 17195 162517 17491
rect 162813 17195 163277 17491
rect 163573 17195 164037 17491
rect 164333 17195 164797 17491
rect 165093 17195 165557 17491
rect 165853 17195 166317 17491
rect 166613 17195 167077 17491
rect 167373 17195 167837 17491
rect 168133 17195 168597 17491
rect 168893 17195 169357 17491
rect 169653 17195 170117 17491
rect 170413 17195 170877 17491
rect 171173 17195 171637 17491
rect 171933 17195 172397 17491
rect 172693 17195 173157 17491
rect 173453 17195 173917 17491
rect 174213 17195 174677 17491
rect 174973 17195 175437 17491
rect 175733 17195 176197 17491
rect 176493 17195 177225 17491
rect 157225 16731 177225 17195
rect 157225 16435 157957 16731
rect 158253 16435 158717 16731
rect 159013 16435 159477 16731
rect 159773 16435 160237 16731
rect 160533 16435 160997 16731
rect 161293 16435 161757 16731
rect 162053 16435 162517 16731
rect 162813 16435 163277 16731
rect 163573 16435 164037 16731
rect 164333 16435 164797 16731
rect 165093 16435 165557 16731
rect 165853 16435 166317 16731
rect 166613 16435 167077 16731
rect 167373 16435 167837 16731
rect 168133 16435 168597 16731
rect 168893 16435 169357 16731
rect 169653 16435 170117 16731
rect 170413 16435 170877 16731
rect 171173 16435 171637 16731
rect 171933 16435 172397 16731
rect 172693 16435 173157 16731
rect 173453 16435 173917 16731
rect 174213 16435 174677 16731
rect 174973 16435 175437 16731
rect 175733 16435 176197 16731
rect 176493 16435 177225 16731
rect 157225 15971 177225 16435
rect 157225 15675 157957 15971
rect 158253 15675 158717 15971
rect 159013 15675 159477 15971
rect 159773 15675 160237 15971
rect 160533 15675 160997 15971
rect 161293 15675 161757 15971
rect 162053 15675 162517 15971
rect 162813 15675 163277 15971
rect 163573 15675 164037 15971
rect 164333 15675 164797 15971
rect 165093 15675 165557 15971
rect 165853 15675 166317 15971
rect 166613 15675 167077 15971
rect 167373 15675 167837 15971
rect 168133 15675 168597 15971
rect 168893 15675 169357 15971
rect 169653 15675 170117 15971
rect 170413 15675 170877 15971
rect 171173 15675 171637 15971
rect 171933 15675 172397 15971
rect 172693 15675 173157 15971
rect 173453 15675 173917 15971
rect 174213 15675 174677 15971
rect 174973 15675 175437 15971
rect 175733 15675 176197 15971
rect 176493 15675 177225 15971
rect 157225 15211 177225 15675
rect 157225 14915 157957 15211
rect 158253 14915 158717 15211
rect 159013 14915 159477 15211
rect 159773 14915 160237 15211
rect 160533 14915 160997 15211
rect 161293 14915 161757 15211
rect 162053 14915 162517 15211
rect 162813 14915 163277 15211
rect 163573 14915 164037 15211
rect 164333 14915 164797 15211
rect 165093 14915 165557 15211
rect 165853 14915 166317 15211
rect 166613 14915 167077 15211
rect 167373 14915 167837 15211
rect 168133 14915 168597 15211
rect 168893 14915 169357 15211
rect 169653 14915 170117 15211
rect 170413 14915 170877 15211
rect 171173 14915 171637 15211
rect 171933 14915 172397 15211
rect 172693 14915 173157 15211
rect 173453 14915 173917 15211
rect 174213 14915 174677 15211
rect 174973 14915 175437 15211
rect 175733 14915 176197 15211
rect 176493 14915 177225 15211
rect 157225 14451 177225 14915
rect 157225 14155 157957 14451
rect 158253 14155 158717 14451
rect 159013 14155 159477 14451
rect 159773 14155 160237 14451
rect 160533 14155 160997 14451
rect 161293 14155 161757 14451
rect 162053 14155 162517 14451
rect 162813 14155 163277 14451
rect 163573 14155 164037 14451
rect 164333 14155 164797 14451
rect 165093 14155 165557 14451
rect 165853 14155 166317 14451
rect 166613 14155 167077 14451
rect 167373 14155 167837 14451
rect 168133 14155 168597 14451
rect 168893 14155 169357 14451
rect 169653 14155 170117 14451
rect 170413 14155 170877 14451
rect 171173 14155 171637 14451
rect 171933 14155 172397 14451
rect 172693 14155 173157 14451
rect 173453 14155 173917 14451
rect 174213 14155 174677 14451
rect 174973 14155 175437 14451
rect 175733 14155 176197 14451
rect 176493 14155 177225 14451
rect 157225 13691 177225 14155
rect 157225 13395 157957 13691
rect 158253 13395 158717 13691
rect 159013 13395 159477 13691
rect 159773 13395 160237 13691
rect 160533 13395 160997 13691
rect 161293 13395 161757 13691
rect 162053 13395 162517 13691
rect 162813 13395 163277 13691
rect 163573 13395 164037 13691
rect 164333 13395 164797 13691
rect 165093 13395 165557 13691
rect 165853 13395 166317 13691
rect 166613 13395 167077 13691
rect 167373 13395 167837 13691
rect 168133 13395 168597 13691
rect 168893 13395 169357 13691
rect 169653 13395 170117 13691
rect 170413 13395 170877 13691
rect 171173 13395 171637 13691
rect 171933 13395 172397 13691
rect 172693 13395 173157 13691
rect 173453 13395 173917 13691
rect 174213 13395 174677 13691
rect 174973 13395 175437 13691
rect 175733 13395 176197 13691
rect 176493 13395 177225 13691
rect 157225 12931 177225 13395
rect 157225 12635 157957 12931
rect 158253 12635 158717 12931
rect 159013 12635 159477 12931
rect 159773 12635 160237 12931
rect 160533 12635 160997 12931
rect 161293 12635 161757 12931
rect 162053 12635 162517 12931
rect 162813 12635 163277 12931
rect 163573 12635 164037 12931
rect 164333 12635 164797 12931
rect 165093 12635 165557 12931
rect 165853 12635 166317 12931
rect 166613 12635 167077 12931
rect 167373 12635 167837 12931
rect 168133 12635 168597 12931
rect 168893 12635 169357 12931
rect 169653 12635 170117 12931
rect 170413 12635 170877 12931
rect 171173 12635 171637 12931
rect 171933 12635 172397 12931
rect 172693 12635 173157 12931
rect 173453 12635 173917 12931
rect 174213 12635 174677 12931
rect 174973 12635 175437 12931
rect 175733 12635 176197 12931
rect 176493 12635 177225 12931
rect 157225 12171 177225 12635
rect 157225 11875 157957 12171
rect 158253 11875 158717 12171
rect 159013 11875 159477 12171
rect 159773 11875 160237 12171
rect 160533 11875 160997 12171
rect 161293 11875 161757 12171
rect 162053 11875 162517 12171
rect 162813 11875 163277 12171
rect 163573 11875 164037 12171
rect 164333 11875 164797 12171
rect 165093 11875 165557 12171
rect 165853 11875 166317 12171
rect 166613 11875 167077 12171
rect 167373 11875 167837 12171
rect 168133 11875 168597 12171
rect 168893 11875 169357 12171
rect 169653 11875 170117 12171
rect 170413 11875 170877 12171
rect 171173 11875 171637 12171
rect 171933 11875 172397 12171
rect 172693 11875 173157 12171
rect 173453 11875 173917 12171
rect 174213 11875 174677 12171
rect 174973 11875 175437 12171
rect 175733 11875 176197 12171
rect 176493 11875 177225 12171
rect 157225 11411 177225 11875
rect 157225 11115 157957 11411
rect 158253 11115 158717 11411
rect 159013 11115 159477 11411
rect 159773 11115 160237 11411
rect 160533 11115 160997 11411
rect 161293 11115 161757 11411
rect 162053 11115 162517 11411
rect 162813 11115 163277 11411
rect 163573 11115 164037 11411
rect 164333 11115 164797 11411
rect 165093 11115 165557 11411
rect 165853 11115 166317 11411
rect 166613 11115 167077 11411
rect 167373 11115 167837 11411
rect 168133 11115 168597 11411
rect 168893 11115 169357 11411
rect 169653 11115 170117 11411
rect 170413 11115 170877 11411
rect 171173 11115 171637 11411
rect 171933 11115 172397 11411
rect 172693 11115 173157 11411
rect 173453 11115 173917 11411
rect 174213 11115 174677 11411
rect 174973 11115 175437 11411
rect 175733 11115 176197 11411
rect 176493 11115 177225 11411
rect 157225 10651 177225 11115
rect 157225 10355 157957 10651
rect 158253 10355 158717 10651
rect 159013 10355 159477 10651
rect 159773 10355 160237 10651
rect 160533 10355 160997 10651
rect 161293 10355 161757 10651
rect 162053 10355 162517 10651
rect 162813 10355 163277 10651
rect 163573 10355 164037 10651
rect 164333 10355 164797 10651
rect 165093 10355 165557 10651
rect 165853 10355 166317 10651
rect 166613 10355 167077 10651
rect 167373 10355 167837 10651
rect 168133 10355 168597 10651
rect 168893 10355 169357 10651
rect 169653 10355 170117 10651
rect 170413 10355 170877 10651
rect 171173 10355 171637 10651
rect 171933 10355 172397 10651
rect 172693 10355 173157 10651
rect 173453 10355 173917 10651
rect 174213 10355 174677 10651
rect 174973 10355 175437 10651
rect 175733 10355 176197 10651
rect 176493 10355 177225 10651
rect 157225 9891 177225 10355
rect 157225 9595 157957 9891
rect 158253 9595 158717 9891
rect 159013 9595 159477 9891
rect 159773 9595 160237 9891
rect 160533 9595 160997 9891
rect 161293 9595 161757 9891
rect 162053 9595 162517 9891
rect 162813 9595 163277 9891
rect 163573 9595 164037 9891
rect 164333 9595 164797 9891
rect 165093 9595 165557 9891
rect 165853 9595 166317 9891
rect 166613 9595 167077 9891
rect 167373 9595 167837 9891
rect 168133 9595 168597 9891
rect 168893 9595 169357 9891
rect 169653 9595 170117 9891
rect 170413 9595 170877 9891
rect 171173 9595 171637 9891
rect 171933 9595 172397 9891
rect 172693 9595 173157 9891
rect 173453 9595 173917 9891
rect 174213 9595 174677 9891
rect 174973 9595 175437 9891
rect 175733 9595 176197 9891
rect 176493 9595 177225 9891
rect 157225 9131 177225 9595
rect 157225 8835 157957 9131
rect 158253 8835 158717 9131
rect 159013 8835 159477 9131
rect 159773 8835 160237 9131
rect 160533 8835 160997 9131
rect 161293 8835 161757 9131
rect 162053 8835 162517 9131
rect 162813 8835 163277 9131
rect 163573 8835 164037 9131
rect 164333 8835 164797 9131
rect 165093 8835 165557 9131
rect 165853 8835 166317 9131
rect 166613 8835 167077 9131
rect 167373 8835 167837 9131
rect 168133 8835 168597 9131
rect 168893 8835 169357 9131
rect 169653 8835 170117 9131
rect 170413 8835 170877 9131
rect 171173 8835 171637 9131
rect 171933 8835 172397 9131
rect 172693 8835 173157 9131
rect 173453 8835 173917 9131
rect 174213 8835 174677 9131
rect 174973 8835 175437 9131
rect 175733 8835 176197 9131
rect 176493 8835 177225 9131
rect 157225 8371 177225 8835
rect 157225 8075 157957 8371
rect 158253 8075 158717 8371
rect 159013 8075 159477 8371
rect 159773 8075 160237 8371
rect 160533 8075 160997 8371
rect 161293 8075 161757 8371
rect 162053 8075 162517 8371
rect 162813 8075 163277 8371
rect 163573 8075 164037 8371
rect 164333 8075 164797 8371
rect 165093 8075 165557 8371
rect 165853 8075 166317 8371
rect 166613 8075 167077 8371
rect 167373 8075 167837 8371
rect 168133 8075 168597 8371
rect 168893 8075 169357 8371
rect 169653 8075 170117 8371
rect 170413 8075 170877 8371
rect 171173 8075 171637 8371
rect 171933 8075 172397 8371
rect 172693 8075 173157 8371
rect 173453 8075 173917 8371
rect 174213 8075 174677 8371
rect 174973 8075 175437 8371
rect 175733 8075 176197 8371
rect 176493 8075 177225 8371
rect 157225 7611 177225 8075
rect 157225 7315 157957 7611
rect 158253 7315 158717 7611
rect 159013 7315 159477 7611
rect 159773 7315 160237 7611
rect 160533 7315 160997 7611
rect 161293 7315 161757 7611
rect 162053 7315 162517 7611
rect 162813 7315 163277 7611
rect 163573 7315 164037 7611
rect 164333 7315 164797 7611
rect 165093 7315 165557 7611
rect 165853 7315 166317 7611
rect 166613 7315 167077 7611
rect 167373 7315 167837 7611
rect 168133 7315 168597 7611
rect 168893 7315 169357 7611
rect 169653 7315 170117 7611
rect 170413 7315 170877 7611
rect 171173 7315 171637 7611
rect 171933 7315 172397 7611
rect 172693 7315 173157 7611
rect 173453 7315 173917 7611
rect 174213 7315 174677 7611
rect 174973 7315 175437 7611
rect 175733 7315 176197 7611
rect 176493 7315 177225 7611
rect 157225 6743 177225 7315
rect 186505 28984 211505 29716
rect 186505 28688 187077 28984
rect 187373 28688 187837 28984
rect 188133 28688 188597 28984
rect 188893 28688 189357 28984
rect 189653 28688 190117 28984
rect 190413 28688 190877 28984
rect 191173 28688 191637 28984
rect 191933 28688 192397 28984
rect 192693 28688 193157 28984
rect 193453 28688 193917 28984
rect 194213 28688 194677 28984
rect 194973 28688 195437 28984
rect 195733 28688 196197 28984
rect 196493 28688 196957 28984
rect 197253 28688 197717 28984
rect 198013 28688 198477 28984
rect 198773 28688 199237 28984
rect 199533 28688 199997 28984
rect 200293 28688 200757 28984
rect 201053 28688 201517 28984
rect 201813 28688 202277 28984
rect 202573 28688 203037 28984
rect 203333 28688 203797 28984
rect 204093 28688 204557 28984
rect 204853 28688 205317 28984
rect 205613 28688 206077 28984
rect 206373 28688 206837 28984
rect 207133 28688 207597 28984
rect 207893 28688 208357 28984
rect 208653 28688 209117 28984
rect 209413 28688 209877 28984
rect 210173 28688 210637 28984
rect 210933 28688 211505 28984
rect 186505 28224 211505 28688
rect 186505 27928 187077 28224
rect 187373 27928 187837 28224
rect 188133 27928 188597 28224
rect 188893 27928 189357 28224
rect 189653 27928 190117 28224
rect 190413 27928 190877 28224
rect 191173 27928 191637 28224
rect 191933 27928 192397 28224
rect 192693 27928 193157 28224
rect 193453 27928 193917 28224
rect 194213 27928 194677 28224
rect 194973 27928 195437 28224
rect 195733 27928 196197 28224
rect 196493 27928 196957 28224
rect 197253 27928 197717 28224
rect 198013 27928 198477 28224
rect 198773 27928 199237 28224
rect 199533 27928 199997 28224
rect 200293 27928 200757 28224
rect 201053 27928 201517 28224
rect 201813 27928 202277 28224
rect 202573 27928 203037 28224
rect 203333 27928 203797 28224
rect 204093 27928 204557 28224
rect 204853 27928 205317 28224
rect 205613 27928 206077 28224
rect 206373 27928 206837 28224
rect 207133 27928 207597 28224
rect 207893 27928 208357 28224
rect 208653 27928 209117 28224
rect 209413 27928 209877 28224
rect 210173 27928 210637 28224
rect 210933 27928 211505 28224
rect 186505 27464 211505 27928
rect 186505 27168 187077 27464
rect 187373 27168 187837 27464
rect 188133 27168 188597 27464
rect 188893 27168 189357 27464
rect 189653 27168 190117 27464
rect 190413 27168 190877 27464
rect 191173 27168 191637 27464
rect 191933 27168 192397 27464
rect 192693 27168 193157 27464
rect 193453 27168 193917 27464
rect 194213 27168 194677 27464
rect 194973 27168 195437 27464
rect 195733 27168 196197 27464
rect 196493 27168 196957 27464
rect 197253 27168 197717 27464
rect 198013 27168 198477 27464
rect 198773 27168 199237 27464
rect 199533 27168 199997 27464
rect 200293 27168 200757 27464
rect 201053 27168 201517 27464
rect 201813 27168 202277 27464
rect 202573 27168 203037 27464
rect 203333 27168 203797 27464
rect 204093 27168 204557 27464
rect 204853 27168 205317 27464
rect 205613 27168 206077 27464
rect 206373 27168 206837 27464
rect 207133 27168 207597 27464
rect 207893 27168 208357 27464
rect 208653 27168 209117 27464
rect 209413 27168 209877 27464
rect 210173 27168 210637 27464
rect 210933 27168 211505 27464
rect 186505 26704 211505 27168
rect 186505 26408 187077 26704
rect 187373 26408 187837 26704
rect 188133 26408 188597 26704
rect 188893 26408 189357 26704
rect 189653 26408 190117 26704
rect 190413 26408 190877 26704
rect 191173 26408 191637 26704
rect 191933 26408 192397 26704
rect 192693 26408 193157 26704
rect 193453 26408 193917 26704
rect 194213 26408 194677 26704
rect 194973 26408 195437 26704
rect 195733 26408 196197 26704
rect 196493 26408 196957 26704
rect 197253 26408 197717 26704
rect 198013 26408 198477 26704
rect 198773 26408 199237 26704
rect 199533 26408 199997 26704
rect 200293 26408 200757 26704
rect 201053 26408 201517 26704
rect 201813 26408 202277 26704
rect 202573 26408 203037 26704
rect 203333 26408 203797 26704
rect 204093 26408 204557 26704
rect 204853 26408 205317 26704
rect 205613 26408 206077 26704
rect 206373 26408 206837 26704
rect 207133 26408 207597 26704
rect 207893 26408 208357 26704
rect 208653 26408 209117 26704
rect 209413 26408 209877 26704
rect 210173 26408 210637 26704
rect 210933 26408 211505 26704
rect 186505 25944 211505 26408
rect 186505 25648 187077 25944
rect 187373 25648 187837 25944
rect 188133 25648 188597 25944
rect 188893 25648 189357 25944
rect 189653 25648 190117 25944
rect 190413 25648 190877 25944
rect 191173 25648 191637 25944
rect 191933 25648 192397 25944
rect 192693 25648 193157 25944
rect 193453 25648 193917 25944
rect 194213 25648 194677 25944
rect 194973 25648 195437 25944
rect 195733 25648 196197 25944
rect 196493 25648 196957 25944
rect 197253 25648 197717 25944
rect 198013 25648 198477 25944
rect 198773 25648 199237 25944
rect 199533 25648 199997 25944
rect 200293 25648 200757 25944
rect 201053 25648 201517 25944
rect 201813 25648 202277 25944
rect 202573 25648 203037 25944
rect 203333 25648 203797 25944
rect 204093 25648 204557 25944
rect 204853 25648 205317 25944
rect 205613 25648 206077 25944
rect 206373 25648 206837 25944
rect 207133 25648 207597 25944
rect 207893 25648 208357 25944
rect 208653 25648 209117 25944
rect 209413 25648 209877 25944
rect 210173 25648 210637 25944
rect 210933 25648 211505 25944
rect 186505 25184 211505 25648
rect 186505 24888 187077 25184
rect 187373 24888 187837 25184
rect 188133 24888 188597 25184
rect 188893 24888 189357 25184
rect 189653 24888 190117 25184
rect 190413 24888 190877 25184
rect 191173 24888 191637 25184
rect 191933 24888 192397 25184
rect 192693 24888 193157 25184
rect 193453 24888 193917 25184
rect 194213 24888 194677 25184
rect 194973 24888 195437 25184
rect 195733 24888 196197 25184
rect 196493 24888 196957 25184
rect 197253 24888 197717 25184
rect 198013 24888 198477 25184
rect 198773 24888 199237 25184
rect 199533 24888 199997 25184
rect 200293 24888 200757 25184
rect 201053 24888 201517 25184
rect 201813 24888 202277 25184
rect 202573 24888 203037 25184
rect 203333 24888 203797 25184
rect 204093 24888 204557 25184
rect 204853 24888 205317 25184
rect 205613 24888 206077 25184
rect 206373 24888 206837 25184
rect 207133 24888 207597 25184
rect 207893 24888 208357 25184
rect 208653 24888 209117 25184
rect 209413 24888 209877 25184
rect 210173 24888 210637 25184
rect 210933 24888 211505 25184
rect 186505 24424 211505 24888
rect 186505 24128 187077 24424
rect 187373 24128 187837 24424
rect 188133 24128 188597 24424
rect 188893 24128 189357 24424
rect 189653 24128 190117 24424
rect 190413 24128 190877 24424
rect 191173 24128 191637 24424
rect 191933 24128 192397 24424
rect 192693 24128 193157 24424
rect 193453 24128 193917 24424
rect 194213 24128 194677 24424
rect 194973 24128 195437 24424
rect 195733 24128 196197 24424
rect 196493 24128 196957 24424
rect 197253 24128 197717 24424
rect 198013 24128 198477 24424
rect 198773 24128 199237 24424
rect 199533 24128 199997 24424
rect 200293 24128 200757 24424
rect 201053 24128 201517 24424
rect 201813 24128 202277 24424
rect 202573 24128 203037 24424
rect 203333 24128 203797 24424
rect 204093 24128 204557 24424
rect 204853 24128 205317 24424
rect 205613 24128 206077 24424
rect 206373 24128 206837 24424
rect 207133 24128 207597 24424
rect 207893 24128 208357 24424
rect 208653 24128 209117 24424
rect 209413 24128 209877 24424
rect 210173 24128 210637 24424
rect 210933 24128 211505 24424
rect 186505 23664 211505 24128
rect 186505 23368 187077 23664
rect 187373 23368 187837 23664
rect 188133 23368 188597 23664
rect 188893 23368 189357 23664
rect 189653 23368 190117 23664
rect 190413 23368 190877 23664
rect 191173 23368 191637 23664
rect 191933 23368 192397 23664
rect 192693 23368 193157 23664
rect 193453 23368 193917 23664
rect 194213 23368 194677 23664
rect 194973 23368 195437 23664
rect 195733 23368 196197 23664
rect 196493 23368 196957 23664
rect 197253 23368 197717 23664
rect 198013 23368 198477 23664
rect 198773 23368 199237 23664
rect 199533 23368 199997 23664
rect 200293 23368 200757 23664
rect 201053 23368 201517 23664
rect 201813 23368 202277 23664
rect 202573 23368 203037 23664
rect 203333 23368 203797 23664
rect 204093 23368 204557 23664
rect 204853 23368 205317 23664
rect 205613 23368 206077 23664
rect 206373 23368 206837 23664
rect 207133 23368 207597 23664
rect 207893 23368 208357 23664
rect 208653 23368 209117 23664
rect 209413 23368 209877 23664
rect 210173 23368 210637 23664
rect 210933 23368 211505 23664
rect 186505 22904 211505 23368
rect 186505 22608 187077 22904
rect 187373 22608 187837 22904
rect 188133 22608 188597 22904
rect 188893 22608 189357 22904
rect 189653 22608 190117 22904
rect 190413 22608 190877 22904
rect 191173 22608 191637 22904
rect 191933 22608 192397 22904
rect 192693 22608 193157 22904
rect 193453 22608 193917 22904
rect 194213 22608 194677 22904
rect 194973 22608 195437 22904
rect 195733 22608 196197 22904
rect 196493 22608 196957 22904
rect 197253 22608 197717 22904
rect 198013 22608 198477 22904
rect 198773 22608 199237 22904
rect 199533 22608 199997 22904
rect 200293 22608 200757 22904
rect 201053 22608 201517 22904
rect 201813 22608 202277 22904
rect 202573 22608 203037 22904
rect 203333 22608 203797 22904
rect 204093 22608 204557 22904
rect 204853 22608 205317 22904
rect 205613 22608 206077 22904
rect 206373 22608 206837 22904
rect 207133 22608 207597 22904
rect 207893 22608 208357 22904
rect 208653 22608 209117 22904
rect 209413 22608 209877 22904
rect 210173 22608 210637 22904
rect 210933 22608 211505 22904
rect 186505 22144 211505 22608
rect 186505 21848 187077 22144
rect 187373 21848 187837 22144
rect 188133 21848 188597 22144
rect 188893 21848 189357 22144
rect 189653 21848 190117 22144
rect 190413 21848 190877 22144
rect 191173 21848 191637 22144
rect 191933 21848 192397 22144
rect 192693 21848 193157 22144
rect 193453 21848 193917 22144
rect 194213 21848 194677 22144
rect 194973 21848 195437 22144
rect 195733 21848 196197 22144
rect 196493 21848 196957 22144
rect 197253 21848 197717 22144
rect 198013 21848 198477 22144
rect 198773 21848 199237 22144
rect 199533 21848 199997 22144
rect 200293 21848 200757 22144
rect 201053 21848 201517 22144
rect 201813 21848 202277 22144
rect 202573 21848 203037 22144
rect 203333 21848 203797 22144
rect 204093 21848 204557 22144
rect 204853 21848 205317 22144
rect 205613 21848 206077 22144
rect 206373 21848 206837 22144
rect 207133 21848 207597 22144
rect 207893 21848 208357 22144
rect 208653 21848 209117 22144
rect 209413 21848 209877 22144
rect 210173 21848 210637 22144
rect 210933 21848 211505 22144
rect 186505 21384 211505 21848
rect 186505 21088 187077 21384
rect 187373 21088 187837 21384
rect 188133 21088 188597 21384
rect 188893 21088 189357 21384
rect 189653 21088 190117 21384
rect 190413 21088 190877 21384
rect 191173 21088 191637 21384
rect 191933 21088 192397 21384
rect 192693 21088 193157 21384
rect 193453 21088 193917 21384
rect 194213 21088 194677 21384
rect 194973 21088 195437 21384
rect 195733 21088 196197 21384
rect 196493 21088 196957 21384
rect 197253 21088 197717 21384
rect 198013 21088 198477 21384
rect 198773 21088 199237 21384
rect 199533 21088 199997 21384
rect 200293 21088 200757 21384
rect 201053 21088 201517 21384
rect 201813 21088 202277 21384
rect 202573 21088 203037 21384
rect 203333 21088 203797 21384
rect 204093 21088 204557 21384
rect 204853 21088 205317 21384
rect 205613 21088 206077 21384
rect 206373 21088 206837 21384
rect 207133 21088 207597 21384
rect 207893 21088 208357 21384
rect 208653 21088 209117 21384
rect 209413 21088 209877 21384
rect 210173 21088 210637 21384
rect 210933 21088 211505 21384
rect 186505 20624 211505 21088
rect 186505 20328 187077 20624
rect 187373 20328 187837 20624
rect 188133 20328 188597 20624
rect 188893 20328 189357 20624
rect 189653 20328 190117 20624
rect 190413 20328 190877 20624
rect 191173 20328 191637 20624
rect 191933 20328 192397 20624
rect 192693 20328 193157 20624
rect 193453 20328 193917 20624
rect 194213 20328 194677 20624
rect 194973 20328 195437 20624
rect 195733 20328 196197 20624
rect 196493 20328 196957 20624
rect 197253 20328 197717 20624
rect 198013 20328 198477 20624
rect 198773 20328 199237 20624
rect 199533 20328 199997 20624
rect 200293 20328 200757 20624
rect 201053 20328 201517 20624
rect 201813 20328 202277 20624
rect 202573 20328 203037 20624
rect 203333 20328 203797 20624
rect 204093 20328 204557 20624
rect 204853 20328 205317 20624
rect 205613 20328 206077 20624
rect 206373 20328 206837 20624
rect 207133 20328 207597 20624
rect 207893 20328 208357 20624
rect 208653 20328 209117 20624
rect 209413 20328 209877 20624
rect 210173 20328 210637 20624
rect 210933 20328 211505 20624
rect 186505 19864 211505 20328
rect 186505 19568 187077 19864
rect 187373 19568 187837 19864
rect 188133 19568 188597 19864
rect 188893 19568 189357 19864
rect 189653 19568 190117 19864
rect 190413 19568 190877 19864
rect 191173 19568 191637 19864
rect 191933 19568 192397 19864
rect 192693 19568 193157 19864
rect 193453 19568 193917 19864
rect 194213 19568 194677 19864
rect 194973 19568 195437 19864
rect 195733 19568 196197 19864
rect 196493 19568 196957 19864
rect 197253 19568 197717 19864
rect 198013 19568 198477 19864
rect 198773 19568 199237 19864
rect 199533 19568 199997 19864
rect 200293 19568 200757 19864
rect 201053 19568 201517 19864
rect 201813 19568 202277 19864
rect 202573 19568 203037 19864
rect 203333 19568 203797 19864
rect 204093 19568 204557 19864
rect 204853 19568 205317 19864
rect 205613 19568 206077 19864
rect 206373 19568 206837 19864
rect 207133 19568 207597 19864
rect 207893 19568 208357 19864
rect 208653 19568 209117 19864
rect 209413 19568 209877 19864
rect 210173 19568 210637 19864
rect 210933 19568 211505 19864
rect 186505 19104 211505 19568
rect 186505 18808 187077 19104
rect 187373 18808 187837 19104
rect 188133 18808 188597 19104
rect 188893 18808 189357 19104
rect 189653 18808 190117 19104
rect 190413 18808 190877 19104
rect 191173 18808 191637 19104
rect 191933 18808 192397 19104
rect 192693 18808 193157 19104
rect 193453 18808 193917 19104
rect 194213 18808 194677 19104
rect 194973 18808 195437 19104
rect 195733 18808 196197 19104
rect 196493 18808 196957 19104
rect 197253 18808 197717 19104
rect 198013 18808 198477 19104
rect 198773 18808 199237 19104
rect 199533 18808 199997 19104
rect 200293 18808 200757 19104
rect 201053 18808 201517 19104
rect 201813 18808 202277 19104
rect 202573 18808 203037 19104
rect 203333 18808 203797 19104
rect 204093 18808 204557 19104
rect 204853 18808 205317 19104
rect 205613 18808 206077 19104
rect 206373 18808 206837 19104
rect 207133 18808 207597 19104
rect 207893 18808 208357 19104
rect 208653 18808 209117 19104
rect 209413 18808 209877 19104
rect 210173 18808 210637 19104
rect 210933 18808 211505 19104
rect 186505 18344 211505 18808
rect 186505 18048 187077 18344
rect 187373 18048 187837 18344
rect 188133 18048 188597 18344
rect 188893 18048 189357 18344
rect 189653 18048 190117 18344
rect 190413 18048 190877 18344
rect 191173 18048 191637 18344
rect 191933 18048 192397 18344
rect 192693 18048 193157 18344
rect 193453 18048 193917 18344
rect 194213 18048 194677 18344
rect 194973 18048 195437 18344
rect 195733 18048 196197 18344
rect 196493 18048 196957 18344
rect 197253 18048 197717 18344
rect 198013 18048 198477 18344
rect 198773 18048 199237 18344
rect 199533 18048 199997 18344
rect 200293 18048 200757 18344
rect 201053 18048 201517 18344
rect 201813 18048 202277 18344
rect 202573 18048 203037 18344
rect 203333 18048 203797 18344
rect 204093 18048 204557 18344
rect 204853 18048 205317 18344
rect 205613 18048 206077 18344
rect 206373 18048 206837 18344
rect 207133 18048 207597 18344
rect 207893 18048 208357 18344
rect 208653 18048 209117 18344
rect 209413 18048 209877 18344
rect 210173 18048 210637 18344
rect 210933 18048 211505 18344
rect 186505 17584 211505 18048
rect 186505 17288 187077 17584
rect 187373 17288 187837 17584
rect 188133 17288 188597 17584
rect 188893 17288 189357 17584
rect 189653 17288 190117 17584
rect 190413 17288 190877 17584
rect 191173 17288 191637 17584
rect 191933 17288 192397 17584
rect 192693 17288 193157 17584
rect 193453 17288 193917 17584
rect 194213 17288 194677 17584
rect 194973 17288 195437 17584
rect 195733 17288 196197 17584
rect 196493 17288 196957 17584
rect 197253 17288 197717 17584
rect 198013 17288 198477 17584
rect 198773 17288 199237 17584
rect 199533 17288 199997 17584
rect 200293 17288 200757 17584
rect 201053 17288 201517 17584
rect 201813 17288 202277 17584
rect 202573 17288 203037 17584
rect 203333 17288 203797 17584
rect 204093 17288 204557 17584
rect 204853 17288 205317 17584
rect 205613 17288 206077 17584
rect 206373 17288 206837 17584
rect 207133 17288 207597 17584
rect 207893 17288 208357 17584
rect 208653 17288 209117 17584
rect 209413 17288 209877 17584
rect 210173 17288 210637 17584
rect 210933 17288 211505 17584
rect 186505 16824 211505 17288
rect 186505 16528 187077 16824
rect 187373 16528 187837 16824
rect 188133 16528 188597 16824
rect 188893 16528 189357 16824
rect 189653 16528 190117 16824
rect 190413 16528 190877 16824
rect 191173 16528 191637 16824
rect 191933 16528 192397 16824
rect 192693 16528 193157 16824
rect 193453 16528 193917 16824
rect 194213 16528 194677 16824
rect 194973 16528 195437 16824
rect 195733 16528 196197 16824
rect 196493 16528 196957 16824
rect 197253 16528 197717 16824
rect 198013 16528 198477 16824
rect 198773 16528 199237 16824
rect 199533 16528 199997 16824
rect 200293 16528 200757 16824
rect 201053 16528 201517 16824
rect 201813 16528 202277 16824
rect 202573 16528 203037 16824
rect 203333 16528 203797 16824
rect 204093 16528 204557 16824
rect 204853 16528 205317 16824
rect 205613 16528 206077 16824
rect 206373 16528 206837 16824
rect 207133 16528 207597 16824
rect 207893 16528 208357 16824
rect 208653 16528 209117 16824
rect 209413 16528 209877 16824
rect 210173 16528 210637 16824
rect 210933 16528 211505 16824
rect 186505 16064 211505 16528
rect 186505 15768 187077 16064
rect 187373 15768 187837 16064
rect 188133 15768 188597 16064
rect 188893 15768 189357 16064
rect 189653 15768 190117 16064
rect 190413 15768 190877 16064
rect 191173 15768 191637 16064
rect 191933 15768 192397 16064
rect 192693 15768 193157 16064
rect 193453 15768 193917 16064
rect 194213 15768 194677 16064
rect 194973 15768 195437 16064
rect 195733 15768 196197 16064
rect 196493 15768 196957 16064
rect 197253 15768 197717 16064
rect 198013 15768 198477 16064
rect 198773 15768 199237 16064
rect 199533 15768 199997 16064
rect 200293 15768 200757 16064
rect 201053 15768 201517 16064
rect 201813 15768 202277 16064
rect 202573 15768 203037 16064
rect 203333 15768 203797 16064
rect 204093 15768 204557 16064
rect 204853 15768 205317 16064
rect 205613 15768 206077 16064
rect 206373 15768 206837 16064
rect 207133 15768 207597 16064
rect 207893 15768 208357 16064
rect 208653 15768 209117 16064
rect 209413 15768 209877 16064
rect 210173 15768 210637 16064
rect 210933 15768 211505 16064
rect 186505 15304 211505 15768
rect 186505 15008 187077 15304
rect 187373 15008 187837 15304
rect 188133 15008 188597 15304
rect 188893 15008 189357 15304
rect 189653 15008 190117 15304
rect 190413 15008 190877 15304
rect 191173 15008 191637 15304
rect 191933 15008 192397 15304
rect 192693 15008 193157 15304
rect 193453 15008 193917 15304
rect 194213 15008 194677 15304
rect 194973 15008 195437 15304
rect 195733 15008 196197 15304
rect 196493 15008 196957 15304
rect 197253 15008 197717 15304
rect 198013 15008 198477 15304
rect 198773 15008 199237 15304
rect 199533 15008 199997 15304
rect 200293 15008 200757 15304
rect 201053 15008 201517 15304
rect 201813 15008 202277 15304
rect 202573 15008 203037 15304
rect 203333 15008 203797 15304
rect 204093 15008 204557 15304
rect 204853 15008 205317 15304
rect 205613 15008 206077 15304
rect 206373 15008 206837 15304
rect 207133 15008 207597 15304
rect 207893 15008 208357 15304
rect 208653 15008 209117 15304
rect 209413 15008 209877 15304
rect 210173 15008 210637 15304
rect 210933 15008 211505 15304
rect 186505 14544 211505 15008
rect 186505 14248 187077 14544
rect 187373 14248 187837 14544
rect 188133 14248 188597 14544
rect 188893 14248 189357 14544
rect 189653 14248 190117 14544
rect 190413 14248 190877 14544
rect 191173 14248 191637 14544
rect 191933 14248 192397 14544
rect 192693 14248 193157 14544
rect 193453 14248 193917 14544
rect 194213 14248 194677 14544
rect 194973 14248 195437 14544
rect 195733 14248 196197 14544
rect 196493 14248 196957 14544
rect 197253 14248 197717 14544
rect 198013 14248 198477 14544
rect 198773 14248 199237 14544
rect 199533 14248 199997 14544
rect 200293 14248 200757 14544
rect 201053 14248 201517 14544
rect 201813 14248 202277 14544
rect 202573 14248 203037 14544
rect 203333 14248 203797 14544
rect 204093 14248 204557 14544
rect 204853 14248 205317 14544
rect 205613 14248 206077 14544
rect 206373 14248 206837 14544
rect 207133 14248 207597 14544
rect 207893 14248 208357 14544
rect 208653 14248 209117 14544
rect 209413 14248 209877 14544
rect 210173 14248 210637 14544
rect 210933 14248 211505 14544
rect 186505 13784 211505 14248
rect 186505 13488 187077 13784
rect 187373 13488 187837 13784
rect 188133 13488 188597 13784
rect 188893 13488 189357 13784
rect 189653 13488 190117 13784
rect 190413 13488 190877 13784
rect 191173 13488 191637 13784
rect 191933 13488 192397 13784
rect 192693 13488 193157 13784
rect 193453 13488 193917 13784
rect 194213 13488 194677 13784
rect 194973 13488 195437 13784
rect 195733 13488 196197 13784
rect 196493 13488 196957 13784
rect 197253 13488 197717 13784
rect 198013 13488 198477 13784
rect 198773 13488 199237 13784
rect 199533 13488 199997 13784
rect 200293 13488 200757 13784
rect 201053 13488 201517 13784
rect 201813 13488 202277 13784
rect 202573 13488 203037 13784
rect 203333 13488 203797 13784
rect 204093 13488 204557 13784
rect 204853 13488 205317 13784
rect 205613 13488 206077 13784
rect 206373 13488 206837 13784
rect 207133 13488 207597 13784
rect 207893 13488 208357 13784
rect 208653 13488 209117 13784
rect 209413 13488 209877 13784
rect 210173 13488 210637 13784
rect 210933 13488 211505 13784
rect 186505 13024 211505 13488
rect 186505 12728 187077 13024
rect 187373 12728 187837 13024
rect 188133 12728 188597 13024
rect 188893 12728 189357 13024
rect 189653 12728 190117 13024
rect 190413 12728 190877 13024
rect 191173 12728 191637 13024
rect 191933 12728 192397 13024
rect 192693 12728 193157 13024
rect 193453 12728 193917 13024
rect 194213 12728 194677 13024
rect 194973 12728 195437 13024
rect 195733 12728 196197 13024
rect 196493 12728 196957 13024
rect 197253 12728 197717 13024
rect 198013 12728 198477 13024
rect 198773 12728 199237 13024
rect 199533 12728 199997 13024
rect 200293 12728 200757 13024
rect 201053 12728 201517 13024
rect 201813 12728 202277 13024
rect 202573 12728 203037 13024
rect 203333 12728 203797 13024
rect 204093 12728 204557 13024
rect 204853 12728 205317 13024
rect 205613 12728 206077 13024
rect 206373 12728 206837 13024
rect 207133 12728 207597 13024
rect 207893 12728 208357 13024
rect 208653 12728 209117 13024
rect 209413 12728 209877 13024
rect 210173 12728 210637 13024
rect 210933 12728 211505 13024
rect 186505 12264 211505 12728
rect 186505 11968 187077 12264
rect 187373 11968 187837 12264
rect 188133 11968 188597 12264
rect 188893 11968 189357 12264
rect 189653 11968 190117 12264
rect 190413 11968 190877 12264
rect 191173 11968 191637 12264
rect 191933 11968 192397 12264
rect 192693 11968 193157 12264
rect 193453 11968 193917 12264
rect 194213 11968 194677 12264
rect 194973 11968 195437 12264
rect 195733 11968 196197 12264
rect 196493 11968 196957 12264
rect 197253 11968 197717 12264
rect 198013 11968 198477 12264
rect 198773 11968 199237 12264
rect 199533 11968 199997 12264
rect 200293 11968 200757 12264
rect 201053 11968 201517 12264
rect 201813 11968 202277 12264
rect 202573 11968 203037 12264
rect 203333 11968 203797 12264
rect 204093 11968 204557 12264
rect 204853 11968 205317 12264
rect 205613 11968 206077 12264
rect 206373 11968 206837 12264
rect 207133 11968 207597 12264
rect 207893 11968 208357 12264
rect 208653 11968 209117 12264
rect 209413 11968 209877 12264
rect 210173 11968 210637 12264
rect 210933 11968 211505 12264
rect 186505 11504 211505 11968
rect 186505 11208 187077 11504
rect 187373 11208 187837 11504
rect 188133 11208 188597 11504
rect 188893 11208 189357 11504
rect 189653 11208 190117 11504
rect 190413 11208 190877 11504
rect 191173 11208 191637 11504
rect 191933 11208 192397 11504
rect 192693 11208 193157 11504
rect 193453 11208 193917 11504
rect 194213 11208 194677 11504
rect 194973 11208 195437 11504
rect 195733 11208 196197 11504
rect 196493 11208 196957 11504
rect 197253 11208 197717 11504
rect 198013 11208 198477 11504
rect 198773 11208 199237 11504
rect 199533 11208 199997 11504
rect 200293 11208 200757 11504
rect 201053 11208 201517 11504
rect 201813 11208 202277 11504
rect 202573 11208 203037 11504
rect 203333 11208 203797 11504
rect 204093 11208 204557 11504
rect 204853 11208 205317 11504
rect 205613 11208 206077 11504
rect 206373 11208 206837 11504
rect 207133 11208 207597 11504
rect 207893 11208 208357 11504
rect 208653 11208 209117 11504
rect 209413 11208 209877 11504
rect 210173 11208 210637 11504
rect 210933 11208 211505 11504
rect 186505 10744 211505 11208
rect 186505 10448 187077 10744
rect 187373 10448 187837 10744
rect 188133 10448 188597 10744
rect 188893 10448 189357 10744
rect 189653 10448 190117 10744
rect 190413 10448 190877 10744
rect 191173 10448 191637 10744
rect 191933 10448 192397 10744
rect 192693 10448 193157 10744
rect 193453 10448 193917 10744
rect 194213 10448 194677 10744
rect 194973 10448 195437 10744
rect 195733 10448 196197 10744
rect 196493 10448 196957 10744
rect 197253 10448 197717 10744
rect 198013 10448 198477 10744
rect 198773 10448 199237 10744
rect 199533 10448 199997 10744
rect 200293 10448 200757 10744
rect 201053 10448 201517 10744
rect 201813 10448 202277 10744
rect 202573 10448 203037 10744
rect 203333 10448 203797 10744
rect 204093 10448 204557 10744
rect 204853 10448 205317 10744
rect 205613 10448 206077 10744
rect 206373 10448 206837 10744
rect 207133 10448 207597 10744
rect 207893 10448 208357 10744
rect 208653 10448 209117 10744
rect 209413 10448 209877 10744
rect 210173 10448 210637 10744
rect 210933 10448 211505 10744
rect 186505 9716 211505 10448
<< mimcapcontact >>
rect 114357 30875 114653 31171
rect 115117 30875 115413 31171
rect 115877 30875 116173 31171
rect 116637 30875 116933 31171
rect 117397 30875 117693 31171
rect 118157 30875 118453 31171
rect 118917 30875 119213 31171
rect 119677 30875 119973 31171
rect 120437 30875 120733 31171
rect 121197 30875 121493 31171
rect 121957 30875 122253 31171
rect 122717 30875 123013 31171
rect 123477 30875 123773 31171
rect 124237 30875 124533 31171
rect 124997 30875 125293 31171
rect 125757 30875 126053 31171
rect 126517 30875 126813 31171
rect 127277 30875 127573 31171
rect 128037 30875 128333 31171
rect 128797 30875 129093 31171
rect 129557 30875 129853 31171
rect 130317 30875 130613 31171
rect 131077 30875 131373 31171
rect 131837 30875 132133 31171
rect 132597 30875 132893 31171
rect 114357 30115 114653 30411
rect 115117 30115 115413 30411
rect 115877 30115 116173 30411
rect 116637 30115 116933 30411
rect 117397 30115 117693 30411
rect 118157 30115 118453 30411
rect 118917 30115 119213 30411
rect 119677 30115 119973 30411
rect 120437 30115 120733 30411
rect 121197 30115 121493 30411
rect 121957 30115 122253 30411
rect 122717 30115 123013 30411
rect 123477 30115 123773 30411
rect 124237 30115 124533 30411
rect 124997 30115 125293 30411
rect 125757 30115 126053 30411
rect 126517 30115 126813 30411
rect 127277 30115 127573 30411
rect 128037 30115 128333 30411
rect 128797 30115 129093 30411
rect 129557 30115 129853 30411
rect 130317 30115 130613 30411
rect 131077 30115 131373 30411
rect 131837 30115 132133 30411
rect 132597 30115 132893 30411
rect 114357 29355 114653 29651
rect 115117 29355 115413 29651
rect 115877 29355 116173 29651
rect 116637 29355 116933 29651
rect 117397 29355 117693 29651
rect 118157 29355 118453 29651
rect 118917 29355 119213 29651
rect 119677 29355 119973 29651
rect 120437 29355 120733 29651
rect 121197 29355 121493 29651
rect 121957 29355 122253 29651
rect 122717 29355 123013 29651
rect 123477 29355 123773 29651
rect 124237 29355 124533 29651
rect 124997 29355 125293 29651
rect 125757 29355 126053 29651
rect 126517 29355 126813 29651
rect 127277 29355 127573 29651
rect 128037 29355 128333 29651
rect 128797 29355 129093 29651
rect 129557 29355 129853 29651
rect 130317 29355 130613 29651
rect 131077 29355 131373 29651
rect 131837 29355 132133 29651
rect 132597 29355 132893 29651
rect 114357 28595 114653 28891
rect 115117 28595 115413 28891
rect 115877 28595 116173 28891
rect 116637 28595 116933 28891
rect 117397 28595 117693 28891
rect 118157 28595 118453 28891
rect 118917 28595 119213 28891
rect 119677 28595 119973 28891
rect 120437 28595 120733 28891
rect 121197 28595 121493 28891
rect 121957 28595 122253 28891
rect 122717 28595 123013 28891
rect 123477 28595 123773 28891
rect 124237 28595 124533 28891
rect 124997 28595 125293 28891
rect 125757 28595 126053 28891
rect 126517 28595 126813 28891
rect 127277 28595 127573 28891
rect 128037 28595 128333 28891
rect 128797 28595 129093 28891
rect 129557 28595 129853 28891
rect 130317 28595 130613 28891
rect 131077 28595 131373 28891
rect 131837 28595 132133 28891
rect 132597 28595 132893 28891
rect 114357 27835 114653 28131
rect 115117 27835 115413 28131
rect 115877 27835 116173 28131
rect 116637 27835 116933 28131
rect 117397 27835 117693 28131
rect 118157 27835 118453 28131
rect 118917 27835 119213 28131
rect 119677 27835 119973 28131
rect 120437 27835 120733 28131
rect 121197 27835 121493 28131
rect 121957 27835 122253 28131
rect 122717 27835 123013 28131
rect 123477 27835 123773 28131
rect 124237 27835 124533 28131
rect 124997 27835 125293 28131
rect 125757 27835 126053 28131
rect 126517 27835 126813 28131
rect 127277 27835 127573 28131
rect 128037 27835 128333 28131
rect 128797 27835 129093 28131
rect 129557 27835 129853 28131
rect 130317 27835 130613 28131
rect 131077 27835 131373 28131
rect 131837 27835 132133 28131
rect 132597 27835 132893 28131
rect 114357 27075 114653 27371
rect 115117 27075 115413 27371
rect 115877 27075 116173 27371
rect 116637 27075 116933 27371
rect 117397 27075 117693 27371
rect 118157 27075 118453 27371
rect 118917 27075 119213 27371
rect 119677 27075 119973 27371
rect 120437 27075 120733 27371
rect 121197 27075 121493 27371
rect 121957 27075 122253 27371
rect 122717 27075 123013 27371
rect 123477 27075 123773 27371
rect 124237 27075 124533 27371
rect 124997 27075 125293 27371
rect 125757 27075 126053 27371
rect 126517 27075 126813 27371
rect 127277 27075 127573 27371
rect 128037 27075 128333 27371
rect 128797 27075 129093 27371
rect 129557 27075 129853 27371
rect 130317 27075 130613 27371
rect 131077 27075 131373 27371
rect 131837 27075 132133 27371
rect 132597 27075 132893 27371
rect 114357 26315 114653 26611
rect 115117 26315 115413 26611
rect 115877 26315 116173 26611
rect 116637 26315 116933 26611
rect 117397 26315 117693 26611
rect 118157 26315 118453 26611
rect 118917 26315 119213 26611
rect 119677 26315 119973 26611
rect 120437 26315 120733 26611
rect 121197 26315 121493 26611
rect 121957 26315 122253 26611
rect 122717 26315 123013 26611
rect 123477 26315 123773 26611
rect 124237 26315 124533 26611
rect 124997 26315 125293 26611
rect 125757 26315 126053 26611
rect 126517 26315 126813 26611
rect 127277 26315 127573 26611
rect 128037 26315 128333 26611
rect 128797 26315 129093 26611
rect 129557 26315 129853 26611
rect 130317 26315 130613 26611
rect 131077 26315 131373 26611
rect 131837 26315 132133 26611
rect 132597 26315 132893 26611
rect 114357 25555 114653 25851
rect 115117 25555 115413 25851
rect 115877 25555 116173 25851
rect 116637 25555 116933 25851
rect 117397 25555 117693 25851
rect 118157 25555 118453 25851
rect 118917 25555 119213 25851
rect 119677 25555 119973 25851
rect 120437 25555 120733 25851
rect 121197 25555 121493 25851
rect 121957 25555 122253 25851
rect 122717 25555 123013 25851
rect 123477 25555 123773 25851
rect 124237 25555 124533 25851
rect 124997 25555 125293 25851
rect 125757 25555 126053 25851
rect 126517 25555 126813 25851
rect 127277 25555 127573 25851
rect 128037 25555 128333 25851
rect 128797 25555 129093 25851
rect 129557 25555 129853 25851
rect 130317 25555 130613 25851
rect 131077 25555 131373 25851
rect 131837 25555 132133 25851
rect 132597 25555 132893 25851
rect 114357 24795 114653 25091
rect 115117 24795 115413 25091
rect 115877 24795 116173 25091
rect 116637 24795 116933 25091
rect 117397 24795 117693 25091
rect 118157 24795 118453 25091
rect 118917 24795 119213 25091
rect 119677 24795 119973 25091
rect 120437 24795 120733 25091
rect 121197 24795 121493 25091
rect 121957 24795 122253 25091
rect 122717 24795 123013 25091
rect 123477 24795 123773 25091
rect 124237 24795 124533 25091
rect 124997 24795 125293 25091
rect 125757 24795 126053 25091
rect 126517 24795 126813 25091
rect 127277 24795 127573 25091
rect 128037 24795 128333 25091
rect 128797 24795 129093 25091
rect 129557 24795 129853 25091
rect 130317 24795 130613 25091
rect 131077 24795 131373 25091
rect 131837 24795 132133 25091
rect 132597 24795 132893 25091
rect 114357 24035 114653 24331
rect 115117 24035 115413 24331
rect 115877 24035 116173 24331
rect 116637 24035 116933 24331
rect 117397 24035 117693 24331
rect 118157 24035 118453 24331
rect 118917 24035 119213 24331
rect 119677 24035 119973 24331
rect 120437 24035 120733 24331
rect 121197 24035 121493 24331
rect 121957 24035 122253 24331
rect 122717 24035 123013 24331
rect 123477 24035 123773 24331
rect 124237 24035 124533 24331
rect 124997 24035 125293 24331
rect 125757 24035 126053 24331
rect 126517 24035 126813 24331
rect 127277 24035 127573 24331
rect 128037 24035 128333 24331
rect 128797 24035 129093 24331
rect 129557 24035 129853 24331
rect 130317 24035 130613 24331
rect 131077 24035 131373 24331
rect 131837 24035 132133 24331
rect 132597 24035 132893 24331
rect 114357 23275 114653 23571
rect 115117 23275 115413 23571
rect 115877 23275 116173 23571
rect 116637 23275 116933 23571
rect 117397 23275 117693 23571
rect 118157 23275 118453 23571
rect 118917 23275 119213 23571
rect 119677 23275 119973 23571
rect 120437 23275 120733 23571
rect 121197 23275 121493 23571
rect 121957 23275 122253 23571
rect 122717 23275 123013 23571
rect 123477 23275 123773 23571
rect 124237 23275 124533 23571
rect 124997 23275 125293 23571
rect 125757 23275 126053 23571
rect 126517 23275 126813 23571
rect 127277 23275 127573 23571
rect 128037 23275 128333 23571
rect 128797 23275 129093 23571
rect 129557 23275 129853 23571
rect 130317 23275 130613 23571
rect 131077 23275 131373 23571
rect 131837 23275 132133 23571
rect 132597 23275 132893 23571
rect 114357 22515 114653 22811
rect 115117 22515 115413 22811
rect 115877 22515 116173 22811
rect 116637 22515 116933 22811
rect 117397 22515 117693 22811
rect 118157 22515 118453 22811
rect 118917 22515 119213 22811
rect 119677 22515 119973 22811
rect 120437 22515 120733 22811
rect 121197 22515 121493 22811
rect 121957 22515 122253 22811
rect 122717 22515 123013 22811
rect 123477 22515 123773 22811
rect 124237 22515 124533 22811
rect 124997 22515 125293 22811
rect 125757 22515 126053 22811
rect 126517 22515 126813 22811
rect 127277 22515 127573 22811
rect 128037 22515 128333 22811
rect 128797 22515 129093 22811
rect 129557 22515 129853 22811
rect 130317 22515 130613 22811
rect 131077 22515 131373 22811
rect 131837 22515 132133 22811
rect 132597 22515 132893 22811
rect 114357 21755 114653 22051
rect 115117 21755 115413 22051
rect 115877 21755 116173 22051
rect 116637 21755 116933 22051
rect 117397 21755 117693 22051
rect 118157 21755 118453 22051
rect 118917 21755 119213 22051
rect 119677 21755 119973 22051
rect 120437 21755 120733 22051
rect 121197 21755 121493 22051
rect 121957 21755 122253 22051
rect 122717 21755 123013 22051
rect 123477 21755 123773 22051
rect 124237 21755 124533 22051
rect 124997 21755 125293 22051
rect 125757 21755 126053 22051
rect 126517 21755 126813 22051
rect 127277 21755 127573 22051
rect 128037 21755 128333 22051
rect 128797 21755 129093 22051
rect 129557 21755 129853 22051
rect 130317 21755 130613 22051
rect 131077 21755 131373 22051
rect 131837 21755 132133 22051
rect 132597 21755 132893 22051
rect 114357 20995 114653 21291
rect 115117 20995 115413 21291
rect 115877 20995 116173 21291
rect 116637 20995 116933 21291
rect 117397 20995 117693 21291
rect 118157 20995 118453 21291
rect 118917 20995 119213 21291
rect 119677 20995 119973 21291
rect 120437 20995 120733 21291
rect 121197 20995 121493 21291
rect 121957 20995 122253 21291
rect 122717 20995 123013 21291
rect 123477 20995 123773 21291
rect 124237 20995 124533 21291
rect 124997 20995 125293 21291
rect 125757 20995 126053 21291
rect 126517 20995 126813 21291
rect 127277 20995 127573 21291
rect 128037 20995 128333 21291
rect 128797 20995 129093 21291
rect 129557 20995 129853 21291
rect 130317 20995 130613 21291
rect 131077 20995 131373 21291
rect 131837 20995 132133 21291
rect 132597 20995 132893 21291
rect 114357 20235 114653 20531
rect 115117 20235 115413 20531
rect 115877 20235 116173 20531
rect 116637 20235 116933 20531
rect 117397 20235 117693 20531
rect 118157 20235 118453 20531
rect 118917 20235 119213 20531
rect 119677 20235 119973 20531
rect 120437 20235 120733 20531
rect 121197 20235 121493 20531
rect 121957 20235 122253 20531
rect 122717 20235 123013 20531
rect 123477 20235 123773 20531
rect 124237 20235 124533 20531
rect 124997 20235 125293 20531
rect 125757 20235 126053 20531
rect 126517 20235 126813 20531
rect 127277 20235 127573 20531
rect 128037 20235 128333 20531
rect 128797 20235 129093 20531
rect 129557 20235 129853 20531
rect 130317 20235 130613 20531
rect 131077 20235 131373 20531
rect 131837 20235 132133 20531
rect 132597 20235 132893 20531
rect 114357 19475 114653 19771
rect 115117 19475 115413 19771
rect 115877 19475 116173 19771
rect 116637 19475 116933 19771
rect 117397 19475 117693 19771
rect 118157 19475 118453 19771
rect 118917 19475 119213 19771
rect 119677 19475 119973 19771
rect 120437 19475 120733 19771
rect 121197 19475 121493 19771
rect 121957 19475 122253 19771
rect 122717 19475 123013 19771
rect 123477 19475 123773 19771
rect 124237 19475 124533 19771
rect 124997 19475 125293 19771
rect 125757 19475 126053 19771
rect 126517 19475 126813 19771
rect 127277 19475 127573 19771
rect 128037 19475 128333 19771
rect 128797 19475 129093 19771
rect 129557 19475 129853 19771
rect 130317 19475 130613 19771
rect 131077 19475 131373 19771
rect 131837 19475 132133 19771
rect 132597 19475 132893 19771
rect 114357 18715 114653 19011
rect 115117 18715 115413 19011
rect 115877 18715 116173 19011
rect 116637 18715 116933 19011
rect 117397 18715 117693 19011
rect 118157 18715 118453 19011
rect 118917 18715 119213 19011
rect 119677 18715 119973 19011
rect 120437 18715 120733 19011
rect 121197 18715 121493 19011
rect 121957 18715 122253 19011
rect 122717 18715 123013 19011
rect 123477 18715 123773 19011
rect 124237 18715 124533 19011
rect 124997 18715 125293 19011
rect 125757 18715 126053 19011
rect 126517 18715 126813 19011
rect 127277 18715 127573 19011
rect 128037 18715 128333 19011
rect 128797 18715 129093 19011
rect 129557 18715 129853 19011
rect 130317 18715 130613 19011
rect 131077 18715 131373 19011
rect 131837 18715 132133 19011
rect 132597 18715 132893 19011
rect 114357 17955 114653 18251
rect 115117 17955 115413 18251
rect 115877 17955 116173 18251
rect 116637 17955 116933 18251
rect 117397 17955 117693 18251
rect 118157 17955 118453 18251
rect 118917 17955 119213 18251
rect 119677 17955 119973 18251
rect 120437 17955 120733 18251
rect 121197 17955 121493 18251
rect 121957 17955 122253 18251
rect 122717 17955 123013 18251
rect 123477 17955 123773 18251
rect 124237 17955 124533 18251
rect 124997 17955 125293 18251
rect 125757 17955 126053 18251
rect 126517 17955 126813 18251
rect 127277 17955 127573 18251
rect 128037 17955 128333 18251
rect 128797 17955 129093 18251
rect 129557 17955 129853 18251
rect 130317 17955 130613 18251
rect 131077 17955 131373 18251
rect 131837 17955 132133 18251
rect 132597 17955 132893 18251
rect 114357 17195 114653 17491
rect 115117 17195 115413 17491
rect 115877 17195 116173 17491
rect 116637 17195 116933 17491
rect 117397 17195 117693 17491
rect 118157 17195 118453 17491
rect 118917 17195 119213 17491
rect 119677 17195 119973 17491
rect 120437 17195 120733 17491
rect 121197 17195 121493 17491
rect 121957 17195 122253 17491
rect 122717 17195 123013 17491
rect 123477 17195 123773 17491
rect 124237 17195 124533 17491
rect 124997 17195 125293 17491
rect 125757 17195 126053 17491
rect 126517 17195 126813 17491
rect 127277 17195 127573 17491
rect 128037 17195 128333 17491
rect 128797 17195 129093 17491
rect 129557 17195 129853 17491
rect 130317 17195 130613 17491
rect 131077 17195 131373 17491
rect 131837 17195 132133 17491
rect 132597 17195 132893 17491
rect 114357 16435 114653 16731
rect 115117 16435 115413 16731
rect 115877 16435 116173 16731
rect 116637 16435 116933 16731
rect 117397 16435 117693 16731
rect 118157 16435 118453 16731
rect 118917 16435 119213 16731
rect 119677 16435 119973 16731
rect 120437 16435 120733 16731
rect 121197 16435 121493 16731
rect 121957 16435 122253 16731
rect 122717 16435 123013 16731
rect 123477 16435 123773 16731
rect 124237 16435 124533 16731
rect 124997 16435 125293 16731
rect 125757 16435 126053 16731
rect 126517 16435 126813 16731
rect 127277 16435 127573 16731
rect 128037 16435 128333 16731
rect 128797 16435 129093 16731
rect 129557 16435 129853 16731
rect 130317 16435 130613 16731
rect 131077 16435 131373 16731
rect 131837 16435 132133 16731
rect 132597 16435 132893 16731
rect 114357 15675 114653 15971
rect 115117 15675 115413 15971
rect 115877 15675 116173 15971
rect 116637 15675 116933 15971
rect 117397 15675 117693 15971
rect 118157 15675 118453 15971
rect 118917 15675 119213 15971
rect 119677 15675 119973 15971
rect 120437 15675 120733 15971
rect 121197 15675 121493 15971
rect 121957 15675 122253 15971
rect 122717 15675 123013 15971
rect 123477 15675 123773 15971
rect 124237 15675 124533 15971
rect 124997 15675 125293 15971
rect 125757 15675 126053 15971
rect 126517 15675 126813 15971
rect 127277 15675 127573 15971
rect 128037 15675 128333 15971
rect 128797 15675 129093 15971
rect 129557 15675 129853 15971
rect 130317 15675 130613 15971
rect 131077 15675 131373 15971
rect 131837 15675 132133 15971
rect 132597 15675 132893 15971
rect 114357 14915 114653 15211
rect 115117 14915 115413 15211
rect 115877 14915 116173 15211
rect 116637 14915 116933 15211
rect 117397 14915 117693 15211
rect 118157 14915 118453 15211
rect 118917 14915 119213 15211
rect 119677 14915 119973 15211
rect 120437 14915 120733 15211
rect 121197 14915 121493 15211
rect 121957 14915 122253 15211
rect 122717 14915 123013 15211
rect 123477 14915 123773 15211
rect 124237 14915 124533 15211
rect 124997 14915 125293 15211
rect 125757 14915 126053 15211
rect 126517 14915 126813 15211
rect 127277 14915 127573 15211
rect 128037 14915 128333 15211
rect 128797 14915 129093 15211
rect 129557 14915 129853 15211
rect 130317 14915 130613 15211
rect 131077 14915 131373 15211
rect 131837 14915 132133 15211
rect 132597 14915 132893 15211
rect 114357 14155 114653 14451
rect 115117 14155 115413 14451
rect 115877 14155 116173 14451
rect 116637 14155 116933 14451
rect 117397 14155 117693 14451
rect 118157 14155 118453 14451
rect 118917 14155 119213 14451
rect 119677 14155 119973 14451
rect 120437 14155 120733 14451
rect 121197 14155 121493 14451
rect 121957 14155 122253 14451
rect 122717 14155 123013 14451
rect 123477 14155 123773 14451
rect 124237 14155 124533 14451
rect 124997 14155 125293 14451
rect 125757 14155 126053 14451
rect 126517 14155 126813 14451
rect 127277 14155 127573 14451
rect 128037 14155 128333 14451
rect 128797 14155 129093 14451
rect 129557 14155 129853 14451
rect 130317 14155 130613 14451
rect 131077 14155 131373 14451
rect 131837 14155 132133 14451
rect 132597 14155 132893 14451
rect 114357 13395 114653 13691
rect 115117 13395 115413 13691
rect 115877 13395 116173 13691
rect 116637 13395 116933 13691
rect 117397 13395 117693 13691
rect 118157 13395 118453 13691
rect 118917 13395 119213 13691
rect 119677 13395 119973 13691
rect 120437 13395 120733 13691
rect 121197 13395 121493 13691
rect 121957 13395 122253 13691
rect 122717 13395 123013 13691
rect 123477 13395 123773 13691
rect 124237 13395 124533 13691
rect 124997 13395 125293 13691
rect 125757 13395 126053 13691
rect 126517 13395 126813 13691
rect 127277 13395 127573 13691
rect 128037 13395 128333 13691
rect 128797 13395 129093 13691
rect 129557 13395 129853 13691
rect 130317 13395 130613 13691
rect 131077 13395 131373 13691
rect 131837 13395 132133 13691
rect 132597 13395 132893 13691
rect 114357 12635 114653 12931
rect 115117 12635 115413 12931
rect 115877 12635 116173 12931
rect 116637 12635 116933 12931
rect 117397 12635 117693 12931
rect 118157 12635 118453 12931
rect 118917 12635 119213 12931
rect 119677 12635 119973 12931
rect 120437 12635 120733 12931
rect 121197 12635 121493 12931
rect 121957 12635 122253 12931
rect 122717 12635 123013 12931
rect 123477 12635 123773 12931
rect 124237 12635 124533 12931
rect 124997 12635 125293 12931
rect 125757 12635 126053 12931
rect 126517 12635 126813 12931
rect 127277 12635 127573 12931
rect 128037 12635 128333 12931
rect 128797 12635 129093 12931
rect 129557 12635 129853 12931
rect 130317 12635 130613 12931
rect 131077 12635 131373 12931
rect 131837 12635 132133 12931
rect 132597 12635 132893 12931
rect 114357 11875 114653 12171
rect 115117 11875 115413 12171
rect 115877 11875 116173 12171
rect 116637 11875 116933 12171
rect 117397 11875 117693 12171
rect 118157 11875 118453 12171
rect 118917 11875 119213 12171
rect 119677 11875 119973 12171
rect 120437 11875 120733 12171
rect 121197 11875 121493 12171
rect 121957 11875 122253 12171
rect 122717 11875 123013 12171
rect 123477 11875 123773 12171
rect 124237 11875 124533 12171
rect 124997 11875 125293 12171
rect 125757 11875 126053 12171
rect 126517 11875 126813 12171
rect 127277 11875 127573 12171
rect 128037 11875 128333 12171
rect 128797 11875 129093 12171
rect 129557 11875 129853 12171
rect 130317 11875 130613 12171
rect 131077 11875 131373 12171
rect 131837 11875 132133 12171
rect 132597 11875 132893 12171
rect 114357 11115 114653 11411
rect 115117 11115 115413 11411
rect 115877 11115 116173 11411
rect 116637 11115 116933 11411
rect 117397 11115 117693 11411
rect 118157 11115 118453 11411
rect 118917 11115 119213 11411
rect 119677 11115 119973 11411
rect 120437 11115 120733 11411
rect 121197 11115 121493 11411
rect 121957 11115 122253 11411
rect 122717 11115 123013 11411
rect 123477 11115 123773 11411
rect 124237 11115 124533 11411
rect 124997 11115 125293 11411
rect 125757 11115 126053 11411
rect 126517 11115 126813 11411
rect 127277 11115 127573 11411
rect 128037 11115 128333 11411
rect 128797 11115 129093 11411
rect 129557 11115 129853 11411
rect 130317 11115 130613 11411
rect 131077 11115 131373 11411
rect 131837 11115 132133 11411
rect 132597 11115 132893 11411
rect 114357 10355 114653 10651
rect 115117 10355 115413 10651
rect 115877 10355 116173 10651
rect 116637 10355 116933 10651
rect 117397 10355 117693 10651
rect 118157 10355 118453 10651
rect 118917 10355 119213 10651
rect 119677 10355 119973 10651
rect 120437 10355 120733 10651
rect 121197 10355 121493 10651
rect 121957 10355 122253 10651
rect 122717 10355 123013 10651
rect 123477 10355 123773 10651
rect 124237 10355 124533 10651
rect 124997 10355 125293 10651
rect 125757 10355 126053 10651
rect 126517 10355 126813 10651
rect 127277 10355 127573 10651
rect 128037 10355 128333 10651
rect 128797 10355 129093 10651
rect 129557 10355 129853 10651
rect 130317 10355 130613 10651
rect 131077 10355 131373 10651
rect 131837 10355 132133 10651
rect 132597 10355 132893 10651
rect 114357 9595 114653 9891
rect 115117 9595 115413 9891
rect 115877 9595 116173 9891
rect 116637 9595 116933 9891
rect 117397 9595 117693 9891
rect 118157 9595 118453 9891
rect 118917 9595 119213 9891
rect 119677 9595 119973 9891
rect 120437 9595 120733 9891
rect 121197 9595 121493 9891
rect 121957 9595 122253 9891
rect 122717 9595 123013 9891
rect 123477 9595 123773 9891
rect 124237 9595 124533 9891
rect 124997 9595 125293 9891
rect 125757 9595 126053 9891
rect 126517 9595 126813 9891
rect 127277 9595 127573 9891
rect 128037 9595 128333 9891
rect 128797 9595 129093 9891
rect 129557 9595 129853 9891
rect 130317 9595 130613 9891
rect 131077 9595 131373 9891
rect 131837 9595 132133 9891
rect 132597 9595 132893 9891
rect 114357 8835 114653 9131
rect 115117 8835 115413 9131
rect 115877 8835 116173 9131
rect 116637 8835 116933 9131
rect 117397 8835 117693 9131
rect 118157 8835 118453 9131
rect 118917 8835 119213 9131
rect 119677 8835 119973 9131
rect 120437 8835 120733 9131
rect 121197 8835 121493 9131
rect 121957 8835 122253 9131
rect 122717 8835 123013 9131
rect 123477 8835 123773 9131
rect 124237 8835 124533 9131
rect 124997 8835 125293 9131
rect 125757 8835 126053 9131
rect 126517 8835 126813 9131
rect 127277 8835 127573 9131
rect 128037 8835 128333 9131
rect 128797 8835 129093 9131
rect 129557 8835 129853 9131
rect 130317 8835 130613 9131
rect 131077 8835 131373 9131
rect 131837 8835 132133 9131
rect 132597 8835 132893 9131
rect 114357 8075 114653 8371
rect 115117 8075 115413 8371
rect 115877 8075 116173 8371
rect 116637 8075 116933 8371
rect 117397 8075 117693 8371
rect 118157 8075 118453 8371
rect 118917 8075 119213 8371
rect 119677 8075 119973 8371
rect 120437 8075 120733 8371
rect 121197 8075 121493 8371
rect 121957 8075 122253 8371
rect 122717 8075 123013 8371
rect 123477 8075 123773 8371
rect 124237 8075 124533 8371
rect 124997 8075 125293 8371
rect 125757 8075 126053 8371
rect 126517 8075 126813 8371
rect 127277 8075 127573 8371
rect 128037 8075 128333 8371
rect 128797 8075 129093 8371
rect 129557 8075 129853 8371
rect 130317 8075 130613 8371
rect 131077 8075 131373 8371
rect 131837 8075 132133 8371
rect 132597 8075 132893 8371
rect 114357 7315 114653 7611
rect 115117 7315 115413 7611
rect 115877 7315 116173 7611
rect 116637 7315 116933 7611
rect 117397 7315 117693 7611
rect 118157 7315 118453 7611
rect 118917 7315 119213 7611
rect 119677 7315 119973 7611
rect 120437 7315 120733 7611
rect 121197 7315 121493 7611
rect 121957 7315 122253 7611
rect 122717 7315 123013 7611
rect 123477 7315 123773 7611
rect 124237 7315 124533 7611
rect 124997 7315 125293 7611
rect 125757 7315 126053 7611
rect 126517 7315 126813 7611
rect 127277 7315 127573 7611
rect 128037 7315 128333 7611
rect 128797 7315 129093 7611
rect 129557 7315 129853 7611
rect 130317 7315 130613 7611
rect 131077 7315 131373 7611
rect 131837 7315 132133 7611
rect 132597 7315 132893 7611
rect 136157 30875 136453 31171
rect 136917 30875 137213 31171
rect 137677 30875 137973 31171
rect 138437 30875 138733 31171
rect 139197 30875 139493 31171
rect 139957 30875 140253 31171
rect 140717 30875 141013 31171
rect 141477 30875 141773 31171
rect 142237 30875 142533 31171
rect 142997 30875 143293 31171
rect 143757 30875 144053 31171
rect 144517 30875 144813 31171
rect 145277 30875 145573 31171
rect 146037 30875 146333 31171
rect 146797 30875 147093 31171
rect 147557 30875 147853 31171
rect 148317 30875 148613 31171
rect 149077 30875 149373 31171
rect 149837 30875 150133 31171
rect 150597 30875 150893 31171
rect 151357 30875 151653 31171
rect 152117 30875 152413 31171
rect 152877 30875 153173 31171
rect 153637 30875 153933 31171
rect 154397 30875 154693 31171
rect 136157 30115 136453 30411
rect 136917 30115 137213 30411
rect 137677 30115 137973 30411
rect 138437 30115 138733 30411
rect 139197 30115 139493 30411
rect 139957 30115 140253 30411
rect 140717 30115 141013 30411
rect 141477 30115 141773 30411
rect 142237 30115 142533 30411
rect 142997 30115 143293 30411
rect 143757 30115 144053 30411
rect 144517 30115 144813 30411
rect 145277 30115 145573 30411
rect 146037 30115 146333 30411
rect 146797 30115 147093 30411
rect 147557 30115 147853 30411
rect 148317 30115 148613 30411
rect 149077 30115 149373 30411
rect 149837 30115 150133 30411
rect 150597 30115 150893 30411
rect 151357 30115 151653 30411
rect 152117 30115 152413 30411
rect 152877 30115 153173 30411
rect 153637 30115 153933 30411
rect 154397 30115 154693 30411
rect 136157 29355 136453 29651
rect 136917 29355 137213 29651
rect 137677 29355 137973 29651
rect 138437 29355 138733 29651
rect 139197 29355 139493 29651
rect 139957 29355 140253 29651
rect 140717 29355 141013 29651
rect 141477 29355 141773 29651
rect 142237 29355 142533 29651
rect 142997 29355 143293 29651
rect 143757 29355 144053 29651
rect 144517 29355 144813 29651
rect 145277 29355 145573 29651
rect 146037 29355 146333 29651
rect 146797 29355 147093 29651
rect 147557 29355 147853 29651
rect 148317 29355 148613 29651
rect 149077 29355 149373 29651
rect 149837 29355 150133 29651
rect 150597 29355 150893 29651
rect 151357 29355 151653 29651
rect 152117 29355 152413 29651
rect 152877 29355 153173 29651
rect 153637 29355 153933 29651
rect 154397 29355 154693 29651
rect 136157 28595 136453 28891
rect 136917 28595 137213 28891
rect 137677 28595 137973 28891
rect 138437 28595 138733 28891
rect 139197 28595 139493 28891
rect 139957 28595 140253 28891
rect 140717 28595 141013 28891
rect 141477 28595 141773 28891
rect 142237 28595 142533 28891
rect 142997 28595 143293 28891
rect 143757 28595 144053 28891
rect 144517 28595 144813 28891
rect 145277 28595 145573 28891
rect 146037 28595 146333 28891
rect 146797 28595 147093 28891
rect 147557 28595 147853 28891
rect 148317 28595 148613 28891
rect 149077 28595 149373 28891
rect 149837 28595 150133 28891
rect 150597 28595 150893 28891
rect 151357 28595 151653 28891
rect 152117 28595 152413 28891
rect 152877 28595 153173 28891
rect 153637 28595 153933 28891
rect 154397 28595 154693 28891
rect 136157 27835 136453 28131
rect 136917 27835 137213 28131
rect 137677 27835 137973 28131
rect 138437 27835 138733 28131
rect 139197 27835 139493 28131
rect 139957 27835 140253 28131
rect 140717 27835 141013 28131
rect 141477 27835 141773 28131
rect 142237 27835 142533 28131
rect 142997 27835 143293 28131
rect 143757 27835 144053 28131
rect 144517 27835 144813 28131
rect 145277 27835 145573 28131
rect 146037 27835 146333 28131
rect 146797 27835 147093 28131
rect 147557 27835 147853 28131
rect 148317 27835 148613 28131
rect 149077 27835 149373 28131
rect 149837 27835 150133 28131
rect 150597 27835 150893 28131
rect 151357 27835 151653 28131
rect 152117 27835 152413 28131
rect 152877 27835 153173 28131
rect 153637 27835 153933 28131
rect 154397 27835 154693 28131
rect 136157 27075 136453 27371
rect 136917 27075 137213 27371
rect 137677 27075 137973 27371
rect 138437 27075 138733 27371
rect 139197 27075 139493 27371
rect 139957 27075 140253 27371
rect 140717 27075 141013 27371
rect 141477 27075 141773 27371
rect 142237 27075 142533 27371
rect 142997 27075 143293 27371
rect 143757 27075 144053 27371
rect 144517 27075 144813 27371
rect 145277 27075 145573 27371
rect 146037 27075 146333 27371
rect 146797 27075 147093 27371
rect 147557 27075 147853 27371
rect 148317 27075 148613 27371
rect 149077 27075 149373 27371
rect 149837 27075 150133 27371
rect 150597 27075 150893 27371
rect 151357 27075 151653 27371
rect 152117 27075 152413 27371
rect 152877 27075 153173 27371
rect 153637 27075 153933 27371
rect 154397 27075 154693 27371
rect 136157 26315 136453 26611
rect 136917 26315 137213 26611
rect 137677 26315 137973 26611
rect 138437 26315 138733 26611
rect 139197 26315 139493 26611
rect 139957 26315 140253 26611
rect 140717 26315 141013 26611
rect 141477 26315 141773 26611
rect 142237 26315 142533 26611
rect 142997 26315 143293 26611
rect 143757 26315 144053 26611
rect 144517 26315 144813 26611
rect 145277 26315 145573 26611
rect 146037 26315 146333 26611
rect 146797 26315 147093 26611
rect 147557 26315 147853 26611
rect 148317 26315 148613 26611
rect 149077 26315 149373 26611
rect 149837 26315 150133 26611
rect 150597 26315 150893 26611
rect 151357 26315 151653 26611
rect 152117 26315 152413 26611
rect 152877 26315 153173 26611
rect 153637 26315 153933 26611
rect 154397 26315 154693 26611
rect 136157 25555 136453 25851
rect 136917 25555 137213 25851
rect 137677 25555 137973 25851
rect 138437 25555 138733 25851
rect 139197 25555 139493 25851
rect 139957 25555 140253 25851
rect 140717 25555 141013 25851
rect 141477 25555 141773 25851
rect 142237 25555 142533 25851
rect 142997 25555 143293 25851
rect 143757 25555 144053 25851
rect 144517 25555 144813 25851
rect 145277 25555 145573 25851
rect 146037 25555 146333 25851
rect 146797 25555 147093 25851
rect 147557 25555 147853 25851
rect 148317 25555 148613 25851
rect 149077 25555 149373 25851
rect 149837 25555 150133 25851
rect 150597 25555 150893 25851
rect 151357 25555 151653 25851
rect 152117 25555 152413 25851
rect 152877 25555 153173 25851
rect 153637 25555 153933 25851
rect 154397 25555 154693 25851
rect 136157 24795 136453 25091
rect 136917 24795 137213 25091
rect 137677 24795 137973 25091
rect 138437 24795 138733 25091
rect 139197 24795 139493 25091
rect 139957 24795 140253 25091
rect 140717 24795 141013 25091
rect 141477 24795 141773 25091
rect 142237 24795 142533 25091
rect 142997 24795 143293 25091
rect 143757 24795 144053 25091
rect 144517 24795 144813 25091
rect 145277 24795 145573 25091
rect 146037 24795 146333 25091
rect 146797 24795 147093 25091
rect 147557 24795 147853 25091
rect 148317 24795 148613 25091
rect 149077 24795 149373 25091
rect 149837 24795 150133 25091
rect 150597 24795 150893 25091
rect 151357 24795 151653 25091
rect 152117 24795 152413 25091
rect 152877 24795 153173 25091
rect 153637 24795 153933 25091
rect 154397 24795 154693 25091
rect 136157 24035 136453 24331
rect 136917 24035 137213 24331
rect 137677 24035 137973 24331
rect 138437 24035 138733 24331
rect 139197 24035 139493 24331
rect 139957 24035 140253 24331
rect 140717 24035 141013 24331
rect 141477 24035 141773 24331
rect 142237 24035 142533 24331
rect 142997 24035 143293 24331
rect 143757 24035 144053 24331
rect 144517 24035 144813 24331
rect 145277 24035 145573 24331
rect 146037 24035 146333 24331
rect 146797 24035 147093 24331
rect 147557 24035 147853 24331
rect 148317 24035 148613 24331
rect 149077 24035 149373 24331
rect 149837 24035 150133 24331
rect 150597 24035 150893 24331
rect 151357 24035 151653 24331
rect 152117 24035 152413 24331
rect 152877 24035 153173 24331
rect 153637 24035 153933 24331
rect 154397 24035 154693 24331
rect 136157 23275 136453 23571
rect 136917 23275 137213 23571
rect 137677 23275 137973 23571
rect 138437 23275 138733 23571
rect 139197 23275 139493 23571
rect 139957 23275 140253 23571
rect 140717 23275 141013 23571
rect 141477 23275 141773 23571
rect 142237 23275 142533 23571
rect 142997 23275 143293 23571
rect 143757 23275 144053 23571
rect 144517 23275 144813 23571
rect 145277 23275 145573 23571
rect 146037 23275 146333 23571
rect 146797 23275 147093 23571
rect 147557 23275 147853 23571
rect 148317 23275 148613 23571
rect 149077 23275 149373 23571
rect 149837 23275 150133 23571
rect 150597 23275 150893 23571
rect 151357 23275 151653 23571
rect 152117 23275 152413 23571
rect 152877 23275 153173 23571
rect 153637 23275 153933 23571
rect 154397 23275 154693 23571
rect 136157 22515 136453 22811
rect 136917 22515 137213 22811
rect 137677 22515 137973 22811
rect 138437 22515 138733 22811
rect 139197 22515 139493 22811
rect 139957 22515 140253 22811
rect 140717 22515 141013 22811
rect 141477 22515 141773 22811
rect 142237 22515 142533 22811
rect 142997 22515 143293 22811
rect 143757 22515 144053 22811
rect 144517 22515 144813 22811
rect 145277 22515 145573 22811
rect 146037 22515 146333 22811
rect 146797 22515 147093 22811
rect 147557 22515 147853 22811
rect 148317 22515 148613 22811
rect 149077 22515 149373 22811
rect 149837 22515 150133 22811
rect 150597 22515 150893 22811
rect 151357 22515 151653 22811
rect 152117 22515 152413 22811
rect 152877 22515 153173 22811
rect 153637 22515 153933 22811
rect 154397 22515 154693 22811
rect 136157 21755 136453 22051
rect 136917 21755 137213 22051
rect 137677 21755 137973 22051
rect 138437 21755 138733 22051
rect 139197 21755 139493 22051
rect 139957 21755 140253 22051
rect 140717 21755 141013 22051
rect 141477 21755 141773 22051
rect 142237 21755 142533 22051
rect 142997 21755 143293 22051
rect 143757 21755 144053 22051
rect 144517 21755 144813 22051
rect 145277 21755 145573 22051
rect 146037 21755 146333 22051
rect 146797 21755 147093 22051
rect 147557 21755 147853 22051
rect 148317 21755 148613 22051
rect 149077 21755 149373 22051
rect 149837 21755 150133 22051
rect 150597 21755 150893 22051
rect 151357 21755 151653 22051
rect 152117 21755 152413 22051
rect 152877 21755 153173 22051
rect 153637 21755 153933 22051
rect 154397 21755 154693 22051
rect 136157 20995 136453 21291
rect 136917 20995 137213 21291
rect 137677 20995 137973 21291
rect 138437 20995 138733 21291
rect 139197 20995 139493 21291
rect 139957 20995 140253 21291
rect 140717 20995 141013 21291
rect 141477 20995 141773 21291
rect 142237 20995 142533 21291
rect 142997 20995 143293 21291
rect 143757 20995 144053 21291
rect 144517 20995 144813 21291
rect 145277 20995 145573 21291
rect 146037 20995 146333 21291
rect 146797 20995 147093 21291
rect 147557 20995 147853 21291
rect 148317 20995 148613 21291
rect 149077 20995 149373 21291
rect 149837 20995 150133 21291
rect 150597 20995 150893 21291
rect 151357 20995 151653 21291
rect 152117 20995 152413 21291
rect 152877 20995 153173 21291
rect 153637 20995 153933 21291
rect 154397 20995 154693 21291
rect 136157 20235 136453 20531
rect 136917 20235 137213 20531
rect 137677 20235 137973 20531
rect 138437 20235 138733 20531
rect 139197 20235 139493 20531
rect 139957 20235 140253 20531
rect 140717 20235 141013 20531
rect 141477 20235 141773 20531
rect 142237 20235 142533 20531
rect 142997 20235 143293 20531
rect 143757 20235 144053 20531
rect 144517 20235 144813 20531
rect 145277 20235 145573 20531
rect 146037 20235 146333 20531
rect 146797 20235 147093 20531
rect 147557 20235 147853 20531
rect 148317 20235 148613 20531
rect 149077 20235 149373 20531
rect 149837 20235 150133 20531
rect 150597 20235 150893 20531
rect 151357 20235 151653 20531
rect 152117 20235 152413 20531
rect 152877 20235 153173 20531
rect 153637 20235 153933 20531
rect 154397 20235 154693 20531
rect 136157 19475 136453 19771
rect 136917 19475 137213 19771
rect 137677 19475 137973 19771
rect 138437 19475 138733 19771
rect 139197 19475 139493 19771
rect 139957 19475 140253 19771
rect 140717 19475 141013 19771
rect 141477 19475 141773 19771
rect 142237 19475 142533 19771
rect 142997 19475 143293 19771
rect 143757 19475 144053 19771
rect 144517 19475 144813 19771
rect 145277 19475 145573 19771
rect 146037 19475 146333 19771
rect 146797 19475 147093 19771
rect 147557 19475 147853 19771
rect 148317 19475 148613 19771
rect 149077 19475 149373 19771
rect 149837 19475 150133 19771
rect 150597 19475 150893 19771
rect 151357 19475 151653 19771
rect 152117 19475 152413 19771
rect 152877 19475 153173 19771
rect 153637 19475 153933 19771
rect 154397 19475 154693 19771
rect 136157 18715 136453 19011
rect 136917 18715 137213 19011
rect 137677 18715 137973 19011
rect 138437 18715 138733 19011
rect 139197 18715 139493 19011
rect 139957 18715 140253 19011
rect 140717 18715 141013 19011
rect 141477 18715 141773 19011
rect 142237 18715 142533 19011
rect 142997 18715 143293 19011
rect 143757 18715 144053 19011
rect 144517 18715 144813 19011
rect 145277 18715 145573 19011
rect 146037 18715 146333 19011
rect 146797 18715 147093 19011
rect 147557 18715 147853 19011
rect 148317 18715 148613 19011
rect 149077 18715 149373 19011
rect 149837 18715 150133 19011
rect 150597 18715 150893 19011
rect 151357 18715 151653 19011
rect 152117 18715 152413 19011
rect 152877 18715 153173 19011
rect 153637 18715 153933 19011
rect 154397 18715 154693 19011
rect 136157 17955 136453 18251
rect 136917 17955 137213 18251
rect 137677 17955 137973 18251
rect 138437 17955 138733 18251
rect 139197 17955 139493 18251
rect 139957 17955 140253 18251
rect 140717 17955 141013 18251
rect 141477 17955 141773 18251
rect 142237 17955 142533 18251
rect 142997 17955 143293 18251
rect 143757 17955 144053 18251
rect 144517 17955 144813 18251
rect 145277 17955 145573 18251
rect 146037 17955 146333 18251
rect 146797 17955 147093 18251
rect 147557 17955 147853 18251
rect 148317 17955 148613 18251
rect 149077 17955 149373 18251
rect 149837 17955 150133 18251
rect 150597 17955 150893 18251
rect 151357 17955 151653 18251
rect 152117 17955 152413 18251
rect 152877 17955 153173 18251
rect 153637 17955 153933 18251
rect 154397 17955 154693 18251
rect 136157 17195 136453 17491
rect 136917 17195 137213 17491
rect 137677 17195 137973 17491
rect 138437 17195 138733 17491
rect 139197 17195 139493 17491
rect 139957 17195 140253 17491
rect 140717 17195 141013 17491
rect 141477 17195 141773 17491
rect 142237 17195 142533 17491
rect 142997 17195 143293 17491
rect 143757 17195 144053 17491
rect 144517 17195 144813 17491
rect 145277 17195 145573 17491
rect 146037 17195 146333 17491
rect 146797 17195 147093 17491
rect 147557 17195 147853 17491
rect 148317 17195 148613 17491
rect 149077 17195 149373 17491
rect 149837 17195 150133 17491
rect 150597 17195 150893 17491
rect 151357 17195 151653 17491
rect 152117 17195 152413 17491
rect 152877 17195 153173 17491
rect 153637 17195 153933 17491
rect 154397 17195 154693 17491
rect 136157 16435 136453 16731
rect 136917 16435 137213 16731
rect 137677 16435 137973 16731
rect 138437 16435 138733 16731
rect 139197 16435 139493 16731
rect 139957 16435 140253 16731
rect 140717 16435 141013 16731
rect 141477 16435 141773 16731
rect 142237 16435 142533 16731
rect 142997 16435 143293 16731
rect 143757 16435 144053 16731
rect 144517 16435 144813 16731
rect 145277 16435 145573 16731
rect 146037 16435 146333 16731
rect 146797 16435 147093 16731
rect 147557 16435 147853 16731
rect 148317 16435 148613 16731
rect 149077 16435 149373 16731
rect 149837 16435 150133 16731
rect 150597 16435 150893 16731
rect 151357 16435 151653 16731
rect 152117 16435 152413 16731
rect 152877 16435 153173 16731
rect 153637 16435 153933 16731
rect 154397 16435 154693 16731
rect 136157 15675 136453 15971
rect 136917 15675 137213 15971
rect 137677 15675 137973 15971
rect 138437 15675 138733 15971
rect 139197 15675 139493 15971
rect 139957 15675 140253 15971
rect 140717 15675 141013 15971
rect 141477 15675 141773 15971
rect 142237 15675 142533 15971
rect 142997 15675 143293 15971
rect 143757 15675 144053 15971
rect 144517 15675 144813 15971
rect 145277 15675 145573 15971
rect 146037 15675 146333 15971
rect 146797 15675 147093 15971
rect 147557 15675 147853 15971
rect 148317 15675 148613 15971
rect 149077 15675 149373 15971
rect 149837 15675 150133 15971
rect 150597 15675 150893 15971
rect 151357 15675 151653 15971
rect 152117 15675 152413 15971
rect 152877 15675 153173 15971
rect 153637 15675 153933 15971
rect 154397 15675 154693 15971
rect 136157 14915 136453 15211
rect 136917 14915 137213 15211
rect 137677 14915 137973 15211
rect 138437 14915 138733 15211
rect 139197 14915 139493 15211
rect 139957 14915 140253 15211
rect 140717 14915 141013 15211
rect 141477 14915 141773 15211
rect 142237 14915 142533 15211
rect 142997 14915 143293 15211
rect 143757 14915 144053 15211
rect 144517 14915 144813 15211
rect 145277 14915 145573 15211
rect 146037 14915 146333 15211
rect 146797 14915 147093 15211
rect 147557 14915 147853 15211
rect 148317 14915 148613 15211
rect 149077 14915 149373 15211
rect 149837 14915 150133 15211
rect 150597 14915 150893 15211
rect 151357 14915 151653 15211
rect 152117 14915 152413 15211
rect 152877 14915 153173 15211
rect 153637 14915 153933 15211
rect 154397 14915 154693 15211
rect 136157 14155 136453 14451
rect 136917 14155 137213 14451
rect 137677 14155 137973 14451
rect 138437 14155 138733 14451
rect 139197 14155 139493 14451
rect 139957 14155 140253 14451
rect 140717 14155 141013 14451
rect 141477 14155 141773 14451
rect 142237 14155 142533 14451
rect 142997 14155 143293 14451
rect 143757 14155 144053 14451
rect 144517 14155 144813 14451
rect 145277 14155 145573 14451
rect 146037 14155 146333 14451
rect 146797 14155 147093 14451
rect 147557 14155 147853 14451
rect 148317 14155 148613 14451
rect 149077 14155 149373 14451
rect 149837 14155 150133 14451
rect 150597 14155 150893 14451
rect 151357 14155 151653 14451
rect 152117 14155 152413 14451
rect 152877 14155 153173 14451
rect 153637 14155 153933 14451
rect 154397 14155 154693 14451
rect 136157 13395 136453 13691
rect 136917 13395 137213 13691
rect 137677 13395 137973 13691
rect 138437 13395 138733 13691
rect 139197 13395 139493 13691
rect 139957 13395 140253 13691
rect 140717 13395 141013 13691
rect 141477 13395 141773 13691
rect 142237 13395 142533 13691
rect 142997 13395 143293 13691
rect 143757 13395 144053 13691
rect 144517 13395 144813 13691
rect 145277 13395 145573 13691
rect 146037 13395 146333 13691
rect 146797 13395 147093 13691
rect 147557 13395 147853 13691
rect 148317 13395 148613 13691
rect 149077 13395 149373 13691
rect 149837 13395 150133 13691
rect 150597 13395 150893 13691
rect 151357 13395 151653 13691
rect 152117 13395 152413 13691
rect 152877 13395 153173 13691
rect 153637 13395 153933 13691
rect 154397 13395 154693 13691
rect 136157 12635 136453 12931
rect 136917 12635 137213 12931
rect 137677 12635 137973 12931
rect 138437 12635 138733 12931
rect 139197 12635 139493 12931
rect 139957 12635 140253 12931
rect 140717 12635 141013 12931
rect 141477 12635 141773 12931
rect 142237 12635 142533 12931
rect 142997 12635 143293 12931
rect 143757 12635 144053 12931
rect 144517 12635 144813 12931
rect 145277 12635 145573 12931
rect 146037 12635 146333 12931
rect 146797 12635 147093 12931
rect 147557 12635 147853 12931
rect 148317 12635 148613 12931
rect 149077 12635 149373 12931
rect 149837 12635 150133 12931
rect 150597 12635 150893 12931
rect 151357 12635 151653 12931
rect 152117 12635 152413 12931
rect 152877 12635 153173 12931
rect 153637 12635 153933 12931
rect 154397 12635 154693 12931
rect 136157 11875 136453 12171
rect 136917 11875 137213 12171
rect 137677 11875 137973 12171
rect 138437 11875 138733 12171
rect 139197 11875 139493 12171
rect 139957 11875 140253 12171
rect 140717 11875 141013 12171
rect 141477 11875 141773 12171
rect 142237 11875 142533 12171
rect 142997 11875 143293 12171
rect 143757 11875 144053 12171
rect 144517 11875 144813 12171
rect 145277 11875 145573 12171
rect 146037 11875 146333 12171
rect 146797 11875 147093 12171
rect 147557 11875 147853 12171
rect 148317 11875 148613 12171
rect 149077 11875 149373 12171
rect 149837 11875 150133 12171
rect 150597 11875 150893 12171
rect 151357 11875 151653 12171
rect 152117 11875 152413 12171
rect 152877 11875 153173 12171
rect 153637 11875 153933 12171
rect 154397 11875 154693 12171
rect 136157 11115 136453 11411
rect 136917 11115 137213 11411
rect 137677 11115 137973 11411
rect 138437 11115 138733 11411
rect 139197 11115 139493 11411
rect 139957 11115 140253 11411
rect 140717 11115 141013 11411
rect 141477 11115 141773 11411
rect 142237 11115 142533 11411
rect 142997 11115 143293 11411
rect 143757 11115 144053 11411
rect 144517 11115 144813 11411
rect 145277 11115 145573 11411
rect 146037 11115 146333 11411
rect 146797 11115 147093 11411
rect 147557 11115 147853 11411
rect 148317 11115 148613 11411
rect 149077 11115 149373 11411
rect 149837 11115 150133 11411
rect 150597 11115 150893 11411
rect 151357 11115 151653 11411
rect 152117 11115 152413 11411
rect 152877 11115 153173 11411
rect 153637 11115 153933 11411
rect 154397 11115 154693 11411
rect 136157 10355 136453 10651
rect 136917 10355 137213 10651
rect 137677 10355 137973 10651
rect 138437 10355 138733 10651
rect 139197 10355 139493 10651
rect 139957 10355 140253 10651
rect 140717 10355 141013 10651
rect 141477 10355 141773 10651
rect 142237 10355 142533 10651
rect 142997 10355 143293 10651
rect 143757 10355 144053 10651
rect 144517 10355 144813 10651
rect 145277 10355 145573 10651
rect 146037 10355 146333 10651
rect 146797 10355 147093 10651
rect 147557 10355 147853 10651
rect 148317 10355 148613 10651
rect 149077 10355 149373 10651
rect 149837 10355 150133 10651
rect 150597 10355 150893 10651
rect 151357 10355 151653 10651
rect 152117 10355 152413 10651
rect 152877 10355 153173 10651
rect 153637 10355 153933 10651
rect 154397 10355 154693 10651
rect 136157 9595 136453 9891
rect 136917 9595 137213 9891
rect 137677 9595 137973 9891
rect 138437 9595 138733 9891
rect 139197 9595 139493 9891
rect 139957 9595 140253 9891
rect 140717 9595 141013 9891
rect 141477 9595 141773 9891
rect 142237 9595 142533 9891
rect 142997 9595 143293 9891
rect 143757 9595 144053 9891
rect 144517 9595 144813 9891
rect 145277 9595 145573 9891
rect 146037 9595 146333 9891
rect 146797 9595 147093 9891
rect 147557 9595 147853 9891
rect 148317 9595 148613 9891
rect 149077 9595 149373 9891
rect 149837 9595 150133 9891
rect 150597 9595 150893 9891
rect 151357 9595 151653 9891
rect 152117 9595 152413 9891
rect 152877 9595 153173 9891
rect 153637 9595 153933 9891
rect 154397 9595 154693 9891
rect 136157 8835 136453 9131
rect 136917 8835 137213 9131
rect 137677 8835 137973 9131
rect 138437 8835 138733 9131
rect 139197 8835 139493 9131
rect 139957 8835 140253 9131
rect 140717 8835 141013 9131
rect 141477 8835 141773 9131
rect 142237 8835 142533 9131
rect 142997 8835 143293 9131
rect 143757 8835 144053 9131
rect 144517 8835 144813 9131
rect 145277 8835 145573 9131
rect 146037 8835 146333 9131
rect 146797 8835 147093 9131
rect 147557 8835 147853 9131
rect 148317 8835 148613 9131
rect 149077 8835 149373 9131
rect 149837 8835 150133 9131
rect 150597 8835 150893 9131
rect 151357 8835 151653 9131
rect 152117 8835 152413 9131
rect 152877 8835 153173 9131
rect 153637 8835 153933 9131
rect 154397 8835 154693 9131
rect 136157 8075 136453 8371
rect 136917 8075 137213 8371
rect 137677 8075 137973 8371
rect 138437 8075 138733 8371
rect 139197 8075 139493 8371
rect 139957 8075 140253 8371
rect 140717 8075 141013 8371
rect 141477 8075 141773 8371
rect 142237 8075 142533 8371
rect 142997 8075 143293 8371
rect 143757 8075 144053 8371
rect 144517 8075 144813 8371
rect 145277 8075 145573 8371
rect 146037 8075 146333 8371
rect 146797 8075 147093 8371
rect 147557 8075 147853 8371
rect 148317 8075 148613 8371
rect 149077 8075 149373 8371
rect 149837 8075 150133 8371
rect 150597 8075 150893 8371
rect 151357 8075 151653 8371
rect 152117 8075 152413 8371
rect 152877 8075 153173 8371
rect 153637 8075 153933 8371
rect 154397 8075 154693 8371
rect 136157 7315 136453 7611
rect 136917 7315 137213 7611
rect 137677 7315 137973 7611
rect 138437 7315 138733 7611
rect 139197 7315 139493 7611
rect 139957 7315 140253 7611
rect 140717 7315 141013 7611
rect 141477 7315 141773 7611
rect 142237 7315 142533 7611
rect 142997 7315 143293 7611
rect 143757 7315 144053 7611
rect 144517 7315 144813 7611
rect 145277 7315 145573 7611
rect 146037 7315 146333 7611
rect 146797 7315 147093 7611
rect 147557 7315 147853 7611
rect 148317 7315 148613 7611
rect 149077 7315 149373 7611
rect 149837 7315 150133 7611
rect 150597 7315 150893 7611
rect 151357 7315 151653 7611
rect 152117 7315 152413 7611
rect 152877 7315 153173 7611
rect 153637 7315 153933 7611
rect 154397 7315 154693 7611
rect 157957 30875 158253 31171
rect 158717 30875 159013 31171
rect 159477 30875 159773 31171
rect 160237 30875 160533 31171
rect 160997 30875 161293 31171
rect 161757 30875 162053 31171
rect 162517 30875 162813 31171
rect 163277 30875 163573 31171
rect 164037 30875 164333 31171
rect 164797 30875 165093 31171
rect 165557 30875 165853 31171
rect 166317 30875 166613 31171
rect 167077 30875 167373 31171
rect 167837 30875 168133 31171
rect 168597 30875 168893 31171
rect 169357 30875 169653 31171
rect 170117 30875 170413 31171
rect 170877 30875 171173 31171
rect 171637 30875 171933 31171
rect 172397 30875 172693 31171
rect 173157 30875 173453 31171
rect 173917 30875 174213 31171
rect 174677 30875 174973 31171
rect 175437 30875 175733 31171
rect 176197 30875 176493 31171
rect 157957 30115 158253 30411
rect 158717 30115 159013 30411
rect 159477 30115 159773 30411
rect 160237 30115 160533 30411
rect 160997 30115 161293 30411
rect 161757 30115 162053 30411
rect 162517 30115 162813 30411
rect 163277 30115 163573 30411
rect 164037 30115 164333 30411
rect 164797 30115 165093 30411
rect 165557 30115 165853 30411
rect 166317 30115 166613 30411
rect 167077 30115 167373 30411
rect 167837 30115 168133 30411
rect 168597 30115 168893 30411
rect 169357 30115 169653 30411
rect 170117 30115 170413 30411
rect 170877 30115 171173 30411
rect 171637 30115 171933 30411
rect 172397 30115 172693 30411
rect 173157 30115 173453 30411
rect 173917 30115 174213 30411
rect 174677 30115 174973 30411
rect 175437 30115 175733 30411
rect 176197 30115 176493 30411
rect 157957 29355 158253 29651
rect 158717 29355 159013 29651
rect 159477 29355 159773 29651
rect 160237 29355 160533 29651
rect 160997 29355 161293 29651
rect 161757 29355 162053 29651
rect 162517 29355 162813 29651
rect 163277 29355 163573 29651
rect 164037 29355 164333 29651
rect 164797 29355 165093 29651
rect 165557 29355 165853 29651
rect 166317 29355 166613 29651
rect 167077 29355 167373 29651
rect 167837 29355 168133 29651
rect 168597 29355 168893 29651
rect 169357 29355 169653 29651
rect 170117 29355 170413 29651
rect 170877 29355 171173 29651
rect 171637 29355 171933 29651
rect 172397 29355 172693 29651
rect 173157 29355 173453 29651
rect 173917 29355 174213 29651
rect 174677 29355 174973 29651
rect 175437 29355 175733 29651
rect 176197 29355 176493 29651
rect 157957 28595 158253 28891
rect 158717 28595 159013 28891
rect 159477 28595 159773 28891
rect 160237 28595 160533 28891
rect 160997 28595 161293 28891
rect 161757 28595 162053 28891
rect 162517 28595 162813 28891
rect 163277 28595 163573 28891
rect 164037 28595 164333 28891
rect 164797 28595 165093 28891
rect 165557 28595 165853 28891
rect 166317 28595 166613 28891
rect 167077 28595 167373 28891
rect 167837 28595 168133 28891
rect 168597 28595 168893 28891
rect 169357 28595 169653 28891
rect 170117 28595 170413 28891
rect 170877 28595 171173 28891
rect 171637 28595 171933 28891
rect 172397 28595 172693 28891
rect 173157 28595 173453 28891
rect 173917 28595 174213 28891
rect 174677 28595 174973 28891
rect 175437 28595 175733 28891
rect 176197 28595 176493 28891
rect 157957 27835 158253 28131
rect 158717 27835 159013 28131
rect 159477 27835 159773 28131
rect 160237 27835 160533 28131
rect 160997 27835 161293 28131
rect 161757 27835 162053 28131
rect 162517 27835 162813 28131
rect 163277 27835 163573 28131
rect 164037 27835 164333 28131
rect 164797 27835 165093 28131
rect 165557 27835 165853 28131
rect 166317 27835 166613 28131
rect 167077 27835 167373 28131
rect 167837 27835 168133 28131
rect 168597 27835 168893 28131
rect 169357 27835 169653 28131
rect 170117 27835 170413 28131
rect 170877 27835 171173 28131
rect 171637 27835 171933 28131
rect 172397 27835 172693 28131
rect 173157 27835 173453 28131
rect 173917 27835 174213 28131
rect 174677 27835 174973 28131
rect 175437 27835 175733 28131
rect 176197 27835 176493 28131
rect 157957 27075 158253 27371
rect 158717 27075 159013 27371
rect 159477 27075 159773 27371
rect 160237 27075 160533 27371
rect 160997 27075 161293 27371
rect 161757 27075 162053 27371
rect 162517 27075 162813 27371
rect 163277 27075 163573 27371
rect 164037 27075 164333 27371
rect 164797 27075 165093 27371
rect 165557 27075 165853 27371
rect 166317 27075 166613 27371
rect 167077 27075 167373 27371
rect 167837 27075 168133 27371
rect 168597 27075 168893 27371
rect 169357 27075 169653 27371
rect 170117 27075 170413 27371
rect 170877 27075 171173 27371
rect 171637 27075 171933 27371
rect 172397 27075 172693 27371
rect 173157 27075 173453 27371
rect 173917 27075 174213 27371
rect 174677 27075 174973 27371
rect 175437 27075 175733 27371
rect 176197 27075 176493 27371
rect 157957 26315 158253 26611
rect 158717 26315 159013 26611
rect 159477 26315 159773 26611
rect 160237 26315 160533 26611
rect 160997 26315 161293 26611
rect 161757 26315 162053 26611
rect 162517 26315 162813 26611
rect 163277 26315 163573 26611
rect 164037 26315 164333 26611
rect 164797 26315 165093 26611
rect 165557 26315 165853 26611
rect 166317 26315 166613 26611
rect 167077 26315 167373 26611
rect 167837 26315 168133 26611
rect 168597 26315 168893 26611
rect 169357 26315 169653 26611
rect 170117 26315 170413 26611
rect 170877 26315 171173 26611
rect 171637 26315 171933 26611
rect 172397 26315 172693 26611
rect 173157 26315 173453 26611
rect 173917 26315 174213 26611
rect 174677 26315 174973 26611
rect 175437 26315 175733 26611
rect 176197 26315 176493 26611
rect 157957 25555 158253 25851
rect 158717 25555 159013 25851
rect 159477 25555 159773 25851
rect 160237 25555 160533 25851
rect 160997 25555 161293 25851
rect 161757 25555 162053 25851
rect 162517 25555 162813 25851
rect 163277 25555 163573 25851
rect 164037 25555 164333 25851
rect 164797 25555 165093 25851
rect 165557 25555 165853 25851
rect 166317 25555 166613 25851
rect 167077 25555 167373 25851
rect 167837 25555 168133 25851
rect 168597 25555 168893 25851
rect 169357 25555 169653 25851
rect 170117 25555 170413 25851
rect 170877 25555 171173 25851
rect 171637 25555 171933 25851
rect 172397 25555 172693 25851
rect 173157 25555 173453 25851
rect 173917 25555 174213 25851
rect 174677 25555 174973 25851
rect 175437 25555 175733 25851
rect 176197 25555 176493 25851
rect 157957 24795 158253 25091
rect 158717 24795 159013 25091
rect 159477 24795 159773 25091
rect 160237 24795 160533 25091
rect 160997 24795 161293 25091
rect 161757 24795 162053 25091
rect 162517 24795 162813 25091
rect 163277 24795 163573 25091
rect 164037 24795 164333 25091
rect 164797 24795 165093 25091
rect 165557 24795 165853 25091
rect 166317 24795 166613 25091
rect 167077 24795 167373 25091
rect 167837 24795 168133 25091
rect 168597 24795 168893 25091
rect 169357 24795 169653 25091
rect 170117 24795 170413 25091
rect 170877 24795 171173 25091
rect 171637 24795 171933 25091
rect 172397 24795 172693 25091
rect 173157 24795 173453 25091
rect 173917 24795 174213 25091
rect 174677 24795 174973 25091
rect 175437 24795 175733 25091
rect 176197 24795 176493 25091
rect 157957 24035 158253 24331
rect 158717 24035 159013 24331
rect 159477 24035 159773 24331
rect 160237 24035 160533 24331
rect 160997 24035 161293 24331
rect 161757 24035 162053 24331
rect 162517 24035 162813 24331
rect 163277 24035 163573 24331
rect 164037 24035 164333 24331
rect 164797 24035 165093 24331
rect 165557 24035 165853 24331
rect 166317 24035 166613 24331
rect 167077 24035 167373 24331
rect 167837 24035 168133 24331
rect 168597 24035 168893 24331
rect 169357 24035 169653 24331
rect 170117 24035 170413 24331
rect 170877 24035 171173 24331
rect 171637 24035 171933 24331
rect 172397 24035 172693 24331
rect 173157 24035 173453 24331
rect 173917 24035 174213 24331
rect 174677 24035 174973 24331
rect 175437 24035 175733 24331
rect 176197 24035 176493 24331
rect 157957 23275 158253 23571
rect 158717 23275 159013 23571
rect 159477 23275 159773 23571
rect 160237 23275 160533 23571
rect 160997 23275 161293 23571
rect 161757 23275 162053 23571
rect 162517 23275 162813 23571
rect 163277 23275 163573 23571
rect 164037 23275 164333 23571
rect 164797 23275 165093 23571
rect 165557 23275 165853 23571
rect 166317 23275 166613 23571
rect 167077 23275 167373 23571
rect 167837 23275 168133 23571
rect 168597 23275 168893 23571
rect 169357 23275 169653 23571
rect 170117 23275 170413 23571
rect 170877 23275 171173 23571
rect 171637 23275 171933 23571
rect 172397 23275 172693 23571
rect 173157 23275 173453 23571
rect 173917 23275 174213 23571
rect 174677 23275 174973 23571
rect 175437 23275 175733 23571
rect 176197 23275 176493 23571
rect 157957 22515 158253 22811
rect 158717 22515 159013 22811
rect 159477 22515 159773 22811
rect 160237 22515 160533 22811
rect 160997 22515 161293 22811
rect 161757 22515 162053 22811
rect 162517 22515 162813 22811
rect 163277 22515 163573 22811
rect 164037 22515 164333 22811
rect 164797 22515 165093 22811
rect 165557 22515 165853 22811
rect 166317 22515 166613 22811
rect 167077 22515 167373 22811
rect 167837 22515 168133 22811
rect 168597 22515 168893 22811
rect 169357 22515 169653 22811
rect 170117 22515 170413 22811
rect 170877 22515 171173 22811
rect 171637 22515 171933 22811
rect 172397 22515 172693 22811
rect 173157 22515 173453 22811
rect 173917 22515 174213 22811
rect 174677 22515 174973 22811
rect 175437 22515 175733 22811
rect 176197 22515 176493 22811
rect 157957 21755 158253 22051
rect 158717 21755 159013 22051
rect 159477 21755 159773 22051
rect 160237 21755 160533 22051
rect 160997 21755 161293 22051
rect 161757 21755 162053 22051
rect 162517 21755 162813 22051
rect 163277 21755 163573 22051
rect 164037 21755 164333 22051
rect 164797 21755 165093 22051
rect 165557 21755 165853 22051
rect 166317 21755 166613 22051
rect 167077 21755 167373 22051
rect 167837 21755 168133 22051
rect 168597 21755 168893 22051
rect 169357 21755 169653 22051
rect 170117 21755 170413 22051
rect 170877 21755 171173 22051
rect 171637 21755 171933 22051
rect 172397 21755 172693 22051
rect 173157 21755 173453 22051
rect 173917 21755 174213 22051
rect 174677 21755 174973 22051
rect 175437 21755 175733 22051
rect 176197 21755 176493 22051
rect 157957 20995 158253 21291
rect 158717 20995 159013 21291
rect 159477 20995 159773 21291
rect 160237 20995 160533 21291
rect 160997 20995 161293 21291
rect 161757 20995 162053 21291
rect 162517 20995 162813 21291
rect 163277 20995 163573 21291
rect 164037 20995 164333 21291
rect 164797 20995 165093 21291
rect 165557 20995 165853 21291
rect 166317 20995 166613 21291
rect 167077 20995 167373 21291
rect 167837 20995 168133 21291
rect 168597 20995 168893 21291
rect 169357 20995 169653 21291
rect 170117 20995 170413 21291
rect 170877 20995 171173 21291
rect 171637 20995 171933 21291
rect 172397 20995 172693 21291
rect 173157 20995 173453 21291
rect 173917 20995 174213 21291
rect 174677 20995 174973 21291
rect 175437 20995 175733 21291
rect 176197 20995 176493 21291
rect 157957 20235 158253 20531
rect 158717 20235 159013 20531
rect 159477 20235 159773 20531
rect 160237 20235 160533 20531
rect 160997 20235 161293 20531
rect 161757 20235 162053 20531
rect 162517 20235 162813 20531
rect 163277 20235 163573 20531
rect 164037 20235 164333 20531
rect 164797 20235 165093 20531
rect 165557 20235 165853 20531
rect 166317 20235 166613 20531
rect 167077 20235 167373 20531
rect 167837 20235 168133 20531
rect 168597 20235 168893 20531
rect 169357 20235 169653 20531
rect 170117 20235 170413 20531
rect 170877 20235 171173 20531
rect 171637 20235 171933 20531
rect 172397 20235 172693 20531
rect 173157 20235 173453 20531
rect 173917 20235 174213 20531
rect 174677 20235 174973 20531
rect 175437 20235 175733 20531
rect 176197 20235 176493 20531
rect 157957 19475 158253 19771
rect 158717 19475 159013 19771
rect 159477 19475 159773 19771
rect 160237 19475 160533 19771
rect 160997 19475 161293 19771
rect 161757 19475 162053 19771
rect 162517 19475 162813 19771
rect 163277 19475 163573 19771
rect 164037 19475 164333 19771
rect 164797 19475 165093 19771
rect 165557 19475 165853 19771
rect 166317 19475 166613 19771
rect 167077 19475 167373 19771
rect 167837 19475 168133 19771
rect 168597 19475 168893 19771
rect 169357 19475 169653 19771
rect 170117 19475 170413 19771
rect 170877 19475 171173 19771
rect 171637 19475 171933 19771
rect 172397 19475 172693 19771
rect 173157 19475 173453 19771
rect 173917 19475 174213 19771
rect 174677 19475 174973 19771
rect 175437 19475 175733 19771
rect 176197 19475 176493 19771
rect 157957 18715 158253 19011
rect 158717 18715 159013 19011
rect 159477 18715 159773 19011
rect 160237 18715 160533 19011
rect 160997 18715 161293 19011
rect 161757 18715 162053 19011
rect 162517 18715 162813 19011
rect 163277 18715 163573 19011
rect 164037 18715 164333 19011
rect 164797 18715 165093 19011
rect 165557 18715 165853 19011
rect 166317 18715 166613 19011
rect 167077 18715 167373 19011
rect 167837 18715 168133 19011
rect 168597 18715 168893 19011
rect 169357 18715 169653 19011
rect 170117 18715 170413 19011
rect 170877 18715 171173 19011
rect 171637 18715 171933 19011
rect 172397 18715 172693 19011
rect 173157 18715 173453 19011
rect 173917 18715 174213 19011
rect 174677 18715 174973 19011
rect 175437 18715 175733 19011
rect 176197 18715 176493 19011
rect 157957 17955 158253 18251
rect 158717 17955 159013 18251
rect 159477 17955 159773 18251
rect 160237 17955 160533 18251
rect 160997 17955 161293 18251
rect 161757 17955 162053 18251
rect 162517 17955 162813 18251
rect 163277 17955 163573 18251
rect 164037 17955 164333 18251
rect 164797 17955 165093 18251
rect 165557 17955 165853 18251
rect 166317 17955 166613 18251
rect 167077 17955 167373 18251
rect 167837 17955 168133 18251
rect 168597 17955 168893 18251
rect 169357 17955 169653 18251
rect 170117 17955 170413 18251
rect 170877 17955 171173 18251
rect 171637 17955 171933 18251
rect 172397 17955 172693 18251
rect 173157 17955 173453 18251
rect 173917 17955 174213 18251
rect 174677 17955 174973 18251
rect 175437 17955 175733 18251
rect 176197 17955 176493 18251
rect 157957 17195 158253 17491
rect 158717 17195 159013 17491
rect 159477 17195 159773 17491
rect 160237 17195 160533 17491
rect 160997 17195 161293 17491
rect 161757 17195 162053 17491
rect 162517 17195 162813 17491
rect 163277 17195 163573 17491
rect 164037 17195 164333 17491
rect 164797 17195 165093 17491
rect 165557 17195 165853 17491
rect 166317 17195 166613 17491
rect 167077 17195 167373 17491
rect 167837 17195 168133 17491
rect 168597 17195 168893 17491
rect 169357 17195 169653 17491
rect 170117 17195 170413 17491
rect 170877 17195 171173 17491
rect 171637 17195 171933 17491
rect 172397 17195 172693 17491
rect 173157 17195 173453 17491
rect 173917 17195 174213 17491
rect 174677 17195 174973 17491
rect 175437 17195 175733 17491
rect 176197 17195 176493 17491
rect 157957 16435 158253 16731
rect 158717 16435 159013 16731
rect 159477 16435 159773 16731
rect 160237 16435 160533 16731
rect 160997 16435 161293 16731
rect 161757 16435 162053 16731
rect 162517 16435 162813 16731
rect 163277 16435 163573 16731
rect 164037 16435 164333 16731
rect 164797 16435 165093 16731
rect 165557 16435 165853 16731
rect 166317 16435 166613 16731
rect 167077 16435 167373 16731
rect 167837 16435 168133 16731
rect 168597 16435 168893 16731
rect 169357 16435 169653 16731
rect 170117 16435 170413 16731
rect 170877 16435 171173 16731
rect 171637 16435 171933 16731
rect 172397 16435 172693 16731
rect 173157 16435 173453 16731
rect 173917 16435 174213 16731
rect 174677 16435 174973 16731
rect 175437 16435 175733 16731
rect 176197 16435 176493 16731
rect 157957 15675 158253 15971
rect 158717 15675 159013 15971
rect 159477 15675 159773 15971
rect 160237 15675 160533 15971
rect 160997 15675 161293 15971
rect 161757 15675 162053 15971
rect 162517 15675 162813 15971
rect 163277 15675 163573 15971
rect 164037 15675 164333 15971
rect 164797 15675 165093 15971
rect 165557 15675 165853 15971
rect 166317 15675 166613 15971
rect 167077 15675 167373 15971
rect 167837 15675 168133 15971
rect 168597 15675 168893 15971
rect 169357 15675 169653 15971
rect 170117 15675 170413 15971
rect 170877 15675 171173 15971
rect 171637 15675 171933 15971
rect 172397 15675 172693 15971
rect 173157 15675 173453 15971
rect 173917 15675 174213 15971
rect 174677 15675 174973 15971
rect 175437 15675 175733 15971
rect 176197 15675 176493 15971
rect 157957 14915 158253 15211
rect 158717 14915 159013 15211
rect 159477 14915 159773 15211
rect 160237 14915 160533 15211
rect 160997 14915 161293 15211
rect 161757 14915 162053 15211
rect 162517 14915 162813 15211
rect 163277 14915 163573 15211
rect 164037 14915 164333 15211
rect 164797 14915 165093 15211
rect 165557 14915 165853 15211
rect 166317 14915 166613 15211
rect 167077 14915 167373 15211
rect 167837 14915 168133 15211
rect 168597 14915 168893 15211
rect 169357 14915 169653 15211
rect 170117 14915 170413 15211
rect 170877 14915 171173 15211
rect 171637 14915 171933 15211
rect 172397 14915 172693 15211
rect 173157 14915 173453 15211
rect 173917 14915 174213 15211
rect 174677 14915 174973 15211
rect 175437 14915 175733 15211
rect 176197 14915 176493 15211
rect 157957 14155 158253 14451
rect 158717 14155 159013 14451
rect 159477 14155 159773 14451
rect 160237 14155 160533 14451
rect 160997 14155 161293 14451
rect 161757 14155 162053 14451
rect 162517 14155 162813 14451
rect 163277 14155 163573 14451
rect 164037 14155 164333 14451
rect 164797 14155 165093 14451
rect 165557 14155 165853 14451
rect 166317 14155 166613 14451
rect 167077 14155 167373 14451
rect 167837 14155 168133 14451
rect 168597 14155 168893 14451
rect 169357 14155 169653 14451
rect 170117 14155 170413 14451
rect 170877 14155 171173 14451
rect 171637 14155 171933 14451
rect 172397 14155 172693 14451
rect 173157 14155 173453 14451
rect 173917 14155 174213 14451
rect 174677 14155 174973 14451
rect 175437 14155 175733 14451
rect 176197 14155 176493 14451
rect 157957 13395 158253 13691
rect 158717 13395 159013 13691
rect 159477 13395 159773 13691
rect 160237 13395 160533 13691
rect 160997 13395 161293 13691
rect 161757 13395 162053 13691
rect 162517 13395 162813 13691
rect 163277 13395 163573 13691
rect 164037 13395 164333 13691
rect 164797 13395 165093 13691
rect 165557 13395 165853 13691
rect 166317 13395 166613 13691
rect 167077 13395 167373 13691
rect 167837 13395 168133 13691
rect 168597 13395 168893 13691
rect 169357 13395 169653 13691
rect 170117 13395 170413 13691
rect 170877 13395 171173 13691
rect 171637 13395 171933 13691
rect 172397 13395 172693 13691
rect 173157 13395 173453 13691
rect 173917 13395 174213 13691
rect 174677 13395 174973 13691
rect 175437 13395 175733 13691
rect 176197 13395 176493 13691
rect 157957 12635 158253 12931
rect 158717 12635 159013 12931
rect 159477 12635 159773 12931
rect 160237 12635 160533 12931
rect 160997 12635 161293 12931
rect 161757 12635 162053 12931
rect 162517 12635 162813 12931
rect 163277 12635 163573 12931
rect 164037 12635 164333 12931
rect 164797 12635 165093 12931
rect 165557 12635 165853 12931
rect 166317 12635 166613 12931
rect 167077 12635 167373 12931
rect 167837 12635 168133 12931
rect 168597 12635 168893 12931
rect 169357 12635 169653 12931
rect 170117 12635 170413 12931
rect 170877 12635 171173 12931
rect 171637 12635 171933 12931
rect 172397 12635 172693 12931
rect 173157 12635 173453 12931
rect 173917 12635 174213 12931
rect 174677 12635 174973 12931
rect 175437 12635 175733 12931
rect 176197 12635 176493 12931
rect 157957 11875 158253 12171
rect 158717 11875 159013 12171
rect 159477 11875 159773 12171
rect 160237 11875 160533 12171
rect 160997 11875 161293 12171
rect 161757 11875 162053 12171
rect 162517 11875 162813 12171
rect 163277 11875 163573 12171
rect 164037 11875 164333 12171
rect 164797 11875 165093 12171
rect 165557 11875 165853 12171
rect 166317 11875 166613 12171
rect 167077 11875 167373 12171
rect 167837 11875 168133 12171
rect 168597 11875 168893 12171
rect 169357 11875 169653 12171
rect 170117 11875 170413 12171
rect 170877 11875 171173 12171
rect 171637 11875 171933 12171
rect 172397 11875 172693 12171
rect 173157 11875 173453 12171
rect 173917 11875 174213 12171
rect 174677 11875 174973 12171
rect 175437 11875 175733 12171
rect 176197 11875 176493 12171
rect 157957 11115 158253 11411
rect 158717 11115 159013 11411
rect 159477 11115 159773 11411
rect 160237 11115 160533 11411
rect 160997 11115 161293 11411
rect 161757 11115 162053 11411
rect 162517 11115 162813 11411
rect 163277 11115 163573 11411
rect 164037 11115 164333 11411
rect 164797 11115 165093 11411
rect 165557 11115 165853 11411
rect 166317 11115 166613 11411
rect 167077 11115 167373 11411
rect 167837 11115 168133 11411
rect 168597 11115 168893 11411
rect 169357 11115 169653 11411
rect 170117 11115 170413 11411
rect 170877 11115 171173 11411
rect 171637 11115 171933 11411
rect 172397 11115 172693 11411
rect 173157 11115 173453 11411
rect 173917 11115 174213 11411
rect 174677 11115 174973 11411
rect 175437 11115 175733 11411
rect 176197 11115 176493 11411
rect 157957 10355 158253 10651
rect 158717 10355 159013 10651
rect 159477 10355 159773 10651
rect 160237 10355 160533 10651
rect 160997 10355 161293 10651
rect 161757 10355 162053 10651
rect 162517 10355 162813 10651
rect 163277 10355 163573 10651
rect 164037 10355 164333 10651
rect 164797 10355 165093 10651
rect 165557 10355 165853 10651
rect 166317 10355 166613 10651
rect 167077 10355 167373 10651
rect 167837 10355 168133 10651
rect 168597 10355 168893 10651
rect 169357 10355 169653 10651
rect 170117 10355 170413 10651
rect 170877 10355 171173 10651
rect 171637 10355 171933 10651
rect 172397 10355 172693 10651
rect 173157 10355 173453 10651
rect 173917 10355 174213 10651
rect 174677 10355 174973 10651
rect 175437 10355 175733 10651
rect 176197 10355 176493 10651
rect 157957 9595 158253 9891
rect 158717 9595 159013 9891
rect 159477 9595 159773 9891
rect 160237 9595 160533 9891
rect 160997 9595 161293 9891
rect 161757 9595 162053 9891
rect 162517 9595 162813 9891
rect 163277 9595 163573 9891
rect 164037 9595 164333 9891
rect 164797 9595 165093 9891
rect 165557 9595 165853 9891
rect 166317 9595 166613 9891
rect 167077 9595 167373 9891
rect 167837 9595 168133 9891
rect 168597 9595 168893 9891
rect 169357 9595 169653 9891
rect 170117 9595 170413 9891
rect 170877 9595 171173 9891
rect 171637 9595 171933 9891
rect 172397 9595 172693 9891
rect 173157 9595 173453 9891
rect 173917 9595 174213 9891
rect 174677 9595 174973 9891
rect 175437 9595 175733 9891
rect 176197 9595 176493 9891
rect 157957 8835 158253 9131
rect 158717 8835 159013 9131
rect 159477 8835 159773 9131
rect 160237 8835 160533 9131
rect 160997 8835 161293 9131
rect 161757 8835 162053 9131
rect 162517 8835 162813 9131
rect 163277 8835 163573 9131
rect 164037 8835 164333 9131
rect 164797 8835 165093 9131
rect 165557 8835 165853 9131
rect 166317 8835 166613 9131
rect 167077 8835 167373 9131
rect 167837 8835 168133 9131
rect 168597 8835 168893 9131
rect 169357 8835 169653 9131
rect 170117 8835 170413 9131
rect 170877 8835 171173 9131
rect 171637 8835 171933 9131
rect 172397 8835 172693 9131
rect 173157 8835 173453 9131
rect 173917 8835 174213 9131
rect 174677 8835 174973 9131
rect 175437 8835 175733 9131
rect 176197 8835 176493 9131
rect 157957 8075 158253 8371
rect 158717 8075 159013 8371
rect 159477 8075 159773 8371
rect 160237 8075 160533 8371
rect 160997 8075 161293 8371
rect 161757 8075 162053 8371
rect 162517 8075 162813 8371
rect 163277 8075 163573 8371
rect 164037 8075 164333 8371
rect 164797 8075 165093 8371
rect 165557 8075 165853 8371
rect 166317 8075 166613 8371
rect 167077 8075 167373 8371
rect 167837 8075 168133 8371
rect 168597 8075 168893 8371
rect 169357 8075 169653 8371
rect 170117 8075 170413 8371
rect 170877 8075 171173 8371
rect 171637 8075 171933 8371
rect 172397 8075 172693 8371
rect 173157 8075 173453 8371
rect 173917 8075 174213 8371
rect 174677 8075 174973 8371
rect 175437 8075 175733 8371
rect 176197 8075 176493 8371
rect 157957 7315 158253 7611
rect 158717 7315 159013 7611
rect 159477 7315 159773 7611
rect 160237 7315 160533 7611
rect 160997 7315 161293 7611
rect 161757 7315 162053 7611
rect 162517 7315 162813 7611
rect 163277 7315 163573 7611
rect 164037 7315 164333 7611
rect 164797 7315 165093 7611
rect 165557 7315 165853 7611
rect 166317 7315 166613 7611
rect 167077 7315 167373 7611
rect 167837 7315 168133 7611
rect 168597 7315 168893 7611
rect 169357 7315 169653 7611
rect 170117 7315 170413 7611
rect 170877 7315 171173 7611
rect 171637 7315 171933 7611
rect 172397 7315 172693 7611
rect 173157 7315 173453 7611
rect 173917 7315 174213 7611
rect 174677 7315 174973 7611
rect 175437 7315 175733 7611
rect 176197 7315 176493 7611
rect 187077 28688 187373 28984
rect 187837 28688 188133 28984
rect 188597 28688 188893 28984
rect 189357 28688 189653 28984
rect 190117 28688 190413 28984
rect 190877 28688 191173 28984
rect 191637 28688 191933 28984
rect 192397 28688 192693 28984
rect 193157 28688 193453 28984
rect 193917 28688 194213 28984
rect 194677 28688 194973 28984
rect 195437 28688 195733 28984
rect 196197 28688 196493 28984
rect 196957 28688 197253 28984
rect 197717 28688 198013 28984
rect 198477 28688 198773 28984
rect 199237 28688 199533 28984
rect 199997 28688 200293 28984
rect 200757 28688 201053 28984
rect 201517 28688 201813 28984
rect 202277 28688 202573 28984
rect 203037 28688 203333 28984
rect 203797 28688 204093 28984
rect 204557 28688 204853 28984
rect 205317 28688 205613 28984
rect 206077 28688 206373 28984
rect 206837 28688 207133 28984
rect 207597 28688 207893 28984
rect 208357 28688 208653 28984
rect 209117 28688 209413 28984
rect 209877 28688 210173 28984
rect 210637 28688 210933 28984
rect 187077 27928 187373 28224
rect 187837 27928 188133 28224
rect 188597 27928 188893 28224
rect 189357 27928 189653 28224
rect 190117 27928 190413 28224
rect 190877 27928 191173 28224
rect 191637 27928 191933 28224
rect 192397 27928 192693 28224
rect 193157 27928 193453 28224
rect 193917 27928 194213 28224
rect 194677 27928 194973 28224
rect 195437 27928 195733 28224
rect 196197 27928 196493 28224
rect 196957 27928 197253 28224
rect 197717 27928 198013 28224
rect 198477 27928 198773 28224
rect 199237 27928 199533 28224
rect 199997 27928 200293 28224
rect 200757 27928 201053 28224
rect 201517 27928 201813 28224
rect 202277 27928 202573 28224
rect 203037 27928 203333 28224
rect 203797 27928 204093 28224
rect 204557 27928 204853 28224
rect 205317 27928 205613 28224
rect 206077 27928 206373 28224
rect 206837 27928 207133 28224
rect 207597 27928 207893 28224
rect 208357 27928 208653 28224
rect 209117 27928 209413 28224
rect 209877 27928 210173 28224
rect 210637 27928 210933 28224
rect 187077 27168 187373 27464
rect 187837 27168 188133 27464
rect 188597 27168 188893 27464
rect 189357 27168 189653 27464
rect 190117 27168 190413 27464
rect 190877 27168 191173 27464
rect 191637 27168 191933 27464
rect 192397 27168 192693 27464
rect 193157 27168 193453 27464
rect 193917 27168 194213 27464
rect 194677 27168 194973 27464
rect 195437 27168 195733 27464
rect 196197 27168 196493 27464
rect 196957 27168 197253 27464
rect 197717 27168 198013 27464
rect 198477 27168 198773 27464
rect 199237 27168 199533 27464
rect 199997 27168 200293 27464
rect 200757 27168 201053 27464
rect 201517 27168 201813 27464
rect 202277 27168 202573 27464
rect 203037 27168 203333 27464
rect 203797 27168 204093 27464
rect 204557 27168 204853 27464
rect 205317 27168 205613 27464
rect 206077 27168 206373 27464
rect 206837 27168 207133 27464
rect 207597 27168 207893 27464
rect 208357 27168 208653 27464
rect 209117 27168 209413 27464
rect 209877 27168 210173 27464
rect 210637 27168 210933 27464
rect 187077 26408 187373 26704
rect 187837 26408 188133 26704
rect 188597 26408 188893 26704
rect 189357 26408 189653 26704
rect 190117 26408 190413 26704
rect 190877 26408 191173 26704
rect 191637 26408 191933 26704
rect 192397 26408 192693 26704
rect 193157 26408 193453 26704
rect 193917 26408 194213 26704
rect 194677 26408 194973 26704
rect 195437 26408 195733 26704
rect 196197 26408 196493 26704
rect 196957 26408 197253 26704
rect 197717 26408 198013 26704
rect 198477 26408 198773 26704
rect 199237 26408 199533 26704
rect 199997 26408 200293 26704
rect 200757 26408 201053 26704
rect 201517 26408 201813 26704
rect 202277 26408 202573 26704
rect 203037 26408 203333 26704
rect 203797 26408 204093 26704
rect 204557 26408 204853 26704
rect 205317 26408 205613 26704
rect 206077 26408 206373 26704
rect 206837 26408 207133 26704
rect 207597 26408 207893 26704
rect 208357 26408 208653 26704
rect 209117 26408 209413 26704
rect 209877 26408 210173 26704
rect 210637 26408 210933 26704
rect 187077 25648 187373 25944
rect 187837 25648 188133 25944
rect 188597 25648 188893 25944
rect 189357 25648 189653 25944
rect 190117 25648 190413 25944
rect 190877 25648 191173 25944
rect 191637 25648 191933 25944
rect 192397 25648 192693 25944
rect 193157 25648 193453 25944
rect 193917 25648 194213 25944
rect 194677 25648 194973 25944
rect 195437 25648 195733 25944
rect 196197 25648 196493 25944
rect 196957 25648 197253 25944
rect 197717 25648 198013 25944
rect 198477 25648 198773 25944
rect 199237 25648 199533 25944
rect 199997 25648 200293 25944
rect 200757 25648 201053 25944
rect 201517 25648 201813 25944
rect 202277 25648 202573 25944
rect 203037 25648 203333 25944
rect 203797 25648 204093 25944
rect 204557 25648 204853 25944
rect 205317 25648 205613 25944
rect 206077 25648 206373 25944
rect 206837 25648 207133 25944
rect 207597 25648 207893 25944
rect 208357 25648 208653 25944
rect 209117 25648 209413 25944
rect 209877 25648 210173 25944
rect 210637 25648 210933 25944
rect 187077 24888 187373 25184
rect 187837 24888 188133 25184
rect 188597 24888 188893 25184
rect 189357 24888 189653 25184
rect 190117 24888 190413 25184
rect 190877 24888 191173 25184
rect 191637 24888 191933 25184
rect 192397 24888 192693 25184
rect 193157 24888 193453 25184
rect 193917 24888 194213 25184
rect 194677 24888 194973 25184
rect 195437 24888 195733 25184
rect 196197 24888 196493 25184
rect 196957 24888 197253 25184
rect 197717 24888 198013 25184
rect 198477 24888 198773 25184
rect 199237 24888 199533 25184
rect 199997 24888 200293 25184
rect 200757 24888 201053 25184
rect 201517 24888 201813 25184
rect 202277 24888 202573 25184
rect 203037 24888 203333 25184
rect 203797 24888 204093 25184
rect 204557 24888 204853 25184
rect 205317 24888 205613 25184
rect 206077 24888 206373 25184
rect 206837 24888 207133 25184
rect 207597 24888 207893 25184
rect 208357 24888 208653 25184
rect 209117 24888 209413 25184
rect 209877 24888 210173 25184
rect 210637 24888 210933 25184
rect 187077 24128 187373 24424
rect 187837 24128 188133 24424
rect 188597 24128 188893 24424
rect 189357 24128 189653 24424
rect 190117 24128 190413 24424
rect 190877 24128 191173 24424
rect 191637 24128 191933 24424
rect 192397 24128 192693 24424
rect 193157 24128 193453 24424
rect 193917 24128 194213 24424
rect 194677 24128 194973 24424
rect 195437 24128 195733 24424
rect 196197 24128 196493 24424
rect 196957 24128 197253 24424
rect 197717 24128 198013 24424
rect 198477 24128 198773 24424
rect 199237 24128 199533 24424
rect 199997 24128 200293 24424
rect 200757 24128 201053 24424
rect 201517 24128 201813 24424
rect 202277 24128 202573 24424
rect 203037 24128 203333 24424
rect 203797 24128 204093 24424
rect 204557 24128 204853 24424
rect 205317 24128 205613 24424
rect 206077 24128 206373 24424
rect 206837 24128 207133 24424
rect 207597 24128 207893 24424
rect 208357 24128 208653 24424
rect 209117 24128 209413 24424
rect 209877 24128 210173 24424
rect 210637 24128 210933 24424
rect 187077 23368 187373 23664
rect 187837 23368 188133 23664
rect 188597 23368 188893 23664
rect 189357 23368 189653 23664
rect 190117 23368 190413 23664
rect 190877 23368 191173 23664
rect 191637 23368 191933 23664
rect 192397 23368 192693 23664
rect 193157 23368 193453 23664
rect 193917 23368 194213 23664
rect 194677 23368 194973 23664
rect 195437 23368 195733 23664
rect 196197 23368 196493 23664
rect 196957 23368 197253 23664
rect 197717 23368 198013 23664
rect 198477 23368 198773 23664
rect 199237 23368 199533 23664
rect 199997 23368 200293 23664
rect 200757 23368 201053 23664
rect 201517 23368 201813 23664
rect 202277 23368 202573 23664
rect 203037 23368 203333 23664
rect 203797 23368 204093 23664
rect 204557 23368 204853 23664
rect 205317 23368 205613 23664
rect 206077 23368 206373 23664
rect 206837 23368 207133 23664
rect 207597 23368 207893 23664
rect 208357 23368 208653 23664
rect 209117 23368 209413 23664
rect 209877 23368 210173 23664
rect 210637 23368 210933 23664
rect 187077 22608 187373 22904
rect 187837 22608 188133 22904
rect 188597 22608 188893 22904
rect 189357 22608 189653 22904
rect 190117 22608 190413 22904
rect 190877 22608 191173 22904
rect 191637 22608 191933 22904
rect 192397 22608 192693 22904
rect 193157 22608 193453 22904
rect 193917 22608 194213 22904
rect 194677 22608 194973 22904
rect 195437 22608 195733 22904
rect 196197 22608 196493 22904
rect 196957 22608 197253 22904
rect 197717 22608 198013 22904
rect 198477 22608 198773 22904
rect 199237 22608 199533 22904
rect 199997 22608 200293 22904
rect 200757 22608 201053 22904
rect 201517 22608 201813 22904
rect 202277 22608 202573 22904
rect 203037 22608 203333 22904
rect 203797 22608 204093 22904
rect 204557 22608 204853 22904
rect 205317 22608 205613 22904
rect 206077 22608 206373 22904
rect 206837 22608 207133 22904
rect 207597 22608 207893 22904
rect 208357 22608 208653 22904
rect 209117 22608 209413 22904
rect 209877 22608 210173 22904
rect 210637 22608 210933 22904
rect 187077 21848 187373 22144
rect 187837 21848 188133 22144
rect 188597 21848 188893 22144
rect 189357 21848 189653 22144
rect 190117 21848 190413 22144
rect 190877 21848 191173 22144
rect 191637 21848 191933 22144
rect 192397 21848 192693 22144
rect 193157 21848 193453 22144
rect 193917 21848 194213 22144
rect 194677 21848 194973 22144
rect 195437 21848 195733 22144
rect 196197 21848 196493 22144
rect 196957 21848 197253 22144
rect 197717 21848 198013 22144
rect 198477 21848 198773 22144
rect 199237 21848 199533 22144
rect 199997 21848 200293 22144
rect 200757 21848 201053 22144
rect 201517 21848 201813 22144
rect 202277 21848 202573 22144
rect 203037 21848 203333 22144
rect 203797 21848 204093 22144
rect 204557 21848 204853 22144
rect 205317 21848 205613 22144
rect 206077 21848 206373 22144
rect 206837 21848 207133 22144
rect 207597 21848 207893 22144
rect 208357 21848 208653 22144
rect 209117 21848 209413 22144
rect 209877 21848 210173 22144
rect 210637 21848 210933 22144
rect 187077 21088 187373 21384
rect 187837 21088 188133 21384
rect 188597 21088 188893 21384
rect 189357 21088 189653 21384
rect 190117 21088 190413 21384
rect 190877 21088 191173 21384
rect 191637 21088 191933 21384
rect 192397 21088 192693 21384
rect 193157 21088 193453 21384
rect 193917 21088 194213 21384
rect 194677 21088 194973 21384
rect 195437 21088 195733 21384
rect 196197 21088 196493 21384
rect 196957 21088 197253 21384
rect 197717 21088 198013 21384
rect 198477 21088 198773 21384
rect 199237 21088 199533 21384
rect 199997 21088 200293 21384
rect 200757 21088 201053 21384
rect 201517 21088 201813 21384
rect 202277 21088 202573 21384
rect 203037 21088 203333 21384
rect 203797 21088 204093 21384
rect 204557 21088 204853 21384
rect 205317 21088 205613 21384
rect 206077 21088 206373 21384
rect 206837 21088 207133 21384
rect 207597 21088 207893 21384
rect 208357 21088 208653 21384
rect 209117 21088 209413 21384
rect 209877 21088 210173 21384
rect 210637 21088 210933 21384
rect 187077 20328 187373 20624
rect 187837 20328 188133 20624
rect 188597 20328 188893 20624
rect 189357 20328 189653 20624
rect 190117 20328 190413 20624
rect 190877 20328 191173 20624
rect 191637 20328 191933 20624
rect 192397 20328 192693 20624
rect 193157 20328 193453 20624
rect 193917 20328 194213 20624
rect 194677 20328 194973 20624
rect 195437 20328 195733 20624
rect 196197 20328 196493 20624
rect 196957 20328 197253 20624
rect 197717 20328 198013 20624
rect 198477 20328 198773 20624
rect 199237 20328 199533 20624
rect 199997 20328 200293 20624
rect 200757 20328 201053 20624
rect 201517 20328 201813 20624
rect 202277 20328 202573 20624
rect 203037 20328 203333 20624
rect 203797 20328 204093 20624
rect 204557 20328 204853 20624
rect 205317 20328 205613 20624
rect 206077 20328 206373 20624
rect 206837 20328 207133 20624
rect 207597 20328 207893 20624
rect 208357 20328 208653 20624
rect 209117 20328 209413 20624
rect 209877 20328 210173 20624
rect 210637 20328 210933 20624
rect 187077 19568 187373 19864
rect 187837 19568 188133 19864
rect 188597 19568 188893 19864
rect 189357 19568 189653 19864
rect 190117 19568 190413 19864
rect 190877 19568 191173 19864
rect 191637 19568 191933 19864
rect 192397 19568 192693 19864
rect 193157 19568 193453 19864
rect 193917 19568 194213 19864
rect 194677 19568 194973 19864
rect 195437 19568 195733 19864
rect 196197 19568 196493 19864
rect 196957 19568 197253 19864
rect 197717 19568 198013 19864
rect 198477 19568 198773 19864
rect 199237 19568 199533 19864
rect 199997 19568 200293 19864
rect 200757 19568 201053 19864
rect 201517 19568 201813 19864
rect 202277 19568 202573 19864
rect 203037 19568 203333 19864
rect 203797 19568 204093 19864
rect 204557 19568 204853 19864
rect 205317 19568 205613 19864
rect 206077 19568 206373 19864
rect 206837 19568 207133 19864
rect 207597 19568 207893 19864
rect 208357 19568 208653 19864
rect 209117 19568 209413 19864
rect 209877 19568 210173 19864
rect 210637 19568 210933 19864
rect 187077 18808 187373 19104
rect 187837 18808 188133 19104
rect 188597 18808 188893 19104
rect 189357 18808 189653 19104
rect 190117 18808 190413 19104
rect 190877 18808 191173 19104
rect 191637 18808 191933 19104
rect 192397 18808 192693 19104
rect 193157 18808 193453 19104
rect 193917 18808 194213 19104
rect 194677 18808 194973 19104
rect 195437 18808 195733 19104
rect 196197 18808 196493 19104
rect 196957 18808 197253 19104
rect 197717 18808 198013 19104
rect 198477 18808 198773 19104
rect 199237 18808 199533 19104
rect 199997 18808 200293 19104
rect 200757 18808 201053 19104
rect 201517 18808 201813 19104
rect 202277 18808 202573 19104
rect 203037 18808 203333 19104
rect 203797 18808 204093 19104
rect 204557 18808 204853 19104
rect 205317 18808 205613 19104
rect 206077 18808 206373 19104
rect 206837 18808 207133 19104
rect 207597 18808 207893 19104
rect 208357 18808 208653 19104
rect 209117 18808 209413 19104
rect 209877 18808 210173 19104
rect 210637 18808 210933 19104
rect 187077 18048 187373 18344
rect 187837 18048 188133 18344
rect 188597 18048 188893 18344
rect 189357 18048 189653 18344
rect 190117 18048 190413 18344
rect 190877 18048 191173 18344
rect 191637 18048 191933 18344
rect 192397 18048 192693 18344
rect 193157 18048 193453 18344
rect 193917 18048 194213 18344
rect 194677 18048 194973 18344
rect 195437 18048 195733 18344
rect 196197 18048 196493 18344
rect 196957 18048 197253 18344
rect 197717 18048 198013 18344
rect 198477 18048 198773 18344
rect 199237 18048 199533 18344
rect 199997 18048 200293 18344
rect 200757 18048 201053 18344
rect 201517 18048 201813 18344
rect 202277 18048 202573 18344
rect 203037 18048 203333 18344
rect 203797 18048 204093 18344
rect 204557 18048 204853 18344
rect 205317 18048 205613 18344
rect 206077 18048 206373 18344
rect 206837 18048 207133 18344
rect 207597 18048 207893 18344
rect 208357 18048 208653 18344
rect 209117 18048 209413 18344
rect 209877 18048 210173 18344
rect 210637 18048 210933 18344
rect 187077 17288 187373 17584
rect 187837 17288 188133 17584
rect 188597 17288 188893 17584
rect 189357 17288 189653 17584
rect 190117 17288 190413 17584
rect 190877 17288 191173 17584
rect 191637 17288 191933 17584
rect 192397 17288 192693 17584
rect 193157 17288 193453 17584
rect 193917 17288 194213 17584
rect 194677 17288 194973 17584
rect 195437 17288 195733 17584
rect 196197 17288 196493 17584
rect 196957 17288 197253 17584
rect 197717 17288 198013 17584
rect 198477 17288 198773 17584
rect 199237 17288 199533 17584
rect 199997 17288 200293 17584
rect 200757 17288 201053 17584
rect 201517 17288 201813 17584
rect 202277 17288 202573 17584
rect 203037 17288 203333 17584
rect 203797 17288 204093 17584
rect 204557 17288 204853 17584
rect 205317 17288 205613 17584
rect 206077 17288 206373 17584
rect 206837 17288 207133 17584
rect 207597 17288 207893 17584
rect 208357 17288 208653 17584
rect 209117 17288 209413 17584
rect 209877 17288 210173 17584
rect 210637 17288 210933 17584
rect 187077 16528 187373 16824
rect 187837 16528 188133 16824
rect 188597 16528 188893 16824
rect 189357 16528 189653 16824
rect 190117 16528 190413 16824
rect 190877 16528 191173 16824
rect 191637 16528 191933 16824
rect 192397 16528 192693 16824
rect 193157 16528 193453 16824
rect 193917 16528 194213 16824
rect 194677 16528 194973 16824
rect 195437 16528 195733 16824
rect 196197 16528 196493 16824
rect 196957 16528 197253 16824
rect 197717 16528 198013 16824
rect 198477 16528 198773 16824
rect 199237 16528 199533 16824
rect 199997 16528 200293 16824
rect 200757 16528 201053 16824
rect 201517 16528 201813 16824
rect 202277 16528 202573 16824
rect 203037 16528 203333 16824
rect 203797 16528 204093 16824
rect 204557 16528 204853 16824
rect 205317 16528 205613 16824
rect 206077 16528 206373 16824
rect 206837 16528 207133 16824
rect 207597 16528 207893 16824
rect 208357 16528 208653 16824
rect 209117 16528 209413 16824
rect 209877 16528 210173 16824
rect 210637 16528 210933 16824
rect 187077 15768 187373 16064
rect 187837 15768 188133 16064
rect 188597 15768 188893 16064
rect 189357 15768 189653 16064
rect 190117 15768 190413 16064
rect 190877 15768 191173 16064
rect 191637 15768 191933 16064
rect 192397 15768 192693 16064
rect 193157 15768 193453 16064
rect 193917 15768 194213 16064
rect 194677 15768 194973 16064
rect 195437 15768 195733 16064
rect 196197 15768 196493 16064
rect 196957 15768 197253 16064
rect 197717 15768 198013 16064
rect 198477 15768 198773 16064
rect 199237 15768 199533 16064
rect 199997 15768 200293 16064
rect 200757 15768 201053 16064
rect 201517 15768 201813 16064
rect 202277 15768 202573 16064
rect 203037 15768 203333 16064
rect 203797 15768 204093 16064
rect 204557 15768 204853 16064
rect 205317 15768 205613 16064
rect 206077 15768 206373 16064
rect 206837 15768 207133 16064
rect 207597 15768 207893 16064
rect 208357 15768 208653 16064
rect 209117 15768 209413 16064
rect 209877 15768 210173 16064
rect 210637 15768 210933 16064
rect 187077 15008 187373 15304
rect 187837 15008 188133 15304
rect 188597 15008 188893 15304
rect 189357 15008 189653 15304
rect 190117 15008 190413 15304
rect 190877 15008 191173 15304
rect 191637 15008 191933 15304
rect 192397 15008 192693 15304
rect 193157 15008 193453 15304
rect 193917 15008 194213 15304
rect 194677 15008 194973 15304
rect 195437 15008 195733 15304
rect 196197 15008 196493 15304
rect 196957 15008 197253 15304
rect 197717 15008 198013 15304
rect 198477 15008 198773 15304
rect 199237 15008 199533 15304
rect 199997 15008 200293 15304
rect 200757 15008 201053 15304
rect 201517 15008 201813 15304
rect 202277 15008 202573 15304
rect 203037 15008 203333 15304
rect 203797 15008 204093 15304
rect 204557 15008 204853 15304
rect 205317 15008 205613 15304
rect 206077 15008 206373 15304
rect 206837 15008 207133 15304
rect 207597 15008 207893 15304
rect 208357 15008 208653 15304
rect 209117 15008 209413 15304
rect 209877 15008 210173 15304
rect 210637 15008 210933 15304
rect 187077 14248 187373 14544
rect 187837 14248 188133 14544
rect 188597 14248 188893 14544
rect 189357 14248 189653 14544
rect 190117 14248 190413 14544
rect 190877 14248 191173 14544
rect 191637 14248 191933 14544
rect 192397 14248 192693 14544
rect 193157 14248 193453 14544
rect 193917 14248 194213 14544
rect 194677 14248 194973 14544
rect 195437 14248 195733 14544
rect 196197 14248 196493 14544
rect 196957 14248 197253 14544
rect 197717 14248 198013 14544
rect 198477 14248 198773 14544
rect 199237 14248 199533 14544
rect 199997 14248 200293 14544
rect 200757 14248 201053 14544
rect 201517 14248 201813 14544
rect 202277 14248 202573 14544
rect 203037 14248 203333 14544
rect 203797 14248 204093 14544
rect 204557 14248 204853 14544
rect 205317 14248 205613 14544
rect 206077 14248 206373 14544
rect 206837 14248 207133 14544
rect 207597 14248 207893 14544
rect 208357 14248 208653 14544
rect 209117 14248 209413 14544
rect 209877 14248 210173 14544
rect 210637 14248 210933 14544
rect 187077 13488 187373 13784
rect 187837 13488 188133 13784
rect 188597 13488 188893 13784
rect 189357 13488 189653 13784
rect 190117 13488 190413 13784
rect 190877 13488 191173 13784
rect 191637 13488 191933 13784
rect 192397 13488 192693 13784
rect 193157 13488 193453 13784
rect 193917 13488 194213 13784
rect 194677 13488 194973 13784
rect 195437 13488 195733 13784
rect 196197 13488 196493 13784
rect 196957 13488 197253 13784
rect 197717 13488 198013 13784
rect 198477 13488 198773 13784
rect 199237 13488 199533 13784
rect 199997 13488 200293 13784
rect 200757 13488 201053 13784
rect 201517 13488 201813 13784
rect 202277 13488 202573 13784
rect 203037 13488 203333 13784
rect 203797 13488 204093 13784
rect 204557 13488 204853 13784
rect 205317 13488 205613 13784
rect 206077 13488 206373 13784
rect 206837 13488 207133 13784
rect 207597 13488 207893 13784
rect 208357 13488 208653 13784
rect 209117 13488 209413 13784
rect 209877 13488 210173 13784
rect 210637 13488 210933 13784
rect 187077 12728 187373 13024
rect 187837 12728 188133 13024
rect 188597 12728 188893 13024
rect 189357 12728 189653 13024
rect 190117 12728 190413 13024
rect 190877 12728 191173 13024
rect 191637 12728 191933 13024
rect 192397 12728 192693 13024
rect 193157 12728 193453 13024
rect 193917 12728 194213 13024
rect 194677 12728 194973 13024
rect 195437 12728 195733 13024
rect 196197 12728 196493 13024
rect 196957 12728 197253 13024
rect 197717 12728 198013 13024
rect 198477 12728 198773 13024
rect 199237 12728 199533 13024
rect 199997 12728 200293 13024
rect 200757 12728 201053 13024
rect 201517 12728 201813 13024
rect 202277 12728 202573 13024
rect 203037 12728 203333 13024
rect 203797 12728 204093 13024
rect 204557 12728 204853 13024
rect 205317 12728 205613 13024
rect 206077 12728 206373 13024
rect 206837 12728 207133 13024
rect 207597 12728 207893 13024
rect 208357 12728 208653 13024
rect 209117 12728 209413 13024
rect 209877 12728 210173 13024
rect 210637 12728 210933 13024
rect 187077 11968 187373 12264
rect 187837 11968 188133 12264
rect 188597 11968 188893 12264
rect 189357 11968 189653 12264
rect 190117 11968 190413 12264
rect 190877 11968 191173 12264
rect 191637 11968 191933 12264
rect 192397 11968 192693 12264
rect 193157 11968 193453 12264
rect 193917 11968 194213 12264
rect 194677 11968 194973 12264
rect 195437 11968 195733 12264
rect 196197 11968 196493 12264
rect 196957 11968 197253 12264
rect 197717 11968 198013 12264
rect 198477 11968 198773 12264
rect 199237 11968 199533 12264
rect 199997 11968 200293 12264
rect 200757 11968 201053 12264
rect 201517 11968 201813 12264
rect 202277 11968 202573 12264
rect 203037 11968 203333 12264
rect 203797 11968 204093 12264
rect 204557 11968 204853 12264
rect 205317 11968 205613 12264
rect 206077 11968 206373 12264
rect 206837 11968 207133 12264
rect 207597 11968 207893 12264
rect 208357 11968 208653 12264
rect 209117 11968 209413 12264
rect 209877 11968 210173 12264
rect 210637 11968 210933 12264
rect 187077 11208 187373 11504
rect 187837 11208 188133 11504
rect 188597 11208 188893 11504
rect 189357 11208 189653 11504
rect 190117 11208 190413 11504
rect 190877 11208 191173 11504
rect 191637 11208 191933 11504
rect 192397 11208 192693 11504
rect 193157 11208 193453 11504
rect 193917 11208 194213 11504
rect 194677 11208 194973 11504
rect 195437 11208 195733 11504
rect 196197 11208 196493 11504
rect 196957 11208 197253 11504
rect 197717 11208 198013 11504
rect 198477 11208 198773 11504
rect 199237 11208 199533 11504
rect 199997 11208 200293 11504
rect 200757 11208 201053 11504
rect 201517 11208 201813 11504
rect 202277 11208 202573 11504
rect 203037 11208 203333 11504
rect 203797 11208 204093 11504
rect 204557 11208 204853 11504
rect 205317 11208 205613 11504
rect 206077 11208 206373 11504
rect 206837 11208 207133 11504
rect 207597 11208 207893 11504
rect 208357 11208 208653 11504
rect 209117 11208 209413 11504
rect 209877 11208 210173 11504
rect 210637 11208 210933 11504
rect 187077 10448 187373 10744
rect 187837 10448 188133 10744
rect 188597 10448 188893 10744
rect 189357 10448 189653 10744
rect 190117 10448 190413 10744
rect 190877 10448 191173 10744
rect 191637 10448 191933 10744
rect 192397 10448 192693 10744
rect 193157 10448 193453 10744
rect 193917 10448 194213 10744
rect 194677 10448 194973 10744
rect 195437 10448 195733 10744
rect 196197 10448 196493 10744
rect 196957 10448 197253 10744
rect 197717 10448 198013 10744
rect 198477 10448 198773 10744
rect 199237 10448 199533 10744
rect 199997 10448 200293 10744
rect 200757 10448 201053 10744
rect 201517 10448 201813 10744
rect 202277 10448 202573 10744
rect 203037 10448 203333 10744
rect 203797 10448 204093 10744
rect 204557 10448 204853 10744
rect 205317 10448 205613 10744
rect 206077 10448 206373 10744
rect 206837 10448 207133 10744
rect 207597 10448 207893 10744
rect 208357 10448 208653 10744
rect 209117 10448 209413 10744
rect 209877 10448 210173 10744
rect 210637 10448 210933 10744
<< metal3 >>
rect 178794 16788 180651 17101
rect 178794 16381 179230 16788
rect 179759 16381 180651 16788
rect 178794 9674 180651 16381
rect 178794 9144 179458 9674
rect 180057 9144 180651 9674
rect 178794 8866 180651 9144
rect 188998 8391 192096 8638
rect 188998 7938 189991 8391
rect 190976 7938 192096 8391
rect 188998 6863 192096 7938
rect 188998 6200 190005 6863
rect 191144 6200 192096 6863
rect 188998 5683 192096 6200
rect 121308 4544 124406 4791
rect 121308 4091 122301 4544
rect 123286 4091 124406 4544
rect 121308 3016 124406 4091
rect 121308 2353 122315 3016
rect 123454 2353 124406 3016
rect 121308 1836 124406 2353
<< via3 >>
rect 179230 16381 179759 16788
rect 189991 7938 190976 8391
rect 122301 4091 123286 4544
<< metal4 >>
rect 113025 31743 134225 32343
rect 113025 6743 113625 31743
rect 133625 6743 134225 31743
rect 113025 5605 134225 6743
rect 113025 5341 113613 5605
rect 113877 5341 114133 5605
rect 114397 5341 114653 5605
rect 114917 5341 115173 5605
rect 115437 5341 115693 5605
rect 115957 5341 116213 5605
rect 116477 5341 116733 5605
rect 116997 5341 117253 5605
rect 117517 5341 117773 5605
rect 118037 5341 118293 5605
rect 118557 5341 118813 5605
rect 119077 5341 119333 5605
rect 119597 5341 119853 5605
rect 120117 5341 120373 5605
rect 120637 5341 120893 5605
rect 121157 5341 121413 5605
rect 121677 5341 121933 5605
rect 122197 5341 122453 5605
rect 122717 5341 122973 5605
rect 123237 5341 123493 5605
rect 123757 5341 124013 5605
rect 124277 5341 124533 5605
rect 124797 5341 125053 5605
rect 125317 5341 125573 5605
rect 125837 5341 126093 5605
rect 126357 5341 126613 5605
rect 126877 5341 127133 5605
rect 127397 5341 127653 5605
rect 127917 5341 128173 5605
rect 128437 5341 128693 5605
rect 128957 5341 129213 5605
rect 129477 5341 129733 5605
rect 129997 5341 130253 5605
rect 130517 5341 130773 5605
rect 131037 5341 131293 5605
rect 131557 5341 131813 5605
rect 132077 5341 132333 5605
rect 132597 5341 132853 5605
rect 133117 5341 133373 5605
rect 133637 5341 134225 5605
rect 113025 4943 134225 5341
rect 134825 31743 156025 32343
rect 134825 6743 135425 31743
rect 155425 6743 156025 31743
rect 134825 5605 156025 6743
rect 134825 5341 135413 5605
rect 135677 5341 135933 5605
rect 136197 5341 136453 5605
rect 136717 5341 136973 5605
rect 137237 5341 137493 5605
rect 137757 5341 138013 5605
rect 138277 5341 138533 5605
rect 138797 5341 139053 5605
rect 139317 5341 139573 5605
rect 139837 5341 140093 5605
rect 140357 5341 140613 5605
rect 140877 5341 141133 5605
rect 141397 5341 141653 5605
rect 141917 5341 142173 5605
rect 142437 5341 142693 5605
rect 142957 5341 143213 5605
rect 143477 5341 143733 5605
rect 143997 5341 144253 5605
rect 144517 5341 144773 5605
rect 145037 5341 145293 5605
rect 145557 5341 145813 5605
rect 146077 5341 146333 5605
rect 146597 5341 146853 5605
rect 147117 5341 147373 5605
rect 147637 5341 147893 5605
rect 148157 5341 148413 5605
rect 148677 5341 148933 5605
rect 149197 5341 149453 5605
rect 149717 5341 149973 5605
rect 150237 5341 150493 5605
rect 150757 5341 151013 5605
rect 151277 5341 151533 5605
rect 151797 5341 152053 5605
rect 152317 5341 152573 5605
rect 152837 5341 153093 5605
rect 153357 5341 153613 5605
rect 153877 5341 154133 5605
rect 154397 5341 154653 5605
rect 154917 5341 155173 5605
rect 155437 5341 156025 5605
rect 134825 4943 156025 5341
rect 156625 31743 177825 32343
rect 156625 6743 157225 31743
rect 177225 6743 177825 31743
rect 185905 29728 213305 30316
rect 185905 29716 212643 29728
rect 178794 19469 180493 20255
rect 178794 18992 179090 19469
rect 179707 18992 180493 19469
rect 178794 16788 180493 18992
rect 178794 16381 179230 16788
rect 179759 16381 180493 16788
rect 178794 15787 180493 16381
rect 185905 9716 186505 29716
rect 211505 29464 212643 29716
rect 212907 29464 213305 29728
rect 211505 29208 213305 29464
rect 211505 28944 212643 29208
rect 212907 28944 213305 29208
rect 211505 28688 213305 28944
rect 211505 28424 212643 28688
rect 212907 28424 213305 28688
rect 211505 28168 213305 28424
rect 211505 27904 212643 28168
rect 212907 27904 213305 28168
rect 211505 27648 213305 27904
rect 211505 27384 212643 27648
rect 212907 27384 213305 27648
rect 211505 27128 213305 27384
rect 211505 26864 212643 27128
rect 212907 26864 213305 27128
rect 211505 26608 213305 26864
rect 211505 26344 212643 26608
rect 212907 26344 213305 26608
rect 211505 26088 213305 26344
rect 211505 25824 212643 26088
rect 212907 25824 213305 26088
rect 211505 25568 213305 25824
rect 211505 25304 212643 25568
rect 212907 25304 213305 25568
rect 211505 25048 213305 25304
rect 211505 24784 212643 25048
rect 212907 24784 213305 25048
rect 211505 24528 213305 24784
rect 211505 24264 212643 24528
rect 212907 24264 213305 24528
rect 211505 24008 213305 24264
rect 211505 23744 212643 24008
rect 212907 23744 213305 24008
rect 211505 23488 213305 23744
rect 211505 23224 212643 23488
rect 212907 23224 213305 23488
rect 211505 22968 213305 23224
rect 211505 22704 212643 22968
rect 212907 22704 213305 22968
rect 211505 22448 213305 22704
rect 211505 22184 212643 22448
rect 212907 22184 213305 22448
rect 211505 21928 213305 22184
rect 211505 21664 212643 21928
rect 212907 21664 213305 21928
rect 211505 21408 213305 21664
rect 211505 21144 212643 21408
rect 212907 21144 213305 21408
rect 211505 20888 213305 21144
rect 211505 20624 212643 20888
rect 212907 20624 213305 20888
rect 211505 20368 213305 20624
rect 211505 20104 212643 20368
rect 212907 20104 213305 20368
rect 211505 19848 213305 20104
rect 211505 19584 212643 19848
rect 212907 19584 213305 19848
rect 211505 19328 213305 19584
rect 211505 19064 212643 19328
rect 212907 19064 213305 19328
rect 211505 18808 213305 19064
rect 211505 18544 212643 18808
rect 212907 18544 213305 18808
rect 211505 18288 213305 18544
rect 211505 18024 212643 18288
rect 212907 18024 213305 18288
rect 211505 17768 213305 18024
rect 211505 17504 212643 17768
rect 212907 17504 213305 17768
rect 211505 17248 213305 17504
rect 211505 16984 212643 17248
rect 212907 16984 213305 17248
rect 211505 16728 213305 16984
rect 211505 16464 212643 16728
rect 212907 16464 213305 16728
rect 211505 16208 213305 16464
rect 211505 15944 212643 16208
rect 212907 15944 213305 16208
rect 211505 15688 213305 15944
rect 211505 15424 212643 15688
rect 212907 15424 213305 15688
rect 211505 15168 213305 15424
rect 211505 14904 212643 15168
rect 212907 14904 213305 15168
rect 211505 14648 213305 14904
rect 211505 14384 212643 14648
rect 212907 14384 213305 14648
rect 211505 14128 213305 14384
rect 211505 13864 212643 14128
rect 212907 13864 213305 14128
rect 211505 13608 213305 13864
rect 211505 13344 212643 13608
rect 212907 13344 213305 13608
rect 211505 13088 213305 13344
rect 211505 12824 212643 13088
rect 212907 12824 213305 13088
rect 211505 12568 213305 12824
rect 211505 12304 212643 12568
rect 212907 12304 213305 12568
rect 211505 12048 213305 12304
rect 211505 11784 212643 12048
rect 212907 11784 213305 12048
rect 211505 11528 213305 11784
rect 211505 11264 212643 11528
rect 212907 11264 213305 11528
rect 211505 11008 213305 11264
rect 211505 10744 212643 11008
rect 212907 10744 213305 11008
rect 211505 10488 213305 10744
rect 211505 10224 212643 10488
rect 212907 10224 213305 10488
rect 211505 9968 213305 10224
rect 211505 9716 212643 9968
rect 185905 9704 212643 9716
rect 212907 9704 213305 9968
rect 185905 9116 213305 9704
rect 189236 8391 191843 9116
rect 189236 7938 189991 8391
rect 190976 7938 191843 8391
rect 189236 7379 191843 7938
rect 156625 5605 177825 6743
rect 156625 5341 157213 5605
rect 157477 5341 157733 5605
rect 157997 5341 158253 5605
rect 158517 5341 158773 5605
rect 159037 5341 159293 5605
rect 159557 5341 159813 5605
rect 160077 5341 160333 5605
rect 160597 5341 160853 5605
rect 161117 5341 161373 5605
rect 161637 5341 161893 5605
rect 162157 5341 162413 5605
rect 162677 5341 162933 5605
rect 163197 5341 163453 5605
rect 163717 5341 163973 5605
rect 164237 5341 164493 5605
rect 164757 5341 165013 5605
rect 165277 5341 165533 5605
rect 165797 5341 166053 5605
rect 166317 5341 166573 5605
rect 166837 5341 167093 5605
rect 167357 5341 167613 5605
rect 167877 5341 168133 5605
rect 168397 5341 168653 5605
rect 168917 5341 169173 5605
rect 169437 5341 169693 5605
rect 169957 5341 170213 5605
rect 170477 5341 170733 5605
rect 170997 5341 171253 5605
rect 171517 5341 171773 5605
rect 172037 5341 172293 5605
rect 172557 5341 172813 5605
rect 173077 5341 173333 5605
rect 173597 5341 173853 5605
rect 174117 5341 174373 5605
rect 174637 5341 174893 5605
rect 175157 5341 175413 5605
rect 175677 5341 175933 5605
rect 176197 5341 176453 5605
rect 176717 5341 176973 5605
rect 177237 5341 177825 5605
rect 156625 4943 177825 5341
rect 121546 4544 124153 4943
rect 121546 4091 122301 4544
rect 123286 4091 124153 4544
rect 121546 3532 124153 4091
<< via4 >>
rect 113613 5341 113877 5605
rect 114133 5341 114397 5605
rect 114653 5341 114917 5605
rect 115173 5341 115437 5605
rect 115693 5341 115957 5605
rect 116213 5341 116477 5605
rect 116733 5341 116997 5605
rect 117253 5341 117517 5605
rect 117773 5341 118037 5605
rect 118293 5341 118557 5605
rect 118813 5341 119077 5605
rect 119333 5341 119597 5605
rect 119853 5341 120117 5605
rect 120373 5341 120637 5605
rect 120893 5341 121157 5605
rect 121413 5341 121677 5605
rect 121933 5341 122197 5605
rect 122453 5341 122717 5605
rect 122973 5341 123237 5605
rect 123493 5341 123757 5605
rect 124013 5341 124277 5605
rect 124533 5341 124797 5605
rect 125053 5341 125317 5605
rect 125573 5341 125837 5605
rect 126093 5341 126357 5605
rect 126613 5341 126877 5605
rect 127133 5341 127397 5605
rect 127653 5341 127917 5605
rect 128173 5341 128437 5605
rect 128693 5341 128957 5605
rect 129213 5341 129477 5605
rect 129733 5341 129997 5605
rect 130253 5341 130517 5605
rect 130773 5341 131037 5605
rect 131293 5341 131557 5605
rect 131813 5341 132077 5605
rect 132333 5341 132597 5605
rect 132853 5341 133117 5605
rect 133373 5341 133637 5605
rect 135413 5341 135677 5605
rect 135933 5341 136197 5605
rect 136453 5341 136717 5605
rect 136973 5341 137237 5605
rect 137493 5341 137757 5605
rect 138013 5341 138277 5605
rect 138533 5341 138797 5605
rect 139053 5341 139317 5605
rect 139573 5341 139837 5605
rect 140093 5341 140357 5605
rect 140613 5341 140877 5605
rect 141133 5341 141397 5605
rect 141653 5341 141917 5605
rect 142173 5341 142437 5605
rect 142693 5341 142957 5605
rect 143213 5341 143477 5605
rect 143733 5341 143997 5605
rect 144253 5341 144517 5605
rect 144773 5341 145037 5605
rect 145293 5341 145557 5605
rect 145813 5341 146077 5605
rect 146333 5341 146597 5605
rect 146853 5341 147117 5605
rect 147373 5341 147637 5605
rect 147893 5341 148157 5605
rect 148413 5341 148677 5605
rect 148933 5341 149197 5605
rect 149453 5341 149717 5605
rect 149973 5341 150237 5605
rect 150493 5341 150757 5605
rect 151013 5341 151277 5605
rect 151533 5341 151797 5605
rect 152053 5341 152317 5605
rect 152573 5341 152837 5605
rect 153093 5341 153357 5605
rect 153613 5341 153877 5605
rect 154133 5341 154397 5605
rect 154653 5341 154917 5605
rect 155173 5341 155437 5605
rect 179090 18992 179707 19469
rect 212643 29464 212907 29728
rect 212643 28944 212907 29208
rect 212643 28424 212907 28688
rect 212643 27904 212907 28168
rect 212643 27384 212907 27648
rect 212643 26864 212907 27128
rect 212643 26344 212907 26608
rect 212643 25824 212907 26088
rect 212643 25304 212907 25568
rect 212643 24784 212907 25048
rect 212643 24264 212907 24528
rect 212643 23744 212907 24008
rect 212643 23224 212907 23488
rect 212643 22704 212907 22968
rect 212643 22184 212907 22448
rect 212643 21664 212907 21928
rect 212643 21144 212907 21408
rect 212643 20624 212907 20888
rect 212643 20104 212907 20368
rect 212643 19584 212907 19848
rect 212643 19064 212907 19328
rect 212643 18544 212907 18808
rect 212643 18024 212907 18288
rect 212643 17504 212907 17768
rect 212643 16984 212907 17248
rect 212643 16464 212907 16728
rect 212643 15944 212907 16208
rect 212643 15424 212907 15688
rect 212643 14904 212907 15168
rect 212643 14384 212907 14648
rect 212643 13864 212907 14128
rect 212643 13344 212907 13608
rect 212643 12824 212907 13088
rect 212643 12304 212907 12568
rect 212643 11784 212907 12048
rect 212643 11264 212907 11528
rect 212643 10744 212907 11008
rect 212643 10224 212907 10488
rect 212643 9704 212907 9968
rect 157213 5341 157477 5605
rect 157733 5341 157997 5605
rect 158253 5341 158517 5605
rect 158773 5341 159037 5605
rect 159293 5341 159557 5605
rect 159813 5341 160077 5605
rect 160333 5341 160597 5605
rect 160853 5341 161117 5605
rect 161373 5341 161637 5605
rect 161893 5341 162157 5605
rect 162413 5341 162677 5605
rect 162933 5341 163197 5605
rect 163453 5341 163717 5605
rect 163973 5341 164237 5605
rect 164493 5341 164757 5605
rect 165013 5341 165277 5605
rect 165533 5341 165797 5605
rect 166053 5341 166317 5605
rect 166573 5341 166837 5605
rect 167093 5341 167357 5605
rect 167613 5341 167877 5605
rect 168133 5341 168397 5605
rect 168653 5341 168917 5605
rect 169173 5341 169437 5605
rect 169693 5341 169957 5605
rect 170213 5341 170477 5605
rect 170733 5341 170997 5605
rect 171253 5341 171517 5605
rect 171773 5341 172037 5605
rect 172293 5341 172557 5605
rect 172813 5341 173077 5605
rect 173333 5341 173597 5605
rect 173853 5341 174117 5605
rect 174373 5341 174637 5605
rect 174893 5341 175157 5605
rect 175413 5341 175677 5605
rect 175933 5341 176197 5605
rect 176453 5341 176717 5605
rect 176973 5341 177237 5605
<< metal5 >>
rect 114025 31171 133225 31343
rect 114025 30875 114357 31171
rect 114653 30875 115117 31171
rect 115413 30875 115877 31171
rect 116173 30875 116637 31171
rect 116933 30875 117397 31171
rect 117693 30875 118157 31171
rect 118453 30875 118917 31171
rect 119213 30875 119677 31171
rect 119973 30875 120437 31171
rect 120733 30875 121197 31171
rect 121493 30875 121957 31171
rect 122253 30875 122717 31171
rect 123013 30875 123477 31171
rect 123773 30875 124237 31171
rect 124533 30875 124997 31171
rect 125293 30875 125757 31171
rect 126053 30875 126517 31171
rect 126813 30875 127277 31171
rect 127573 30875 128037 31171
rect 128333 30875 128797 31171
rect 129093 30875 129557 31171
rect 129853 30875 130317 31171
rect 130613 30875 131077 31171
rect 131373 30875 131837 31171
rect 132133 30875 132597 31171
rect 132893 30875 133225 31171
rect 114025 30411 133225 30875
rect 114025 30115 114357 30411
rect 114653 30115 115117 30411
rect 115413 30115 115877 30411
rect 116173 30115 116637 30411
rect 116933 30115 117397 30411
rect 117693 30115 118157 30411
rect 118453 30115 118917 30411
rect 119213 30115 119677 30411
rect 119973 30115 120437 30411
rect 120733 30115 121197 30411
rect 121493 30115 121957 30411
rect 122253 30115 122717 30411
rect 123013 30115 123477 30411
rect 123773 30115 124237 30411
rect 124533 30115 124997 30411
rect 125293 30115 125757 30411
rect 126053 30115 126517 30411
rect 126813 30115 127277 30411
rect 127573 30115 128037 30411
rect 128333 30115 128797 30411
rect 129093 30115 129557 30411
rect 129853 30115 130317 30411
rect 130613 30115 131077 30411
rect 131373 30115 131837 30411
rect 132133 30115 132597 30411
rect 132893 30115 133225 30411
rect 114025 29651 133225 30115
rect 114025 29355 114357 29651
rect 114653 29355 115117 29651
rect 115413 29355 115877 29651
rect 116173 29355 116637 29651
rect 116933 29355 117397 29651
rect 117693 29355 118157 29651
rect 118453 29355 118917 29651
rect 119213 29355 119677 29651
rect 119973 29355 120437 29651
rect 120733 29355 121197 29651
rect 121493 29355 121957 29651
rect 122253 29355 122717 29651
rect 123013 29355 123477 29651
rect 123773 29355 124237 29651
rect 124533 29355 124997 29651
rect 125293 29355 125757 29651
rect 126053 29355 126517 29651
rect 126813 29355 127277 29651
rect 127573 29355 128037 29651
rect 128333 29355 128797 29651
rect 129093 29355 129557 29651
rect 129853 29355 130317 29651
rect 130613 29355 131077 29651
rect 131373 29355 131837 29651
rect 132133 29355 132597 29651
rect 132893 29355 133225 29651
rect 114025 28891 133225 29355
rect 114025 28595 114357 28891
rect 114653 28595 115117 28891
rect 115413 28595 115877 28891
rect 116173 28595 116637 28891
rect 116933 28595 117397 28891
rect 117693 28595 118157 28891
rect 118453 28595 118917 28891
rect 119213 28595 119677 28891
rect 119973 28595 120437 28891
rect 120733 28595 121197 28891
rect 121493 28595 121957 28891
rect 122253 28595 122717 28891
rect 123013 28595 123477 28891
rect 123773 28595 124237 28891
rect 124533 28595 124997 28891
rect 125293 28595 125757 28891
rect 126053 28595 126517 28891
rect 126813 28595 127277 28891
rect 127573 28595 128037 28891
rect 128333 28595 128797 28891
rect 129093 28595 129557 28891
rect 129853 28595 130317 28891
rect 130613 28595 131077 28891
rect 131373 28595 131837 28891
rect 132133 28595 132597 28891
rect 132893 28595 133225 28891
rect 114025 28131 133225 28595
rect 114025 27835 114357 28131
rect 114653 27835 115117 28131
rect 115413 27835 115877 28131
rect 116173 27835 116637 28131
rect 116933 27835 117397 28131
rect 117693 27835 118157 28131
rect 118453 27835 118917 28131
rect 119213 27835 119677 28131
rect 119973 27835 120437 28131
rect 120733 27835 121197 28131
rect 121493 27835 121957 28131
rect 122253 27835 122717 28131
rect 123013 27835 123477 28131
rect 123773 27835 124237 28131
rect 124533 27835 124997 28131
rect 125293 27835 125757 28131
rect 126053 27835 126517 28131
rect 126813 27835 127277 28131
rect 127573 27835 128037 28131
rect 128333 27835 128797 28131
rect 129093 27835 129557 28131
rect 129853 27835 130317 28131
rect 130613 27835 131077 28131
rect 131373 27835 131837 28131
rect 132133 27835 132597 28131
rect 132893 27835 133225 28131
rect 114025 27371 133225 27835
rect 114025 27075 114357 27371
rect 114653 27075 115117 27371
rect 115413 27075 115877 27371
rect 116173 27075 116637 27371
rect 116933 27075 117397 27371
rect 117693 27075 118157 27371
rect 118453 27075 118917 27371
rect 119213 27075 119677 27371
rect 119973 27075 120437 27371
rect 120733 27075 121197 27371
rect 121493 27075 121957 27371
rect 122253 27075 122717 27371
rect 123013 27075 123477 27371
rect 123773 27075 124237 27371
rect 124533 27075 124997 27371
rect 125293 27075 125757 27371
rect 126053 27075 126517 27371
rect 126813 27075 127277 27371
rect 127573 27075 128037 27371
rect 128333 27075 128797 27371
rect 129093 27075 129557 27371
rect 129853 27075 130317 27371
rect 130613 27075 131077 27371
rect 131373 27075 131837 27371
rect 132133 27075 132597 27371
rect 132893 27075 133225 27371
rect 114025 26611 133225 27075
rect 114025 26315 114357 26611
rect 114653 26315 115117 26611
rect 115413 26315 115877 26611
rect 116173 26315 116637 26611
rect 116933 26315 117397 26611
rect 117693 26315 118157 26611
rect 118453 26315 118917 26611
rect 119213 26315 119677 26611
rect 119973 26315 120437 26611
rect 120733 26315 121197 26611
rect 121493 26315 121957 26611
rect 122253 26315 122717 26611
rect 123013 26315 123477 26611
rect 123773 26315 124237 26611
rect 124533 26315 124997 26611
rect 125293 26315 125757 26611
rect 126053 26315 126517 26611
rect 126813 26315 127277 26611
rect 127573 26315 128037 26611
rect 128333 26315 128797 26611
rect 129093 26315 129557 26611
rect 129853 26315 130317 26611
rect 130613 26315 131077 26611
rect 131373 26315 131837 26611
rect 132133 26315 132597 26611
rect 132893 26315 133225 26611
rect 114025 25851 133225 26315
rect 114025 25555 114357 25851
rect 114653 25555 115117 25851
rect 115413 25555 115877 25851
rect 116173 25555 116637 25851
rect 116933 25555 117397 25851
rect 117693 25555 118157 25851
rect 118453 25555 118917 25851
rect 119213 25555 119677 25851
rect 119973 25555 120437 25851
rect 120733 25555 121197 25851
rect 121493 25555 121957 25851
rect 122253 25555 122717 25851
rect 123013 25555 123477 25851
rect 123773 25555 124237 25851
rect 124533 25555 124997 25851
rect 125293 25555 125757 25851
rect 126053 25555 126517 25851
rect 126813 25555 127277 25851
rect 127573 25555 128037 25851
rect 128333 25555 128797 25851
rect 129093 25555 129557 25851
rect 129853 25555 130317 25851
rect 130613 25555 131077 25851
rect 131373 25555 131837 25851
rect 132133 25555 132597 25851
rect 132893 25555 133225 25851
rect 114025 25091 133225 25555
rect 114025 24795 114357 25091
rect 114653 24795 115117 25091
rect 115413 24795 115877 25091
rect 116173 24795 116637 25091
rect 116933 24795 117397 25091
rect 117693 24795 118157 25091
rect 118453 24795 118917 25091
rect 119213 24795 119677 25091
rect 119973 24795 120437 25091
rect 120733 24795 121197 25091
rect 121493 24795 121957 25091
rect 122253 24795 122717 25091
rect 123013 24795 123477 25091
rect 123773 24795 124237 25091
rect 124533 24795 124997 25091
rect 125293 24795 125757 25091
rect 126053 24795 126517 25091
rect 126813 24795 127277 25091
rect 127573 24795 128037 25091
rect 128333 24795 128797 25091
rect 129093 24795 129557 25091
rect 129853 24795 130317 25091
rect 130613 24795 131077 25091
rect 131373 24795 131837 25091
rect 132133 24795 132597 25091
rect 132893 24795 133225 25091
rect 114025 24331 133225 24795
rect 114025 24035 114357 24331
rect 114653 24035 115117 24331
rect 115413 24035 115877 24331
rect 116173 24035 116637 24331
rect 116933 24035 117397 24331
rect 117693 24035 118157 24331
rect 118453 24035 118917 24331
rect 119213 24035 119677 24331
rect 119973 24035 120437 24331
rect 120733 24035 121197 24331
rect 121493 24035 121957 24331
rect 122253 24035 122717 24331
rect 123013 24035 123477 24331
rect 123773 24035 124237 24331
rect 124533 24035 124997 24331
rect 125293 24035 125757 24331
rect 126053 24035 126517 24331
rect 126813 24035 127277 24331
rect 127573 24035 128037 24331
rect 128333 24035 128797 24331
rect 129093 24035 129557 24331
rect 129853 24035 130317 24331
rect 130613 24035 131077 24331
rect 131373 24035 131837 24331
rect 132133 24035 132597 24331
rect 132893 24035 133225 24331
rect 114025 23571 133225 24035
rect 114025 23275 114357 23571
rect 114653 23275 115117 23571
rect 115413 23275 115877 23571
rect 116173 23275 116637 23571
rect 116933 23275 117397 23571
rect 117693 23275 118157 23571
rect 118453 23275 118917 23571
rect 119213 23275 119677 23571
rect 119973 23275 120437 23571
rect 120733 23275 121197 23571
rect 121493 23275 121957 23571
rect 122253 23275 122717 23571
rect 123013 23275 123477 23571
rect 123773 23275 124237 23571
rect 124533 23275 124997 23571
rect 125293 23275 125757 23571
rect 126053 23275 126517 23571
rect 126813 23275 127277 23571
rect 127573 23275 128037 23571
rect 128333 23275 128797 23571
rect 129093 23275 129557 23571
rect 129853 23275 130317 23571
rect 130613 23275 131077 23571
rect 131373 23275 131837 23571
rect 132133 23275 132597 23571
rect 132893 23275 133225 23571
rect 114025 22811 133225 23275
rect 114025 22515 114357 22811
rect 114653 22515 115117 22811
rect 115413 22515 115877 22811
rect 116173 22515 116637 22811
rect 116933 22515 117397 22811
rect 117693 22515 118157 22811
rect 118453 22515 118917 22811
rect 119213 22515 119677 22811
rect 119973 22515 120437 22811
rect 120733 22515 121197 22811
rect 121493 22515 121957 22811
rect 122253 22515 122717 22811
rect 123013 22515 123477 22811
rect 123773 22515 124237 22811
rect 124533 22515 124997 22811
rect 125293 22515 125757 22811
rect 126053 22515 126517 22811
rect 126813 22515 127277 22811
rect 127573 22515 128037 22811
rect 128333 22515 128797 22811
rect 129093 22515 129557 22811
rect 129853 22515 130317 22811
rect 130613 22515 131077 22811
rect 131373 22515 131837 22811
rect 132133 22515 132597 22811
rect 132893 22515 133225 22811
rect 114025 22051 133225 22515
rect 114025 21755 114357 22051
rect 114653 21755 115117 22051
rect 115413 21755 115877 22051
rect 116173 21755 116637 22051
rect 116933 21755 117397 22051
rect 117693 21755 118157 22051
rect 118453 21755 118917 22051
rect 119213 21755 119677 22051
rect 119973 21755 120437 22051
rect 120733 21755 121197 22051
rect 121493 21755 121957 22051
rect 122253 21755 122717 22051
rect 123013 21755 123477 22051
rect 123773 21755 124237 22051
rect 124533 21755 124997 22051
rect 125293 21755 125757 22051
rect 126053 21755 126517 22051
rect 126813 21755 127277 22051
rect 127573 21755 128037 22051
rect 128333 21755 128797 22051
rect 129093 21755 129557 22051
rect 129853 21755 130317 22051
rect 130613 21755 131077 22051
rect 131373 21755 131837 22051
rect 132133 21755 132597 22051
rect 132893 21755 133225 22051
rect 114025 21291 133225 21755
rect 114025 20995 114357 21291
rect 114653 20995 115117 21291
rect 115413 20995 115877 21291
rect 116173 20995 116637 21291
rect 116933 20995 117397 21291
rect 117693 20995 118157 21291
rect 118453 20995 118917 21291
rect 119213 20995 119677 21291
rect 119973 20995 120437 21291
rect 120733 20995 121197 21291
rect 121493 20995 121957 21291
rect 122253 20995 122717 21291
rect 123013 20995 123477 21291
rect 123773 20995 124237 21291
rect 124533 20995 124997 21291
rect 125293 20995 125757 21291
rect 126053 20995 126517 21291
rect 126813 20995 127277 21291
rect 127573 20995 128037 21291
rect 128333 20995 128797 21291
rect 129093 20995 129557 21291
rect 129853 20995 130317 21291
rect 130613 20995 131077 21291
rect 131373 20995 131837 21291
rect 132133 20995 132597 21291
rect 132893 20995 133225 21291
rect 114025 20531 133225 20995
rect 114025 20235 114357 20531
rect 114653 20235 115117 20531
rect 115413 20235 115877 20531
rect 116173 20235 116637 20531
rect 116933 20235 117397 20531
rect 117693 20235 118157 20531
rect 118453 20235 118917 20531
rect 119213 20235 119677 20531
rect 119973 20235 120437 20531
rect 120733 20235 121197 20531
rect 121493 20235 121957 20531
rect 122253 20235 122717 20531
rect 123013 20235 123477 20531
rect 123773 20235 124237 20531
rect 124533 20235 124997 20531
rect 125293 20235 125757 20531
rect 126053 20235 126517 20531
rect 126813 20235 127277 20531
rect 127573 20235 128037 20531
rect 128333 20235 128797 20531
rect 129093 20235 129557 20531
rect 129853 20235 130317 20531
rect 130613 20235 131077 20531
rect 131373 20235 131837 20531
rect 132133 20235 132597 20531
rect 132893 20235 133225 20531
rect 114025 19773 133225 20235
rect 135825 31171 155025 31343
rect 135825 30875 136157 31171
rect 136453 30875 136917 31171
rect 137213 30875 137677 31171
rect 137973 30875 138437 31171
rect 138733 30875 139197 31171
rect 139493 30875 139957 31171
rect 140253 30875 140717 31171
rect 141013 30875 141477 31171
rect 141773 30875 142237 31171
rect 142533 30875 142997 31171
rect 143293 30875 143757 31171
rect 144053 30875 144517 31171
rect 144813 30875 145277 31171
rect 145573 30875 146037 31171
rect 146333 30875 146797 31171
rect 147093 30875 147557 31171
rect 147853 30875 148317 31171
rect 148613 30875 149077 31171
rect 149373 30875 149837 31171
rect 150133 30875 150597 31171
rect 150893 30875 151357 31171
rect 151653 30875 152117 31171
rect 152413 30875 152877 31171
rect 153173 30875 153637 31171
rect 153933 30875 154397 31171
rect 154693 30875 155025 31171
rect 135825 30411 155025 30875
rect 135825 30115 136157 30411
rect 136453 30115 136917 30411
rect 137213 30115 137677 30411
rect 137973 30115 138437 30411
rect 138733 30115 139197 30411
rect 139493 30115 139957 30411
rect 140253 30115 140717 30411
rect 141013 30115 141477 30411
rect 141773 30115 142237 30411
rect 142533 30115 142997 30411
rect 143293 30115 143757 30411
rect 144053 30115 144517 30411
rect 144813 30115 145277 30411
rect 145573 30115 146037 30411
rect 146333 30115 146797 30411
rect 147093 30115 147557 30411
rect 147853 30115 148317 30411
rect 148613 30115 149077 30411
rect 149373 30115 149837 30411
rect 150133 30115 150597 30411
rect 150893 30115 151357 30411
rect 151653 30115 152117 30411
rect 152413 30115 152877 30411
rect 153173 30115 153637 30411
rect 153933 30115 154397 30411
rect 154693 30115 155025 30411
rect 135825 29651 155025 30115
rect 135825 29355 136157 29651
rect 136453 29355 136917 29651
rect 137213 29355 137677 29651
rect 137973 29355 138437 29651
rect 138733 29355 139197 29651
rect 139493 29355 139957 29651
rect 140253 29355 140717 29651
rect 141013 29355 141477 29651
rect 141773 29355 142237 29651
rect 142533 29355 142997 29651
rect 143293 29355 143757 29651
rect 144053 29355 144517 29651
rect 144813 29355 145277 29651
rect 145573 29355 146037 29651
rect 146333 29355 146797 29651
rect 147093 29355 147557 29651
rect 147853 29355 148317 29651
rect 148613 29355 149077 29651
rect 149373 29355 149837 29651
rect 150133 29355 150597 29651
rect 150893 29355 151357 29651
rect 151653 29355 152117 29651
rect 152413 29355 152877 29651
rect 153173 29355 153637 29651
rect 153933 29355 154397 29651
rect 154693 29355 155025 29651
rect 135825 28891 155025 29355
rect 135825 28595 136157 28891
rect 136453 28595 136917 28891
rect 137213 28595 137677 28891
rect 137973 28595 138437 28891
rect 138733 28595 139197 28891
rect 139493 28595 139957 28891
rect 140253 28595 140717 28891
rect 141013 28595 141477 28891
rect 141773 28595 142237 28891
rect 142533 28595 142997 28891
rect 143293 28595 143757 28891
rect 144053 28595 144517 28891
rect 144813 28595 145277 28891
rect 145573 28595 146037 28891
rect 146333 28595 146797 28891
rect 147093 28595 147557 28891
rect 147853 28595 148317 28891
rect 148613 28595 149077 28891
rect 149373 28595 149837 28891
rect 150133 28595 150597 28891
rect 150893 28595 151357 28891
rect 151653 28595 152117 28891
rect 152413 28595 152877 28891
rect 153173 28595 153637 28891
rect 153933 28595 154397 28891
rect 154693 28595 155025 28891
rect 135825 28131 155025 28595
rect 135825 27835 136157 28131
rect 136453 27835 136917 28131
rect 137213 27835 137677 28131
rect 137973 27835 138437 28131
rect 138733 27835 139197 28131
rect 139493 27835 139957 28131
rect 140253 27835 140717 28131
rect 141013 27835 141477 28131
rect 141773 27835 142237 28131
rect 142533 27835 142997 28131
rect 143293 27835 143757 28131
rect 144053 27835 144517 28131
rect 144813 27835 145277 28131
rect 145573 27835 146037 28131
rect 146333 27835 146797 28131
rect 147093 27835 147557 28131
rect 147853 27835 148317 28131
rect 148613 27835 149077 28131
rect 149373 27835 149837 28131
rect 150133 27835 150597 28131
rect 150893 27835 151357 28131
rect 151653 27835 152117 28131
rect 152413 27835 152877 28131
rect 153173 27835 153637 28131
rect 153933 27835 154397 28131
rect 154693 27835 155025 28131
rect 135825 27371 155025 27835
rect 135825 27075 136157 27371
rect 136453 27075 136917 27371
rect 137213 27075 137677 27371
rect 137973 27075 138437 27371
rect 138733 27075 139197 27371
rect 139493 27075 139957 27371
rect 140253 27075 140717 27371
rect 141013 27075 141477 27371
rect 141773 27075 142237 27371
rect 142533 27075 142997 27371
rect 143293 27075 143757 27371
rect 144053 27075 144517 27371
rect 144813 27075 145277 27371
rect 145573 27075 146037 27371
rect 146333 27075 146797 27371
rect 147093 27075 147557 27371
rect 147853 27075 148317 27371
rect 148613 27075 149077 27371
rect 149373 27075 149837 27371
rect 150133 27075 150597 27371
rect 150893 27075 151357 27371
rect 151653 27075 152117 27371
rect 152413 27075 152877 27371
rect 153173 27075 153637 27371
rect 153933 27075 154397 27371
rect 154693 27075 155025 27371
rect 135825 26611 155025 27075
rect 135825 26315 136157 26611
rect 136453 26315 136917 26611
rect 137213 26315 137677 26611
rect 137973 26315 138437 26611
rect 138733 26315 139197 26611
rect 139493 26315 139957 26611
rect 140253 26315 140717 26611
rect 141013 26315 141477 26611
rect 141773 26315 142237 26611
rect 142533 26315 142997 26611
rect 143293 26315 143757 26611
rect 144053 26315 144517 26611
rect 144813 26315 145277 26611
rect 145573 26315 146037 26611
rect 146333 26315 146797 26611
rect 147093 26315 147557 26611
rect 147853 26315 148317 26611
rect 148613 26315 149077 26611
rect 149373 26315 149837 26611
rect 150133 26315 150597 26611
rect 150893 26315 151357 26611
rect 151653 26315 152117 26611
rect 152413 26315 152877 26611
rect 153173 26315 153637 26611
rect 153933 26315 154397 26611
rect 154693 26315 155025 26611
rect 135825 25851 155025 26315
rect 135825 25555 136157 25851
rect 136453 25555 136917 25851
rect 137213 25555 137677 25851
rect 137973 25555 138437 25851
rect 138733 25555 139197 25851
rect 139493 25555 139957 25851
rect 140253 25555 140717 25851
rect 141013 25555 141477 25851
rect 141773 25555 142237 25851
rect 142533 25555 142997 25851
rect 143293 25555 143757 25851
rect 144053 25555 144517 25851
rect 144813 25555 145277 25851
rect 145573 25555 146037 25851
rect 146333 25555 146797 25851
rect 147093 25555 147557 25851
rect 147853 25555 148317 25851
rect 148613 25555 149077 25851
rect 149373 25555 149837 25851
rect 150133 25555 150597 25851
rect 150893 25555 151357 25851
rect 151653 25555 152117 25851
rect 152413 25555 152877 25851
rect 153173 25555 153637 25851
rect 153933 25555 154397 25851
rect 154693 25555 155025 25851
rect 135825 25091 155025 25555
rect 135825 24795 136157 25091
rect 136453 24795 136917 25091
rect 137213 24795 137677 25091
rect 137973 24795 138437 25091
rect 138733 24795 139197 25091
rect 139493 24795 139957 25091
rect 140253 24795 140717 25091
rect 141013 24795 141477 25091
rect 141773 24795 142237 25091
rect 142533 24795 142997 25091
rect 143293 24795 143757 25091
rect 144053 24795 144517 25091
rect 144813 24795 145277 25091
rect 145573 24795 146037 25091
rect 146333 24795 146797 25091
rect 147093 24795 147557 25091
rect 147853 24795 148317 25091
rect 148613 24795 149077 25091
rect 149373 24795 149837 25091
rect 150133 24795 150597 25091
rect 150893 24795 151357 25091
rect 151653 24795 152117 25091
rect 152413 24795 152877 25091
rect 153173 24795 153637 25091
rect 153933 24795 154397 25091
rect 154693 24795 155025 25091
rect 135825 24331 155025 24795
rect 135825 24035 136157 24331
rect 136453 24035 136917 24331
rect 137213 24035 137677 24331
rect 137973 24035 138437 24331
rect 138733 24035 139197 24331
rect 139493 24035 139957 24331
rect 140253 24035 140717 24331
rect 141013 24035 141477 24331
rect 141773 24035 142237 24331
rect 142533 24035 142997 24331
rect 143293 24035 143757 24331
rect 144053 24035 144517 24331
rect 144813 24035 145277 24331
rect 145573 24035 146037 24331
rect 146333 24035 146797 24331
rect 147093 24035 147557 24331
rect 147853 24035 148317 24331
rect 148613 24035 149077 24331
rect 149373 24035 149837 24331
rect 150133 24035 150597 24331
rect 150893 24035 151357 24331
rect 151653 24035 152117 24331
rect 152413 24035 152877 24331
rect 153173 24035 153637 24331
rect 153933 24035 154397 24331
rect 154693 24035 155025 24331
rect 135825 23571 155025 24035
rect 135825 23275 136157 23571
rect 136453 23275 136917 23571
rect 137213 23275 137677 23571
rect 137973 23275 138437 23571
rect 138733 23275 139197 23571
rect 139493 23275 139957 23571
rect 140253 23275 140717 23571
rect 141013 23275 141477 23571
rect 141773 23275 142237 23571
rect 142533 23275 142997 23571
rect 143293 23275 143757 23571
rect 144053 23275 144517 23571
rect 144813 23275 145277 23571
rect 145573 23275 146037 23571
rect 146333 23275 146797 23571
rect 147093 23275 147557 23571
rect 147853 23275 148317 23571
rect 148613 23275 149077 23571
rect 149373 23275 149837 23571
rect 150133 23275 150597 23571
rect 150893 23275 151357 23571
rect 151653 23275 152117 23571
rect 152413 23275 152877 23571
rect 153173 23275 153637 23571
rect 153933 23275 154397 23571
rect 154693 23275 155025 23571
rect 135825 22811 155025 23275
rect 135825 22515 136157 22811
rect 136453 22515 136917 22811
rect 137213 22515 137677 22811
rect 137973 22515 138437 22811
rect 138733 22515 139197 22811
rect 139493 22515 139957 22811
rect 140253 22515 140717 22811
rect 141013 22515 141477 22811
rect 141773 22515 142237 22811
rect 142533 22515 142997 22811
rect 143293 22515 143757 22811
rect 144053 22515 144517 22811
rect 144813 22515 145277 22811
rect 145573 22515 146037 22811
rect 146333 22515 146797 22811
rect 147093 22515 147557 22811
rect 147853 22515 148317 22811
rect 148613 22515 149077 22811
rect 149373 22515 149837 22811
rect 150133 22515 150597 22811
rect 150893 22515 151357 22811
rect 151653 22515 152117 22811
rect 152413 22515 152877 22811
rect 153173 22515 153637 22811
rect 153933 22515 154397 22811
rect 154693 22515 155025 22811
rect 135825 22051 155025 22515
rect 135825 21755 136157 22051
rect 136453 21755 136917 22051
rect 137213 21755 137677 22051
rect 137973 21755 138437 22051
rect 138733 21755 139197 22051
rect 139493 21755 139957 22051
rect 140253 21755 140717 22051
rect 141013 21755 141477 22051
rect 141773 21755 142237 22051
rect 142533 21755 142997 22051
rect 143293 21755 143757 22051
rect 144053 21755 144517 22051
rect 144813 21755 145277 22051
rect 145573 21755 146037 22051
rect 146333 21755 146797 22051
rect 147093 21755 147557 22051
rect 147853 21755 148317 22051
rect 148613 21755 149077 22051
rect 149373 21755 149837 22051
rect 150133 21755 150597 22051
rect 150893 21755 151357 22051
rect 151653 21755 152117 22051
rect 152413 21755 152877 22051
rect 153173 21755 153637 22051
rect 153933 21755 154397 22051
rect 154693 21755 155025 22051
rect 135825 21291 155025 21755
rect 135825 20995 136157 21291
rect 136453 20995 136917 21291
rect 137213 20995 137677 21291
rect 137973 20995 138437 21291
rect 138733 20995 139197 21291
rect 139493 20995 139957 21291
rect 140253 20995 140717 21291
rect 141013 20995 141477 21291
rect 141773 20995 142237 21291
rect 142533 20995 142997 21291
rect 143293 20995 143757 21291
rect 144053 20995 144517 21291
rect 144813 20995 145277 21291
rect 145573 20995 146037 21291
rect 146333 20995 146797 21291
rect 147093 20995 147557 21291
rect 147853 20995 148317 21291
rect 148613 20995 149077 21291
rect 149373 20995 149837 21291
rect 150133 20995 150597 21291
rect 150893 20995 151357 21291
rect 151653 20995 152117 21291
rect 152413 20995 152877 21291
rect 153173 20995 153637 21291
rect 153933 20995 154397 21291
rect 154693 20995 155025 21291
rect 135825 20531 155025 20995
rect 135825 20235 136157 20531
rect 136453 20235 136917 20531
rect 137213 20235 137677 20531
rect 137973 20235 138437 20531
rect 138733 20235 139197 20531
rect 139493 20235 139957 20531
rect 140253 20235 140717 20531
rect 141013 20235 141477 20531
rect 141773 20235 142237 20531
rect 142533 20235 142997 20531
rect 143293 20235 143757 20531
rect 144053 20235 144517 20531
rect 144813 20235 145277 20531
rect 145573 20235 146037 20531
rect 146333 20235 146797 20531
rect 147093 20235 147557 20531
rect 147853 20235 148317 20531
rect 148613 20235 149077 20531
rect 149373 20235 149837 20531
rect 150133 20235 150597 20531
rect 150893 20235 151357 20531
rect 151653 20235 152117 20531
rect 152413 20235 152877 20531
rect 153173 20235 153637 20531
rect 153933 20235 154397 20531
rect 154693 20235 155025 20531
rect 135825 19773 155025 20235
rect 157625 31171 176825 31343
rect 157625 30875 157957 31171
rect 158253 30875 158717 31171
rect 159013 30875 159477 31171
rect 159773 30875 160237 31171
rect 160533 30875 160997 31171
rect 161293 30875 161757 31171
rect 162053 30875 162517 31171
rect 162813 30875 163277 31171
rect 163573 30875 164037 31171
rect 164333 30875 164797 31171
rect 165093 30875 165557 31171
rect 165853 30875 166317 31171
rect 166613 30875 167077 31171
rect 167373 30875 167837 31171
rect 168133 30875 168597 31171
rect 168893 30875 169357 31171
rect 169653 30875 170117 31171
rect 170413 30875 170877 31171
rect 171173 30875 171637 31171
rect 171933 30875 172397 31171
rect 172693 30875 173157 31171
rect 173453 30875 173917 31171
rect 174213 30875 174677 31171
rect 174973 30875 175437 31171
rect 175733 30875 176197 31171
rect 176493 30875 176825 31171
rect 157625 30411 176825 30875
rect 157625 30115 157957 30411
rect 158253 30115 158717 30411
rect 159013 30115 159477 30411
rect 159773 30115 160237 30411
rect 160533 30115 160997 30411
rect 161293 30115 161757 30411
rect 162053 30115 162517 30411
rect 162813 30115 163277 30411
rect 163573 30115 164037 30411
rect 164333 30115 164797 30411
rect 165093 30115 165557 30411
rect 165853 30115 166317 30411
rect 166613 30115 167077 30411
rect 167373 30115 167837 30411
rect 168133 30115 168597 30411
rect 168893 30115 169357 30411
rect 169653 30115 170117 30411
rect 170413 30115 170877 30411
rect 171173 30115 171637 30411
rect 171933 30115 172397 30411
rect 172693 30115 173157 30411
rect 173453 30115 173917 30411
rect 174213 30115 174677 30411
rect 174973 30115 175437 30411
rect 175733 30115 176197 30411
rect 176493 30115 176825 30411
rect 157625 29651 176825 30115
rect 157625 29355 157957 29651
rect 158253 29355 158717 29651
rect 159013 29355 159477 29651
rect 159773 29355 160237 29651
rect 160533 29355 160997 29651
rect 161293 29355 161757 29651
rect 162053 29355 162517 29651
rect 162813 29355 163277 29651
rect 163573 29355 164037 29651
rect 164333 29355 164797 29651
rect 165093 29355 165557 29651
rect 165853 29355 166317 29651
rect 166613 29355 167077 29651
rect 167373 29355 167837 29651
rect 168133 29355 168597 29651
rect 168893 29355 169357 29651
rect 169653 29355 170117 29651
rect 170413 29355 170877 29651
rect 171173 29355 171637 29651
rect 171933 29355 172397 29651
rect 172693 29355 173157 29651
rect 173453 29355 173917 29651
rect 174213 29355 174677 29651
rect 174973 29355 175437 29651
rect 175733 29355 176197 29651
rect 176493 29355 176825 29651
rect 157625 28891 176825 29355
rect 212555 29728 212995 30031
rect 212555 29464 212643 29728
rect 212907 29464 212995 29728
rect 157625 28595 157957 28891
rect 158253 28595 158717 28891
rect 159013 28595 159477 28891
rect 159773 28595 160237 28891
rect 160533 28595 160997 28891
rect 161293 28595 161757 28891
rect 162053 28595 162517 28891
rect 162813 28595 163277 28891
rect 163573 28595 164037 28891
rect 164333 28595 164797 28891
rect 165093 28595 165557 28891
rect 165853 28595 166317 28891
rect 166613 28595 167077 28891
rect 167373 28595 167837 28891
rect 168133 28595 168597 28891
rect 168893 28595 169357 28891
rect 169653 28595 170117 28891
rect 170413 28595 170877 28891
rect 171173 28595 171637 28891
rect 171933 28595 172397 28891
rect 172693 28595 173157 28891
rect 173453 28595 173917 28891
rect 174213 28595 174677 28891
rect 174973 28595 175437 28891
rect 175733 28595 176197 28891
rect 176493 28595 176825 28891
rect 157625 28131 176825 28595
rect 157625 27835 157957 28131
rect 158253 27835 158717 28131
rect 159013 27835 159477 28131
rect 159773 27835 160237 28131
rect 160533 27835 160997 28131
rect 161293 27835 161757 28131
rect 162053 27835 162517 28131
rect 162813 27835 163277 28131
rect 163573 27835 164037 28131
rect 164333 27835 164797 28131
rect 165093 27835 165557 28131
rect 165853 27835 166317 28131
rect 166613 27835 167077 28131
rect 167373 27835 167837 28131
rect 168133 27835 168597 28131
rect 168893 27835 169357 28131
rect 169653 27835 170117 28131
rect 170413 27835 170877 28131
rect 171173 27835 171637 28131
rect 171933 27835 172397 28131
rect 172693 27835 173157 28131
rect 173453 27835 173917 28131
rect 174213 27835 174677 28131
rect 174973 27835 175437 28131
rect 175733 27835 176197 28131
rect 176493 27835 176825 28131
rect 157625 27371 176825 27835
rect 157625 27075 157957 27371
rect 158253 27075 158717 27371
rect 159013 27075 159477 27371
rect 159773 27075 160237 27371
rect 160533 27075 160997 27371
rect 161293 27075 161757 27371
rect 162053 27075 162517 27371
rect 162813 27075 163277 27371
rect 163573 27075 164037 27371
rect 164333 27075 164797 27371
rect 165093 27075 165557 27371
rect 165853 27075 166317 27371
rect 166613 27075 167077 27371
rect 167373 27075 167837 27371
rect 168133 27075 168597 27371
rect 168893 27075 169357 27371
rect 169653 27075 170117 27371
rect 170413 27075 170877 27371
rect 171173 27075 171637 27371
rect 171933 27075 172397 27371
rect 172693 27075 173157 27371
rect 173453 27075 173917 27371
rect 174213 27075 174677 27371
rect 174973 27075 175437 27371
rect 175733 27075 176197 27371
rect 176493 27075 176825 27371
rect 157625 26611 176825 27075
rect 157625 26315 157957 26611
rect 158253 26315 158717 26611
rect 159013 26315 159477 26611
rect 159773 26315 160237 26611
rect 160533 26315 160997 26611
rect 161293 26315 161757 26611
rect 162053 26315 162517 26611
rect 162813 26315 163277 26611
rect 163573 26315 164037 26611
rect 164333 26315 164797 26611
rect 165093 26315 165557 26611
rect 165853 26315 166317 26611
rect 166613 26315 167077 26611
rect 167373 26315 167837 26611
rect 168133 26315 168597 26611
rect 168893 26315 169357 26611
rect 169653 26315 170117 26611
rect 170413 26315 170877 26611
rect 171173 26315 171637 26611
rect 171933 26315 172397 26611
rect 172693 26315 173157 26611
rect 173453 26315 173917 26611
rect 174213 26315 174677 26611
rect 174973 26315 175437 26611
rect 175733 26315 176197 26611
rect 176493 26315 176825 26611
rect 157625 25851 176825 26315
rect 157625 25555 157957 25851
rect 158253 25555 158717 25851
rect 159013 25555 159477 25851
rect 159773 25555 160237 25851
rect 160533 25555 160997 25851
rect 161293 25555 161757 25851
rect 162053 25555 162517 25851
rect 162813 25555 163277 25851
rect 163573 25555 164037 25851
rect 164333 25555 164797 25851
rect 165093 25555 165557 25851
rect 165853 25555 166317 25851
rect 166613 25555 167077 25851
rect 167373 25555 167837 25851
rect 168133 25555 168597 25851
rect 168893 25555 169357 25851
rect 169653 25555 170117 25851
rect 170413 25555 170877 25851
rect 171173 25555 171637 25851
rect 171933 25555 172397 25851
rect 172693 25555 173157 25851
rect 173453 25555 173917 25851
rect 174213 25555 174677 25851
rect 174973 25555 175437 25851
rect 175733 25555 176197 25851
rect 176493 25555 176825 25851
rect 157625 25091 176825 25555
rect 157625 24795 157957 25091
rect 158253 24795 158717 25091
rect 159013 24795 159477 25091
rect 159773 24795 160237 25091
rect 160533 24795 160997 25091
rect 161293 24795 161757 25091
rect 162053 24795 162517 25091
rect 162813 24795 163277 25091
rect 163573 24795 164037 25091
rect 164333 24795 164797 25091
rect 165093 24795 165557 25091
rect 165853 24795 166317 25091
rect 166613 24795 167077 25091
rect 167373 24795 167837 25091
rect 168133 24795 168597 25091
rect 168893 24795 169357 25091
rect 169653 24795 170117 25091
rect 170413 24795 170877 25091
rect 171173 24795 171637 25091
rect 171933 24795 172397 25091
rect 172693 24795 173157 25091
rect 173453 24795 173917 25091
rect 174213 24795 174677 25091
rect 174973 24795 175437 25091
rect 175733 24795 176197 25091
rect 176493 24795 176825 25091
rect 157625 24331 176825 24795
rect 157625 24035 157957 24331
rect 158253 24035 158717 24331
rect 159013 24035 159477 24331
rect 159773 24035 160237 24331
rect 160533 24035 160997 24331
rect 161293 24035 161757 24331
rect 162053 24035 162517 24331
rect 162813 24035 163277 24331
rect 163573 24035 164037 24331
rect 164333 24035 164797 24331
rect 165093 24035 165557 24331
rect 165853 24035 166317 24331
rect 166613 24035 167077 24331
rect 167373 24035 167837 24331
rect 168133 24035 168597 24331
rect 168893 24035 169357 24331
rect 169653 24035 170117 24331
rect 170413 24035 170877 24331
rect 171173 24035 171637 24331
rect 171933 24035 172397 24331
rect 172693 24035 173157 24331
rect 173453 24035 173917 24331
rect 174213 24035 174677 24331
rect 174973 24035 175437 24331
rect 175733 24035 176197 24331
rect 176493 24035 176825 24331
rect 157625 23571 176825 24035
rect 157625 23275 157957 23571
rect 158253 23275 158717 23571
rect 159013 23275 159477 23571
rect 159773 23275 160237 23571
rect 160533 23275 160997 23571
rect 161293 23275 161757 23571
rect 162053 23275 162517 23571
rect 162813 23275 163277 23571
rect 163573 23275 164037 23571
rect 164333 23275 164797 23571
rect 165093 23275 165557 23571
rect 165853 23275 166317 23571
rect 166613 23275 167077 23571
rect 167373 23275 167837 23571
rect 168133 23275 168597 23571
rect 168893 23275 169357 23571
rect 169653 23275 170117 23571
rect 170413 23275 170877 23571
rect 171173 23275 171637 23571
rect 171933 23275 172397 23571
rect 172693 23275 173157 23571
rect 173453 23275 173917 23571
rect 174213 23275 174677 23571
rect 174973 23275 175437 23571
rect 175733 23275 176197 23571
rect 176493 23275 176825 23571
rect 157625 22811 176825 23275
rect 157625 22515 157957 22811
rect 158253 22515 158717 22811
rect 159013 22515 159477 22811
rect 159773 22515 160237 22811
rect 160533 22515 160997 22811
rect 161293 22515 161757 22811
rect 162053 22515 162517 22811
rect 162813 22515 163277 22811
rect 163573 22515 164037 22811
rect 164333 22515 164797 22811
rect 165093 22515 165557 22811
rect 165853 22515 166317 22811
rect 166613 22515 167077 22811
rect 167373 22515 167837 22811
rect 168133 22515 168597 22811
rect 168893 22515 169357 22811
rect 169653 22515 170117 22811
rect 170413 22515 170877 22811
rect 171173 22515 171637 22811
rect 171933 22515 172397 22811
rect 172693 22515 173157 22811
rect 173453 22515 173917 22811
rect 174213 22515 174677 22811
rect 174973 22515 175437 22811
rect 175733 22515 176197 22811
rect 176493 22515 176825 22811
rect 157625 22051 176825 22515
rect 157625 21755 157957 22051
rect 158253 21755 158717 22051
rect 159013 21755 159477 22051
rect 159773 21755 160237 22051
rect 160533 21755 160997 22051
rect 161293 21755 161757 22051
rect 162053 21755 162517 22051
rect 162813 21755 163277 22051
rect 163573 21755 164037 22051
rect 164333 21755 164797 22051
rect 165093 21755 165557 22051
rect 165853 21755 166317 22051
rect 166613 21755 167077 22051
rect 167373 21755 167837 22051
rect 168133 21755 168597 22051
rect 168893 21755 169357 22051
rect 169653 21755 170117 22051
rect 170413 21755 170877 22051
rect 171173 21755 171637 22051
rect 171933 21755 172397 22051
rect 172693 21755 173157 22051
rect 173453 21755 173917 22051
rect 174213 21755 174677 22051
rect 174973 21755 175437 22051
rect 175733 21755 176197 22051
rect 176493 21755 176825 22051
rect 157625 21291 176825 21755
rect 157625 20995 157957 21291
rect 158253 20995 158717 21291
rect 159013 20995 159477 21291
rect 159773 20995 160237 21291
rect 160533 20995 160997 21291
rect 161293 20995 161757 21291
rect 162053 20995 162517 21291
rect 162813 20995 163277 21291
rect 163573 20995 164037 21291
rect 164333 20995 164797 21291
rect 165093 20995 165557 21291
rect 165853 20995 166317 21291
rect 166613 20995 167077 21291
rect 167373 20995 167837 21291
rect 168133 20995 168597 21291
rect 168893 20995 169357 21291
rect 169653 20995 170117 21291
rect 170413 20995 170877 21291
rect 171173 20995 171637 21291
rect 171933 20995 172397 21291
rect 172693 20995 173157 21291
rect 173453 20995 173917 21291
rect 174213 20995 174677 21291
rect 174973 20995 175437 21291
rect 175733 20995 176197 21291
rect 176493 20995 176825 21291
rect 157625 20531 176825 20995
rect 157625 20235 157957 20531
rect 158253 20235 158717 20531
rect 159013 20235 159477 20531
rect 159773 20235 160237 20531
rect 160533 20235 160997 20531
rect 161293 20235 161757 20531
rect 162053 20235 162517 20531
rect 162813 20235 163277 20531
rect 163573 20235 164037 20531
rect 164333 20235 164797 20531
rect 165093 20235 165557 20531
rect 165853 20235 166317 20531
rect 166613 20235 167077 20531
rect 167373 20235 167837 20531
rect 168133 20235 168597 20531
rect 168893 20235 169357 20531
rect 169653 20235 170117 20531
rect 170413 20235 170877 20531
rect 171173 20235 171637 20531
rect 171933 20235 172397 20531
rect 172693 20235 173157 20531
rect 173453 20235 173917 20531
rect 174213 20235 174677 20531
rect 174973 20235 175437 20531
rect 175733 20235 176197 20531
rect 176493 20235 176825 20531
rect 157625 19773 176825 20235
rect 186905 28984 211105 29316
rect 186905 28688 187077 28984
rect 187373 28688 187837 28984
rect 188133 28688 188597 28984
rect 188893 28688 189357 28984
rect 189653 28688 190117 28984
rect 190413 28688 190877 28984
rect 191173 28688 191637 28984
rect 191933 28688 192397 28984
rect 192693 28688 193157 28984
rect 193453 28688 193917 28984
rect 194213 28688 194677 28984
rect 194973 28688 195437 28984
rect 195733 28688 196197 28984
rect 196493 28688 196957 28984
rect 197253 28688 197717 28984
rect 198013 28688 198477 28984
rect 198773 28688 199237 28984
rect 199533 28688 199997 28984
rect 200293 28688 200757 28984
rect 201053 28688 201517 28984
rect 201813 28688 202277 28984
rect 202573 28688 203037 28984
rect 203333 28688 203797 28984
rect 204093 28688 204557 28984
rect 204853 28688 205317 28984
rect 205613 28688 206077 28984
rect 206373 28688 206837 28984
rect 207133 28688 207597 28984
rect 207893 28688 208357 28984
rect 208653 28688 209117 28984
rect 209413 28688 209877 28984
rect 210173 28688 210637 28984
rect 210933 28688 211105 28984
rect 186905 28224 211105 28688
rect 186905 27928 187077 28224
rect 187373 27928 187837 28224
rect 188133 27928 188597 28224
rect 188893 27928 189357 28224
rect 189653 27928 190117 28224
rect 190413 27928 190877 28224
rect 191173 27928 191637 28224
rect 191933 27928 192397 28224
rect 192693 27928 193157 28224
rect 193453 27928 193917 28224
rect 194213 27928 194677 28224
rect 194973 27928 195437 28224
rect 195733 27928 196197 28224
rect 196493 27928 196957 28224
rect 197253 27928 197717 28224
rect 198013 27928 198477 28224
rect 198773 27928 199237 28224
rect 199533 27928 199997 28224
rect 200293 27928 200757 28224
rect 201053 27928 201517 28224
rect 201813 27928 202277 28224
rect 202573 27928 203037 28224
rect 203333 27928 203797 28224
rect 204093 27928 204557 28224
rect 204853 27928 205317 28224
rect 205613 27928 206077 28224
rect 206373 27928 206837 28224
rect 207133 27928 207597 28224
rect 207893 27928 208357 28224
rect 208653 27928 209117 28224
rect 209413 27928 209877 28224
rect 210173 27928 210637 28224
rect 210933 27928 211105 28224
rect 186905 27464 211105 27928
rect 186905 27168 187077 27464
rect 187373 27168 187837 27464
rect 188133 27168 188597 27464
rect 188893 27168 189357 27464
rect 189653 27168 190117 27464
rect 190413 27168 190877 27464
rect 191173 27168 191637 27464
rect 191933 27168 192397 27464
rect 192693 27168 193157 27464
rect 193453 27168 193917 27464
rect 194213 27168 194677 27464
rect 194973 27168 195437 27464
rect 195733 27168 196197 27464
rect 196493 27168 196957 27464
rect 197253 27168 197717 27464
rect 198013 27168 198477 27464
rect 198773 27168 199237 27464
rect 199533 27168 199997 27464
rect 200293 27168 200757 27464
rect 201053 27168 201517 27464
rect 201813 27168 202277 27464
rect 202573 27168 203037 27464
rect 203333 27168 203797 27464
rect 204093 27168 204557 27464
rect 204853 27168 205317 27464
rect 205613 27168 206077 27464
rect 206373 27168 206837 27464
rect 207133 27168 207597 27464
rect 207893 27168 208357 27464
rect 208653 27168 209117 27464
rect 209413 27168 209877 27464
rect 210173 27168 210637 27464
rect 210933 27168 211105 27464
rect 186905 26704 211105 27168
rect 186905 26408 187077 26704
rect 187373 26408 187837 26704
rect 188133 26408 188597 26704
rect 188893 26408 189357 26704
rect 189653 26408 190117 26704
rect 190413 26408 190877 26704
rect 191173 26408 191637 26704
rect 191933 26408 192397 26704
rect 192693 26408 193157 26704
rect 193453 26408 193917 26704
rect 194213 26408 194677 26704
rect 194973 26408 195437 26704
rect 195733 26408 196197 26704
rect 196493 26408 196957 26704
rect 197253 26408 197717 26704
rect 198013 26408 198477 26704
rect 198773 26408 199237 26704
rect 199533 26408 199997 26704
rect 200293 26408 200757 26704
rect 201053 26408 201517 26704
rect 201813 26408 202277 26704
rect 202573 26408 203037 26704
rect 203333 26408 203797 26704
rect 204093 26408 204557 26704
rect 204853 26408 205317 26704
rect 205613 26408 206077 26704
rect 206373 26408 206837 26704
rect 207133 26408 207597 26704
rect 207893 26408 208357 26704
rect 208653 26408 209117 26704
rect 209413 26408 209877 26704
rect 210173 26408 210637 26704
rect 210933 26408 211105 26704
rect 186905 25944 211105 26408
rect 186905 25648 187077 25944
rect 187373 25648 187837 25944
rect 188133 25648 188597 25944
rect 188893 25648 189357 25944
rect 189653 25648 190117 25944
rect 190413 25648 190877 25944
rect 191173 25648 191637 25944
rect 191933 25648 192397 25944
rect 192693 25648 193157 25944
rect 193453 25648 193917 25944
rect 194213 25648 194677 25944
rect 194973 25648 195437 25944
rect 195733 25648 196197 25944
rect 196493 25648 196957 25944
rect 197253 25648 197717 25944
rect 198013 25648 198477 25944
rect 198773 25648 199237 25944
rect 199533 25648 199997 25944
rect 200293 25648 200757 25944
rect 201053 25648 201517 25944
rect 201813 25648 202277 25944
rect 202573 25648 203037 25944
rect 203333 25648 203797 25944
rect 204093 25648 204557 25944
rect 204853 25648 205317 25944
rect 205613 25648 206077 25944
rect 206373 25648 206837 25944
rect 207133 25648 207597 25944
rect 207893 25648 208357 25944
rect 208653 25648 209117 25944
rect 209413 25648 209877 25944
rect 210173 25648 210637 25944
rect 210933 25648 211105 25944
rect 186905 25184 211105 25648
rect 186905 24888 187077 25184
rect 187373 24888 187837 25184
rect 188133 24888 188597 25184
rect 188893 24888 189357 25184
rect 189653 24888 190117 25184
rect 190413 24888 190877 25184
rect 191173 24888 191637 25184
rect 191933 24888 192397 25184
rect 192693 24888 193157 25184
rect 193453 24888 193917 25184
rect 194213 24888 194677 25184
rect 194973 24888 195437 25184
rect 195733 24888 196197 25184
rect 196493 24888 196957 25184
rect 197253 24888 197717 25184
rect 198013 24888 198477 25184
rect 198773 24888 199237 25184
rect 199533 24888 199997 25184
rect 200293 24888 200757 25184
rect 201053 24888 201517 25184
rect 201813 24888 202277 25184
rect 202573 24888 203037 25184
rect 203333 24888 203797 25184
rect 204093 24888 204557 25184
rect 204853 24888 205317 25184
rect 205613 24888 206077 25184
rect 206373 24888 206837 25184
rect 207133 24888 207597 25184
rect 207893 24888 208357 25184
rect 208653 24888 209117 25184
rect 209413 24888 209877 25184
rect 210173 24888 210637 25184
rect 210933 24888 211105 25184
rect 186905 24424 211105 24888
rect 186905 24128 187077 24424
rect 187373 24128 187837 24424
rect 188133 24128 188597 24424
rect 188893 24128 189357 24424
rect 189653 24128 190117 24424
rect 190413 24128 190877 24424
rect 191173 24128 191637 24424
rect 191933 24128 192397 24424
rect 192693 24128 193157 24424
rect 193453 24128 193917 24424
rect 194213 24128 194677 24424
rect 194973 24128 195437 24424
rect 195733 24128 196197 24424
rect 196493 24128 196957 24424
rect 197253 24128 197717 24424
rect 198013 24128 198477 24424
rect 198773 24128 199237 24424
rect 199533 24128 199997 24424
rect 200293 24128 200757 24424
rect 201053 24128 201517 24424
rect 201813 24128 202277 24424
rect 202573 24128 203037 24424
rect 203333 24128 203797 24424
rect 204093 24128 204557 24424
rect 204853 24128 205317 24424
rect 205613 24128 206077 24424
rect 206373 24128 206837 24424
rect 207133 24128 207597 24424
rect 207893 24128 208357 24424
rect 208653 24128 209117 24424
rect 209413 24128 209877 24424
rect 210173 24128 210637 24424
rect 210933 24128 211105 24424
rect 186905 23664 211105 24128
rect 186905 23368 187077 23664
rect 187373 23368 187837 23664
rect 188133 23368 188597 23664
rect 188893 23368 189357 23664
rect 189653 23368 190117 23664
rect 190413 23368 190877 23664
rect 191173 23368 191637 23664
rect 191933 23368 192397 23664
rect 192693 23368 193157 23664
rect 193453 23368 193917 23664
rect 194213 23368 194677 23664
rect 194973 23368 195437 23664
rect 195733 23368 196197 23664
rect 196493 23368 196957 23664
rect 197253 23368 197717 23664
rect 198013 23368 198477 23664
rect 198773 23368 199237 23664
rect 199533 23368 199997 23664
rect 200293 23368 200757 23664
rect 201053 23368 201517 23664
rect 201813 23368 202277 23664
rect 202573 23368 203037 23664
rect 203333 23368 203797 23664
rect 204093 23368 204557 23664
rect 204853 23368 205317 23664
rect 205613 23368 206077 23664
rect 206373 23368 206837 23664
rect 207133 23368 207597 23664
rect 207893 23368 208357 23664
rect 208653 23368 209117 23664
rect 209413 23368 209877 23664
rect 210173 23368 210637 23664
rect 210933 23368 211105 23664
rect 186905 22904 211105 23368
rect 186905 22608 187077 22904
rect 187373 22608 187837 22904
rect 188133 22608 188597 22904
rect 188893 22608 189357 22904
rect 189653 22608 190117 22904
rect 190413 22608 190877 22904
rect 191173 22608 191637 22904
rect 191933 22608 192397 22904
rect 192693 22608 193157 22904
rect 193453 22608 193917 22904
rect 194213 22608 194677 22904
rect 194973 22608 195437 22904
rect 195733 22608 196197 22904
rect 196493 22608 196957 22904
rect 197253 22608 197717 22904
rect 198013 22608 198477 22904
rect 198773 22608 199237 22904
rect 199533 22608 199997 22904
rect 200293 22608 200757 22904
rect 201053 22608 201517 22904
rect 201813 22608 202277 22904
rect 202573 22608 203037 22904
rect 203333 22608 203797 22904
rect 204093 22608 204557 22904
rect 204853 22608 205317 22904
rect 205613 22608 206077 22904
rect 206373 22608 206837 22904
rect 207133 22608 207597 22904
rect 207893 22608 208357 22904
rect 208653 22608 209117 22904
rect 209413 22608 209877 22904
rect 210173 22608 210637 22904
rect 210933 22608 211105 22904
rect 186905 22144 211105 22608
rect 186905 21848 187077 22144
rect 187373 21848 187837 22144
rect 188133 21848 188597 22144
rect 188893 21848 189357 22144
rect 189653 21848 190117 22144
rect 190413 21848 190877 22144
rect 191173 21848 191637 22144
rect 191933 21848 192397 22144
rect 192693 21848 193157 22144
rect 193453 21848 193917 22144
rect 194213 21848 194677 22144
rect 194973 21848 195437 22144
rect 195733 21848 196197 22144
rect 196493 21848 196957 22144
rect 197253 21848 197717 22144
rect 198013 21848 198477 22144
rect 198773 21848 199237 22144
rect 199533 21848 199997 22144
rect 200293 21848 200757 22144
rect 201053 21848 201517 22144
rect 201813 21848 202277 22144
rect 202573 21848 203037 22144
rect 203333 21848 203797 22144
rect 204093 21848 204557 22144
rect 204853 21848 205317 22144
rect 205613 21848 206077 22144
rect 206373 21848 206837 22144
rect 207133 21848 207597 22144
rect 207893 21848 208357 22144
rect 208653 21848 209117 22144
rect 209413 21848 209877 22144
rect 210173 21848 210637 22144
rect 210933 21848 211105 22144
rect 186905 21384 211105 21848
rect 186905 21088 187077 21384
rect 187373 21088 187837 21384
rect 188133 21088 188597 21384
rect 188893 21088 189357 21384
rect 189653 21088 190117 21384
rect 190413 21088 190877 21384
rect 191173 21088 191637 21384
rect 191933 21088 192397 21384
rect 192693 21088 193157 21384
rect 193453 21088 193917 21384
rect 194213 21088 194677 21384
rect 194973 21088 195437 21384
rect 195733 21088 196197 21384
rect 196493 21088 196957 21384
rect 197253 21088 197717 21384
rect 198013 21088 198477 21384
rect 198773 21088 199237 21384
rect 199533 21088 199997 21384
rect 200293 21088 200757 21384
rect 201053 21088 201517 21384
rect 201813 21088 202277 21384
rect 202573 21088 203037 21384
rect 203333 21088 203797 21384
rect 204093 21088 204557 21384
rect 204853 21088 205317 21384
rect 205613 21088 206077 21384
rect 206373 21088 206837 21384
rect 207133 21088 207597 21384
rect 207893 21088 208357 21384
rect 208653 21088 209117 21384
rect 209413 21088 209877 21384
rect 210173 21088 210637 21384
rect 210933 21088 211105 21384
rect 186905 20624 211105 21088
rect 186905 20328 187077 20624
rect 187373 20328 187837 20624
rect 188133 20328 188597 20624
rect 188893 20328 189357 20624
rect 189653 20328 190117 20624
rect 190413 20328 190877 20624
rect 191173 20328 191637 20624
rect 191933 20328 192397 20624
rect 192693 20328 193157 20624
rect 193453 20328 193917 20624
rect 194213 20328 194677 20624
rect 194973 20328 195437 20624
rect 195733 20328 196197 20624
rect 196493 20328 196957 20624
rect 197253 20328 197717 20624
rect 198013 20328 198477 20624
rect 198773 20328 199237 20624
rect 199533 20328 199997 20624
rect 200293 20328 200757 20624
rect 201053 20328 201517 20624
rect 201813 20328 202277 20624
rect 202573 20328 203037 20624
rect 203333 20328 203797 20624
rect 204093 20328 204557 20624
rect 204853 20328 205317 20624
rect 205613 20328 206077 20624
rect 206373 20328 206837 20624
rect 207133 20328 207597 20624
rect 207893 20328 208357 20624
rect 208653 20328 209117 20624
rect 209413 20328 209877 20624
rect 210173 20328 210637 20624
rect 210933 20328 211105 20624
rect 186905 20028 211105 20328
rect 178058 19864 211105 20028
rect 178058 19773 187077 19864
rect 112725 19771 187077 19773
rect 112725 19475 114357 19771
rect 114653 19475 115117 19771
rect 115413 19475 115877 19771
rect 116173 19475 116637 19771
rect 116933 19475 117397 19771
rect 117693 19475 118157 19771
rect 118453 19475 118917 19771
rect 119213 19475 119677 19771
rect 119973 19475 120437 19771
rect 120733 19475 121197 19771
rect 121493 19475 121957 19771
rect 122253 19475 122717 19771
rect 123013 19475 123477 19771
rect 123773 19475 124237 19771
rect 124533 19475 124997 19771
rect 125293 19475 125757 19771
rect 126053 19475 126517 19771
rect 126813 19475 127277 19771
rect 127573 19475 128037 19771
rect 128333 19475 128797 19771
rect 129093 19475 129557 19771
rect 129853 19475 130317 19771
rect 130613 19475 131077 19771
rect 131373 19475 131837 19771
rect 132133 19475 132597 19771
rect 132893 19475 136157 19771
rect 136453 19475 136917 19771
rect 137213 19475 137677 19771
rect 137973 19475 138437 19771
rect 138733 19475 139197 19771
rect 139493 19475 139957 19771
rect 140253 19475 140717 19771
rect 141013 19475 141477 19771
rect 141773 19475 142237 19771
rect 142533 19475 142997 19771
rect 143293 19475 143757 19771
rect 144053 19475 144517 19771
rect 144813 19475 145277 19771
rect 145573 19475 146037 19771
rect 146333 19475 146797 19771
rect 147093 19475 147557 19771
rect 147853 19475 148317 19771
rect 148613 19475 149077 19771
rect 149373 19475 149837 19771
rect 150133 19475 150597 19771
rect 150893 19475 151357 19771
rect 151653 19475 152117 19771
rect 152413 19475 152877 19771
rect 153173 19475 153637 19771
rect 153933 19475 154397 19771
rect 154693 19475 157957 19771
rect 158253 19475 158717 19771
rect 159013 19475 159477 19771
rect 159773 19475 160237 19771
rect 160533 19475 160997 19771
rect 161293 19475 161757 19771
rect 162053 19475 162517 19771
rect 162813 19475 163277 19771
rect 163573 19475 164037 19771
rect 164333 19475 164797 19771
rect 165093 19475 165557 19771
rect 165853 19475 166317 19771
rect 166613 19475 167077 19771
rect 167373 19475 167837 19771
rect 168133 19475 168597 19771
rect 168893 19475 169357 19771
rect 169653 19475 170117 19771
rect 170413 19475 170877 19771
rect 171173 19475 171637 19771
rect 171933 19475 172397 19771
rect 172693 19475 173157 19771
rect 173453 19475 173917 19771
rect 174213 19475 174677 19771
rect 174973 19475 175437 19771
rect 175733 19475 176197 19771
rect 176493 19568 187077 19771
rect 187373 19568 187837 19864
rect 188133 19568 188597 19864
rect 188893 19568 189357 19864
rect 189653 19568 190117 19864
rect 190413 19568 190877 19864
rect 191173 19568 191637 19864
rect 191933 19568 192397 19864
rect 192693 19568 193157 19864
rect 193453 19568 193917 19864
rect 194213 19568 194677 19864
rect 194973 19568 195437 19864
rect 195733 19568 196197 19864
rect 196493 19568 196957 19864
rect 197253 19568 197717 19864
rect 198013 19568 198477 19864
rect 198773 19568 199237 19864
rect 199533 19568 199997 19864
rect 200293 19568 200757 19864
rect 201053 19568 201517 19864
rect 201813 19568 202277 19864
rect 202573 19568 203037 19864
rect 203333 19568 203797 19864
rect 204093 19568 204557 19864
rect 204853 19568 205317 19864
rect 205613 19568 206077 19864
rect 206373 19568 206837 19864
rect 207133 19568 207597 19864
rect 207893 19568 208357 19864
rect 208653 19568 209117 19864
rect 209413 19568 209877 19864
rect 210173 19568 210637 19864
rect 210933 19568 211105 19864
rect 176493 19475 211105 19568
rect 112725 19469 211105 19475
rect 112725 19011 179090 19469
rect 112725 18715 114357 19011
rect 114653 18715 115117 19011
rect 115413 18715 115877 19011
rect 116173 18715 116637 19011
rect 116933 18715 117397 19011
rect 117693 18715 118157 19011
rect 118453 18715 118917 19011
rect 119213 18715 119677 19011
rect 119973 18715 120437 19011
rect 120733 18715 121197 19011
rect 121493 18715 121957 19011
rect 122253 18715 122717 19011
rect 123013 18715 123477 19011
rect 123773 18715 124237 19011
rect 124533 18715 124997 19011
rect 125293 18715 125757 19011
rect 126053 18715 126517 19011
rect 126813 18715 127277 19011
rect 127573 18715 128037 19011
rect 128333 18715 128797 19011
rect 129093 18715 129557 19011
rect 129853 18715 130317 19011
rect 130613 18715 131077 19011
rect 131373 18715 131837 19011
rect 132133 18715 132597 19011
rect 132893 18715 136157 19011
rect 136453 18715 136917 19011
rect 137213 18715 137677 19011
rect 137973 18715 138437 19011
rect 138733 18715 139197 19011
rect 139493 18715 139957 19011
rect 140253 18715 140717 19011
rect 141013 18715 141477 19011
rect 141773 18715 142237 19011
rect 142533 18715 142997 19011
rect 143293 18715 143757 19011
rect 144053 18715 144517 19011
rect 144813 18715 145277 19011
rect 145573 18715 146037 19011
rect 146333 18715 146797 19011
rect 147093 18715 147557 19011
rect 147853 18715 148317 19011
rect 148613 18715 149077 19011
rect 149373 18715 149837 19011
rect 150133 18715 150597 19011
rect 150893 18715 151357 19011
rect 151653 18715 152117 19011
rect 152413 18715 152877 19011
rect 153173 18715 153637 19011
rect 153933 18715 154397 19011
rect 154693 18715 157957 19011
rect 158253 18715 158717 19011
rect 159013 18715 159477 19011
rect 159773 18715 160237 19011
rect 160533 18715 160997 19011
rect 161293 18715 161757 19011
rect 162053 18715 162517 19011
rect 162813 18715 163277 19011
rect 163573 18715 164037 19011
rect 164333 18715 164797 19011
rect 165093 18715 165557 19011
rect 165853 18715 166317 19011
rect 166613 18715 167077 19011
rect 167373 18715 167837 19011
rect 168133 18715 168597 19011
rect 168893 18715 169357 19011
rect 169653 18715 170117 19011
rect 170413 18715 170877 19011
rect 171173 18715 171637 19011
rect 171933 18715 172397 19011
rect 172693 18715 173157 19011
rect 173453 18715 173917 19011
rect 174213 18715 174677 19011
rect 174973 18715 175437 19011
rect 175733 18715 176197 19011
rect 176493 18992 179090 19011
rect 179707 19104 211105 19469
rect 179707 18992 187077 19104
rect 176493 18808 187077 18992
rect 187373 18808 187837 19104
rect 188133 18808 188597 19104
rect 188893 18808 189357 19104
rect 189653 18808 190117 19104
rect 190413 18808 190877 19104
rect 191173 18808 191637 19104
rect 191933 18808 192397 19104
rect 192693 18808 193157 19104
rect 193453 18808 193917 19104
rect 194213 18808 194677 19104
rect 194973 18808 195437 19104
rect 195733 18808 196197 19104
rect 196493 18808 196957 19104
rect 197253 18808 197717 19104
rect 198013 18808 198477 19104
rect 198773 18808 199237 19104
rect 199533 18808 199997 19104
rect 200293 18808 200757 19104
rect 201053 18808 201517 19104
rect 201813 18808 202277 19104
rect 202573 18808 203037 19104
rect 203333 18808 203797 19104
rect 204093 18808 204557 19104
rect 204853 18808 205317 19104
rect 205613 18808 206077 19104
rect 206373 18808 206837 19104
rect 207133 18808 207597 19104
rect 207893 18808 208357 19104
rect 208653 18808 209117 19104
rect 209413 18808 209877 19104
rect 210173 18808 210637 19104
rect 210933 18808 211105 19104
rect 176493 18715 211105 18808
rect 112725 18713 211105 18715
rect 114025 18251 133225 18713
rect 114025 17955 114357 18251
rect 114653 17955 115117 18251
rect 115413 17955 115877 18251
rect 116173 17955 116637 18251
rect 116933 17955 117397 18251
rect 117693 17955 118157 18251
rect 118453 17955 118917 18251
rect 119213 17955 119677 18251
rect 119973 17955 120437 18251
rect 120733 17955 121197 18251
rect 121493 17955 121957 18251
rect 122253 17955 122717 18251
rect 123013 17955 123477 18251
rect 123773 17955 124237 18251
rect 124533 17955 124997 18251
rect 125293 17955 125757 18251
rect 126053 17955 126517 18251
rect 126813 17955 127277 18251
rect 127573 17955 128037 18251
rect 128333 17955 128797 18251
rect 129093 17955 129557 18251
rect 129853 17955 130317 18251
rect 130613 17955 131077 18251
rect 131373 17955 131837 18251
rect 132133 17955 132597 18251
rect 132893 17955 133225 18251
rect 114025 17491 133225 17955
rect 114025 17195 114357 17491
rect 114653 17195 115117 17491
rect 115413 17195 115877 17491
rect 116173 17195 116637 17491
rect 116933 17195 117397 17491
rect 117693 17195 118157 17491
rect 118453 17195 118917 17491
rect 119213 17195 119677 17491
rect 119973 17195 120437 17491
rect 120733 17195 121197 17491
rect 121493 17195 121957 17491
rect 122253 17195 122717 17491
rect 123013 17195 123477 17491
rect 123773 17195 124237 17491
rect 124533 17195 124997 17491
rect 125293 17195 125757 17491
rect 126053 17195 126517 17491
rect 126813 17195 127277 17491
rect 127573 17195 128037 17491
rect 128333 17195 128797 17491
rect 129093 17195 129557 17491
rect 129853 17195 130317 17491
rect 130613 17195 131077 17491
rect 131373 17195 131837 17491
rect 132133 17195 132597 17491
rect 132893 17195 133225 17491
rect 114025 16731 133225 17195
rect 114025 16435 114357 16731
rect 114653 16435 115117 16731
rect 115413 16435 115877 16731
rect 116173 16435 116637 16731
rect 116933 16435 117397 16731
rect 117693 16435 118157 16731
rect 118453 16435 118917 16731
rect 119213 16435 119677 16731
rect 119973 16435 120437 16731
rect 120733 16435 121197 16731
rect 121493 16435 121957 16731
rect 122253 16435 122717 16731
rect 123013 16435 123477 16731
rect 123773 16435 124237 16731
rect 124533 16435 124997 16731
rect 125293 16435 125757 16731
rect 126053 16435 126517 16731
rect 126813 16435 127277 16731
rect 127573 16435 128037 16731
rect 128333 16435 128797 16731
rect 129093 16435 129557 16731
rect 129853 16435 130317 16731
rect 130613 16435 131077 16731
rect 131373 16435 131837 16731
rect 132133 16435 132597 16731
rect 132893 16435 133225 16731
rect 114025 15971 133225 16435
rect 114025 15675 114357 15971
rect 114653 15675 115117 15971
rect 115413 15675 115877 15971
rect 116173 15675 116637 15971
rect 116933 15675 117397 15971
rect 117693 15675 118157 15971
rect 118453 15675 118917 15971
rect 119213 15675 119677 15971
rect 119973 15675 120437 15971
rect 120733 15675 121197 15971
rect 121493 15675 121957 15971
rect 122253 15675 122717 15971
rect 123013 15675 123477 15971
rect 123773 15675 124237 15971
rect 124533 15675 124997 15971
rect 125293 15675 125757 15971
rect 126053 15675 126517 15971
rect 126813 15675 127277 15971
rect 127573 15675 128037 15971
rect 128333 15675 128797 15971
rect 129093 15675 129557 15971
rect 129853 15675 130317 15971
rect 130613 15675 131077 15971
rect 131373 15675 131837 15971
rect 132133 15675 132597 15971
rect 132893 15675 133225 15971
rect 114025 15211 133225 15675
rect 114025 14915 114357 15211
rect 114653 14915 115117 15211
rect 115413 14915 115877 15211
rect 116173 14915 116637 15211
rect 116933 14915 117397 15211
rect 117693 14915 118157 15211
rect 118453 14915 118917 15211
rect 119213 14915 119677 15211
rect 119973 14915 120437 15211
rect 120733 14915 121197 15211
rect 121493 14915 121957 15211
rect 122253 14915 122717 15211
rect 123013 14915 123477 15211
rect 123773 14915 124237 15211
rect 124533 14915 124997 15211
rect 125293 14915 125757 15211
rect 126053 14915 126517 15211
rect 126813 14915 127277 15211
rect 127573 14915 128037 15211
rect 128333 14915 128797 15211
rect 129093 14915 129557 15211
rect 129853 14915 130317 15211
rect 130613 14915 131077 15211
rect 131373 14915 131837 15211
rect 132133 14915 132597 15211
rect 132893 14915 133225 15211
rect 114025 14451 133225 14915
rect 114025 14155 114357 14451
rect 114653 14155 115117 14451
rect 115413 14155 115877 14451
rect 116173 14155 116637 14451
rect 116933 14155 117397 14451
rect 117693 14155 118157 14451
rect 118453 14155 118917 14451
rect 119213 14155 119677 14451
rect 119973 14155 120437 14451
rect 120733 14155 121197 14451
rect 121493 14155 121957 14451
rect 122253 14155 122717 14451
rect 123013 14155 123477 14451
rect 123773 14155 124237 14451
rect 124533 14155 124997 14451
rect 125293 14155 125757 14451
rect 126053 14155 126517 14451
rect 126813 14155 127277 14451
rect 127573 14155 128037 14451
rect 128333 14155 128797 14451
rect 129093 14155 129557 14451
rect 129853 14155 130317 14451
rect 130613 14155 131077 14451
rect 131373 14155 131837 14451
rect 132133 14155 132597 14451
rect 132893 14155 133225 14451
rect 114025 13691 133225 14155
rect 114025 13395 114357 13691
rect 114653 13395 115117 13691
rect 115413 13395 115877 13691
rect 116173 13395 116637 13691
rect 116933 13395 117397 13691
rect 117693 13395 118157 13691
rect 118453 13395 118917 13691
rect 119213 13395 119677 13691
rect 119973 13395 120437 13691
rect 120733 13395 121197 13691
rect 121493 13395 121957 13691
rect 122253 13395 122717 13691
rect 123013 13395 123477 13691
rect 123773 13395 124237 13691
rect 124533 13395 124997 13691
rect 125293 13395 125757 13691
rect 126053 13395 126517 13691
rect 126813 13395 127277 13691
rect 127573 13395 128037 13691
rect 128333 13395 128797 13691
rect 129093 13395 129557 13691
rect 129853 13395 130317 13691
rect 130613 13395 131077 13691
rect 131373 13395 131837 13691
rect 132133 13395 132597 13691
rect 132893 13395 133225 13691
rect 114025 12931 133225 13395
rect 114025 12635 114357 12931
rect 114653 12635 115117 12931
rect 115413 12635 115877 12931
rect 116173 12635 116637 12931
rect 116933 12635 117397 12931
rect 117693 12635 118157 12931
rect 118453 12635 118917 12931
rect 119213 12635 119677 12931
rect 119973 12635 120437 12931
rect 120733 12635 121197 12931
rect 121493 12635 121957 12931
rect 122253 12635 122717 12931
rect 123013 12635 123477 12931
rect 123773 12635 124237 12931
rect 124533 12635 124997 12931
rect 125293 12635 125757 12931
rect 126053 12635 126517 12931
rect 126813 12635 127277 12931
rect 127573 12635 128037 12931
rect 128333 12635 128797 12931
rect 129093 12635 129557 12931
rect 129853 12635 130317 12931
rect 130613 12635 131077 12931
rect 131373 12635 131837 12931
rect 132133 12635 132597 12931
rect 132893 12635 133225 12931
rect 114025 12171 133225 12635
rect 114025 11875 114357 12171
rect 114653 11875 115117 12171
rect 115413 11875 115877 12171
rect 116173 11875 116637 12171
rect 116933 11875 117397 12171
rect 117693 11875 118157 12171
rect 118453 11875 118917 12171
rect 119213 11875 119677 12171
rect 119973 11875 120437 12171
rect 120733 11875 121197 12171
rect 121493 11875 121957 12171
rect 122253 11875 122717 12171
rect 123013 11875 123477 12171
rect 123773 11875 124237 12171
rect 124533 11875 124997 12171
rect 125293 11875 125757 12171
rect 126053 11875 126517 12171
rect 126813 11875 127277 12171
rect 127573 11875 128037 12171
rect 128333 11875 128797 12171
rect 129093 11875 129557 12171
rect 129853 11875 130317 12171
rect 130613 11875 131077 12171
rect 131373 11875 131837 12171
rect 132133 11875 132597 12171
rect 132893 11875 133225 12171
rect 114025 11411 133225 11875
rect 114025 11115 114357 11411
rect 114653 11115 115117 11411
rect 115413 11115 115877 11411
rect 116173 11115 116637 11411
rect 116933 11115 117397 11411
rect 117693 11115 118157 11411
rect 118453 11115 118917 11411
rect 119213 11115 119677 11411
rect 119973 11115 120437 11411
rect 120733 11115 121197 11411
rect 121493 11115 121957 11411
rect 122253 11115 122717 11411
rect 123013 11115 123477 11411
rect 123773 11115 124237 11411
rect 124533 11115 124997 11411
rect 125293 11115 125757 11411
rect 126053 11115 126517 11411
rect 126813 11115 127277 11411
rect 127573 11115 128037 11411
rect 128333 11115 128797 11411
rect 129093 11115 129557 11411
rect 129853 11115 130317 11411
rect 130613 11115 131077 11411
rect 131373 11115 131837 11411
rect 132133 11115 132597 11411
rect 132893 11115 133225 11411
rect 114025 10651 133225 11115
rect 114025 10355 114357 10651
rect 114653 10355 115117 10651
rect 115413 10355 115877 10651
rect 116173 10355 116637 10651
rect 116933 10355 117397 10651
rect 117693 10355 118157 10651
rect 118453 10355 118917 10651
rect 119213 10355 119677 10651
rect 119973 10355 120437 10651
rect 120733 10355 121197 10651
rect 121493 10355 121957 10651
rect 122253 10355 122717 10651
rect 123013 10355 123477 10651
rect 123773 10355 124237 10651
rect 124533 10355 124997 10651
rect 125293 10355 125757 10651
rect 126053 10355 126517 10651
rect 126813 10355 127277 10651
rect 127573 10355 128037 10651
rect 128333 10355 128797 10651
rect 129093 10355 129557 10651
rect 129853 10355 130317 10651
rect 130613 10355 131077 10651
rect 131373 10355 131837 10651
rect 132133 10355 132597 10651
rect 132893 10355 133225 10651
rect 114025 9891 133225 10355
rect 114025 9595 114357 9891
rect 114653 9595 115117 9891
rect 115413 9595 115877 9891
rect 116173 9595 116637 9891
rect 116933 9595 117397 9891
rect 117693 9595 118157 9891
rect 118453 9595 118917 9891
rect 119213 9595 119677 9891
rect 119973 9595 120437 9891
rect 120733 9595 121197 9891
rect 121493 9595 121957 9891
rect 122253 9595 122717 9891
rect 123013 9595 123477 9891
rect 123773 9595 124237 9891
rect 124533 9595 124997 9891
rect 125293 9595 125757 9891
rect 126053 9595 126517 9891
rect 126813 9595 127277 9891
rect 127573 9595 128037 9891
rect 128333 9595 128797 9891
rect 129093 9595 129557 9891
rect 129853 9595 130317 9891
rect 130613 9595 131077 9891
rect 131373 9595 131837 9891
rect 132133 9595 132597 9891
rect 132893 9595 133225 9891
rect 114025 9131 133225 9595
rect 114025 8835 114357 9131
rect 114653 8835 115117 9131
rect 115413 8835 115877 9131
rect 116173 8835 116637 9131
rect 116933 8835 117397 9131
rect 117693 8835 118157 9131
rect 118453 8835 118917 9131
rect 119213 8835 119677 9131
rect 119973 8835 120437 9131
rect 120733 8835 121197 9131
rect 121493 8835 121957 9131
rect 122253 8835 122717 9131
rect 123013 8835 123477 9131
rect 123773 8835 124237 9131
rect 124533 8835 124997 9131
rect 125293 8835 125757 9131
rect 126053 8835 126517 9131
rect 126813 8835 127277 9131
rect 127573 8835 128037 9131
rect 128333 8835 128797 9131
rect 129093 8835 129557 9131
rect 129853 8835 130317 9131
rect 130613 8835 131077 9131
rect 131373 8835 131837 9131
rect 132133 8835 132597 9131
rect 132893 8835 133225 9131
rect 114025 8371 133225 8835
rect 114025 8075 114357 8371
rect 114653 8075 115117 8371
rect 115413 8075 115877 8371
rect 116173 8075 116637 8371
rect 116933 8075 117397 8371
rect 117693 8075 118157 8371
rect 118453 8075 118917 8371
rect 119213 8075 119677 8371
rect 119973 8075 120437 8371
rect 120733 8075 121197 8371
rect 121493 8075 121957 8371
rect 122253 8075 122717 8371
rect 123013 8075 123477 8371
rect 123773 8075 124237 8371
rect 124533 8075 124997 8371
rect 125293 8075 125757 8371
rect 126053 8075 126517 8371
rect 126813 8075 127277 8371
rect 127573 8075 128037 8371
rect 128333 8075 128797 8371
rect 129093 8075 129557 8371
rect 129853 8075 130317 8371
rect 130613 8075 131077 8371
rect 131373 8075 131837 8371
rect 132133 8075 132597 8371
rect 132893 8075 133225 8371
rect 114025 7611 133225 8075
rect 114025 7315 114357 7611
rect 114653 7315 115117 7611
rect 115413 7315 115877 7611
rect 116173 7315 116637 7611
rect 116933 7315 117397 7611
rect 117693 7315 118157 7611
rect 118453 7315 118917 7611
rect 119213 7315 119677 7611
rect 119973 7315 120437 7611
rect 120733 7315 121197 7611
rect 121493 7315 121957 7611
rect 122253 7315 122717 7611
rect 123013 7315 123477 7611
rect 123773 7315 124237 7611
rect 124533 7315 124997 7611
rect 125293 7315 125757 7611
rect 126053 7315 126517 7611
rect 126813 7315 127277 7611
rect 127573 7315 128037 7611
rect 128333 7315 128797 7611
rect 129093 7315 129557 7611
rect 129853 7315 130317 7611
rect 130613 7315 131077 7611
rect 131373 7315 131837 7611
rect 132133 7315 132597 7611
rect 132893 7315 133225 7611
rect 114025 7143 133225 7315
rect 135825 18251 155025 18713
rect 135825 17955 136157 18251
rect 136453 17955 136917 18251
rect 137213 17955 137677 18251
rect 137973 17955 138437 18251
rect 138733 17955 139197 18251
rect 139493 17955 139957 18251
rect 140253 17955 140717 18251
rect 141013 17955 141477 18251
rect 141773 17955 142237 18251
rect 142533 17955 142997 18251
rect 143293 17955 143757 18251
rect 144053 17955 144517 18251
rect 144813 17955 145277 18251
rect 145573 17955 146037 18251
rect 146333 17955 146797 18251
rect 147093 17955 147557 18251
rect 147853 17955 148317 18251
rect 148613 17955 149077 18251
rect 149373 17955 149837 18251
rect 150133 17955 150597 18251
rect 150893 17955 151357 18251
rect 151653 17955 152117 18251
rect 152413 17955 152877 18251
rect 153173 17955 153637 18251
rect 153933 17955 154397 18251
rect 154693 17955 155025 18251
rect 135825 17491 155025 17955
rect 135825 17195 136157 17491
rect 136453 17195 136917 17491
rect 137213 17195 137677 17491
rect 137973 17195 138437 17491
rect 138733 17195 139197 17491
rect 139493 17195 139957 17491
rect 140253 17195 140717 17491
rect 141013 17195 141477 17491
rect 141773 17195 142237 17491
rect 142533 17195 142997 17491
rect 143293 17195 143757 17491
rect 144053 17195 144517 17491
rect 144813 17195 145277 17491
rect 145573 17195 146037 17491
rect 146333 17195 146797 17491
rect 147093 17195 147557 17491
rect 147853 17195 148317 17491
rect 148613 17195 149077 17491
rect 149373 17195 149837 17491
rect 150133 17195 150597 17491
rect 150893 17195 151357 17491
rect 151653 17195 152117 17491
rect 152413 17195 152877 17491
rect 153173 17195 153637 17491
rect 153933 17195 154397 17491
rect 154693 17195 155025 17491
rect 135825 16731 155025 17195
rect 135825 16435 136157 16731
rect 136453 16435 136917 16731
rect 137213 16435 137677 16731
rect 137973 16435 138437 16731
rect 138733 16435 139197 16731
rect 139493 16435 139957 16731
rect 140253 16435 140717 16731
rect 141013 16435 141477 16731
rect 141773 16435 142237 16731
rect 142533 16435 142997 16731
rect 143293 16435 143757 16731
rect 144053 16435 144517 16731
rect 144813 16435 145277 16731
rect 145573 16435 146037 16731
rect 146333 16435 146797 16731
rect 147093 16435 147557 16731
rect 147853 16435 148317 16731
rect 148613 16435 149077 16731
rect 149373 16435 149837 16731
rect 150133 16435 150597 16731
rect 150893 16435 151357 16731
rect 151653 16435 152117 16731
rect 152413 16435 152877 16731
rect 153173 16435 153637 16731
rect 153933 16435 154397 16731
rect 154693 16435 155025 16731
rect 135825 15971 155025 16435
rect 135825 15675 136157 15971
rect 136453 15675 136917 15971
rect 137213 15675 137677 15971
rect 137973 15675 138437 15971
rect 138733 15675 139197 15971
rect 139493 15675 139957 15971
rect 140253 15675 140717 15971
rect 141013 15675 141477 15971
rect 141773 15675 142237 15971
rect 142533 15675 142997 15971
rect 143293 15675 143757 15971
rect 144053 15675 144517 15971
rect 144813 15675 145277 15971
rect 145573 15675 146037 15971
rect 146333 15675 146797 15971
rect 147093 15675 147557 15971
rect 147853 15675 148317 15971
rect 148613 15675 149077 15971
rect 149373 15675 149837 15971
rect 150133 15675 150597 15971
rect 150893 15675 151357 15971
rect 151653 15675 152117 15971
rect 152413 15675 152877 15971
rect 153173 15675 153637 15971
rect 153933 15675 154397 15971
rect 154693 15675 155025 15971
rect 135825 15211 155025 15675
rect 135825 14915 136157 15211
rect 136453 14915 136917 15211
rect 137213 14915 137677 15211
rect 137973 14915 138437 15211
rect 138733 14915 139197 15211
rect 139493 14915 139957 15211
rect 140253 14915 140717 15211
rect 141013 14915 141477 15211
rect 141773 14915 142237 15211
rect 142533 14915 142997 15211
rect 143293 14915 143757 15211
rect 144053 14915 144517 15211
rect 144813 14915 145277 15211
rect 145573 14915 146037 15211
rect 146333 14915 146797 15211
rect 147093 14915 147557 15211
rect 147853 14915 148317 15211
rect 148613 14915 149077 15211
rect 149373 14915 149837 15211
rect 150133 14915 150597 15211
rect 150893 14915 151357 15211
rect 151653 14915 152117 15211
rect 152413 14915 152877 15211
rect 153173 14915 153637 15211
rect 153933 14915 154397 15211
rect 154693 14915 155025 15211
rect 135825 14451 155025 14915
rect 135825 14155 136157 14451
rect 136453 14155 136917 14451
rect 137213 14155 137677 14451
rect 137973 14155 138437 14451
rect 138733 14155 139197 14451
rect 139493 14155 139957 14451
rect 140253 14155 140717 14451
rect 141013 14155 141477 14451
rect 141773 14155 142237 14451
rect 142533 14155 142997 14451
rect 143293 14155 143757 14451
rect 144053 14155 144517 14451
rect 144813 14155 145277 14451
rect 145573 14155 146037 14451
rect 146333 14155 146797 14451
rect 147093 14155 147557 14451
rect 147853 14155 148317 14451
rect 148613 14155 149077 14451
rect 149373 14155 149837 14451
rect 150133 14155 150597 14451
rect 150893 14155 151357 14451
rect 151653 14155 152117 14451
rect 152413 14155 152877 14451
rect 153173 14155 153637 14451
rect 153933 14155 154397 14451
rect 154693 14155 155025 14451
rect 135825 13691 155025 14155
rect 135825 13395 136157 13691
rect 136453 13395 136917 13691
rect 137213 13395 137677 13691
rect 137973 13395 138437 13691
rect 138733 13395 139197 13691
rect 139493 13395 139957 13691
rect 140253 13395 140717 13691
rect 141013 13395 141477 13691
rect 141773 13395 142237 13691
rect 142533 13395 142997 13691
rect 143293 13395 143757 13691
rect 144053 13395 144517 13691
rect 144813 13395 145277 13691
rect 145573 13395 146037 13691
rect 146333 13395 146797 13691
rect 147093 13395 147557 13691
rect 147853 13395 148317 13691
rect 148613 13395 149077 13691
rect 149373 13395 149837 13691
rect 150133 13395 150597 13691
rect 150893 13395 151357 13691
rect 151653 13395 152117 13691
rect 152413 13395 152877 13691
rect 153173 13395 153637 13691
rect 153933 13395 154397 13691
rect 154693 13395 155025 13691
rect 135825 12931 155025 13395
rect 135825 12635 136157 12931
rect 136453 12635 136917 12931
rect 137213 12635 137677 12931
rect 137973 12635 138437 12931
rect 138733 12635 139197 12931
rect 139493 12635 139957 12931
rect 140253 12635 140717 12931
rect 141013 12635 141477 12931
rect 141773 12635 142237 12931
rect 142533 12635 142997 12931
rect 143293 12635 143757 12931
rect 144053 12635 144517 12931
rect 144813 12635 145277 12931
rect 145573 12635 146037 12931
rect 146333 12635 146797 12931
rect 147093 12635 147557 12931
rect 147853 12635 148317 12931
rect 148613 12635 149077 12931
rect 149373 12635 149837 12931
rect 150133 12635 150597 12931
rect 150893 12635 151357 12931
rect 151653 12635 152117 12931
rect 152413 12635 152877 12931
rect 153173 12635 153637 12931
rect 153933 12635 154397 12931
rect 154693 12635 155025 12931
rect 135825 12171 155025 12635
rect 135825 11875 136157 12171
rect 136453 11875 136917 12171
rect 137213 11875 137677 12171
rect 137973 11875 138437 12171
rect 138733 11875 139197 12171
rect 139493 11875 139957 12171
rect 140253 11875 140717 12171
rect 141013 11875 141477 12171
rect 141773 11875 142237 12171
rect 142533 11875 142997 12171
rect 143293 11875 143757 12171
rect 144053 11875 144517 12171
rect 144813 11875 145277 12171
rect 145573 11875 146037 12171
rect 146333 11875 146797 12171
rect 147093 11875 147557 12171
rect 147853 11875 148317 12171
rect 148613 11875 149077 12171
rect 149373 11875 149837 12171
rect 150133 11875 150597 12171
rect 150893 11875 151357 12171
rect 151653 11875 152117 12171
rect 152413 11875 152877 12171
rect 153173 11875 153637 12171
rect 153933 11875 154397 12171
rect 154693 11875 155025 12171
rect 135825 11411 155025 11875
rect 135825 11115 136157 11411
rect 136453 11115 136917 11411
rect 137213 11115 137677 11411
rect 137973 11115 138437 11411
rect 138733 11115 139197 11411
rect 139493 11115 139957 11411
rect 140253 11115 140717 11411
rect 141013 11115 141477 11411
rect 141773 11115 142237 11411
rect 142533 11115 142997 11411
rect 143293 11115 143757 11411
rect 144053 11115 144517 11411
rect 144813 11115 145277 11411
rect 145573 11115 146037 11411
rect 146333 11115 146797 11411
rect 147093 11115 147557 11411
rect 147853 11115 148317 11411
rect 148613 11115 149077 11411
rect 149373 11115 149837 11411
rect 150133 11115 150597 11411
rect 150893 11115 151357 11411
rect 151653 11115 152117 11411
rect 152413 11115 152877 11411
rect 153173 11115 153637 11411
rect 153933 11115 154397 11411
rect 154693 11115 155025 11411
rect 135825 10651 155025 11115
rect 135825 10355 136157 10651
rect 136453 10355 136917 10651
rect 137213 10355 137677 10651
rect 137973 10355 138437 10651
rect 138733 10355 139197 10651
rect 139493 10355 139957 10651
rect 140253 10355 140717 10651
rect 141013 10355 141477 10651
rect 141773 10355 142237 10651
rect 142533 10355 142997 10651
rect 143293 10355 143757 10651
rect 144053 10355 144517 10651
rect 144813 10355 145277 10651
rect 145573 10355 146037 10651
rect 146333 10355 146797 10651
rect 147093 10355 147557 10651
rect 147853 10355 148317 10651
rect 148613 10355 149077 10651
rect 149373 10355 149837 10651
rect 150133 10355 150597 10651
rect 150893 10355 151357 10651
rect 151653 10355 152117 10651
rect 152413 10355 152877 10651
rect 153173 10355 153637 10651
rect 153933 10355 154397 10651
rect 154693 10355 155025 10651
rect 135825 9891 155025 10355
rect 135825 9595 136157 9891
rect 136453 9595 136917 9891
rect 137213 9595 137677 9891
rect 137973 9595 138437 9891
rect 138733 9595 139197 9891
rect 139493 9595 139957 9891
rect 140253 9595 140717 9891
rect 141013 9595 141477 9891
rect 141773 9595 142237 9891
rect 142533 9595 142997 9891
rect 143293 9595 143757 9891
rect 144053 9595 144517 9891
rect 144813 9595 145277 9891
rect 145573 9595 146037 9891
rect 146333 9595 146797 9891
rect 147093 9595 147557 9891
rect 147853 9595 148317 9891
rect 148613 9595 149077 9891
rect 149373 9595 149837 9891
rect 150133 9595 150597 9891
rect 150893 9595 151357 9891
rect 151653 9595 152117 9891
rect 152413 9595 152877 9891
rect 153173 9595 153637 9891
rect 153933 9595 154397 9891
rect 154693 9595 155025 9891
rect 135825 9131 155025 9595
rect 135825 8835 136157 9131
rect 136453 8835 136917 9131
rect 137213 8835 137677 9131
rect 137973 8835 138437 9131
rect 138733 8835 139197 9131
rect 139493 8835 139957 9131
rect 140253 8835 140717 9131
rect 141013 8835 141477 9131
rect 141773 8835 142237 9131
rect 142533 8835 142997 9131
rect 143293 8835 143757 9131
rect 144053 8835 144517 9131
rect 144813 8835 145277 9131
rect 145573 8835 146037 9131
rect 146333 8835 146797 9131
rect 147093 8835 147557 9131
rect 147853 8835 148317 9131
rect 148613 8835 149077 9131
rect 149373 8835 149837 9131
rect 150133 8835 150597 9131
rect 150893 8835 151357 9131
rect 151653 8835 152117 9131
rect 152413 8835 152877 9131
rect 153173 8835 153637 9131
rect 153933 8835 154397 9131
rect 154693 8835 155025 9131
rect 135825 8371 155025 8835
rect 135825 8075 136157 8371
rect 136453 8075 136917 8371
rect 137213 8075 137677 8371
rect 137973 8075 138437 8371
rect 138733 8075 139197 8371
rect 139493 8075 139957 8371
rect 140253 8075 140717 8371
rect 141013 8075 141477 8371
rect 141773 8075 142237 8371
rect 142533 8075 142997 8371
rect 143293 8075 143757 8371
rect 144053 8075 144517 8371
rect 144813 8075 145277 8371
rect 145573 8075 146037 8371
rect 146333 8075 146797 8371
rect 147093 8075 147557 8371
rect 147853 8075 148317 8371
rect 148613 8075 149077 8371
rect 149373 8075 149837 8371
rect 150133 8075 150597 8371
rect 150893 8075 151357 8371
rect 151653 8075 152117 8371
rect 152413 8075 152877 8371
rect 153173 8075 153637 8371
rect 153933 8075 154397 8371
rect 154693 8075 155025 8371
rect 135825 7611 155025 8075
rect 135825 7315 136157 7611
rect 136453 7315 136917 7611
rect 137213 7315 137677 7611
rect 137973 7315 138437 7611
rect 138733 7315 139197 7611
rect 139493 7315 139957 7611
rect 140253 7315 140717 7611
rect 141013 7315 141477 7611
rect 141773 7315 142237 7611
rect 142533 7315 142997 7611
rect 143293 7315 143757 7611
rect 144053 7315 144517 7611
rect 144813 7315 145277 7611
rect 145573 7315 146037 7611
rect 146333 7315 146797 7611
rect 147093 7315 147557 7611
rect 147853 7315 148317 7611
rect 148613 7315 149077 7611
rect 149373 7315 149837 7611
rect 150133 7315 150597 7611
rect 150893 7315 151357 7611
rect 151653 7315 152117 7611
rect 152413 7315 152877 7611
rect 153173 7315 153637 7611
rect 153933 7315 154397 7611
rect 154693 7315 155025 7611
rect 135825 7143 155025 7315
rect 157625 18251 176825 18713
rect 157625 17955 157957 18251
rect 158253 17955 158717 18251
rect 159013 17955 159477 18251
rect 159773 17955 160237 18251
rect 160533 17955 160997 18251
rect 161293 17955 161757 18251
rect 162053 17955 162517 18251
rect 162813 17955 163277 18251
rect 163573 17955 164037 18251
rect 164333 17955 164797 18251
rect 165093 17955 165557 18251
rect 165853 17955 166317 18251
rect 166613 17955 167077 18251
rect 167373 17955 167837 18251
rect 168133 17955 168597 18251
rect 168893 17955 169357 18251
rect 169653 17955 170117 18251
rect 170413 17955 170877 18251
rect 171173 17955 171637 18251
rect 171933 17955 172397 18251
rect 172693 17955 173157 18251
rect 173453 17955 173917 18251
rect 174213 17955 174677 18251
rect 174973 17955 175437 18251
rect 175733 17955 176197 18251
rect 176493 17955 176825 18251
rect 157625 17491 176825 17955
rect 157625 17195 157957 17491
rect 158253 17195 158717 17491
rect 159013 17195 159477 17491
rect 159773 17195 160237 17491
rect 160533 17195 160997 17491
rect 161293 17195 161757 17491
rect 162053 17195 162517 17491
rect 162813 17195 163277 17491
rect 163573 17195 164037 17491
rect 164333 17195 164797 17491
rect 165093 17195 165557 17491
rect 165853 17195 166317 17491
rect 166613 17195 167077 17491
rect 167373 17195 167837 17491
rect 168133 17195 168597 17491
rect 168893 17195 169357 17491
rect 169653 17195 170117 17491
rect 170413 17195 170877 17491
rect 171173 17195 171637 17491
rect 171933 17195 172397 17491
rect 172693 17195 173157 17491
rect 173453 17195 173917 17491
rect 174213 17195 174677 17491
rect 174973 17195 175437 17491
rect 175733 17195 176197 17491
rect 176493 17195 176825 17491
rect 157625 16731 176825 17195
rect 157625 16435 157957 16731
rect 158253 16435 158717 16731
rect 159013 16435 159477 16731
rect 159773 16435 160237 16731
rect 160533 16435 160997 16731
rect 161293 16435 161757 16731
rect 162053 16435 162517 16731
rect 162813 16435 163277 16731
rect 163573 16435 164037 16731
rect 164333 16435 164797 16731
rect 165093 16435 165557 16731
rect 165853 16435 166317 16731
rect 166613 16435 167077 16731
rect 167373 16435 167837 16731
rect 168133 16435 168597 16731
rect 168893 16435 169357 16731
rect 169653 16435 170117 16731
rect 170413 16435 170877 16731
rect 171173 16435 171637 16731
rect 171933 16435 172397 16731
rect 172693 16435 173157 16731
rect 173453 16435 173917 16731
rect 174213 16435 174677 16731
rect 174973 16435 175437 16731
rect 175733 16435 176197 16731
rect 176493 16435 176825 16731
rect 157625 15971 176825 16435
rect 157625 15675 157957 15971
rect 158253 15675 158717 15971
rect 159013 15675 159477 15971
rect 159773 15675 160237 15971
rect 160533 15675 160997 15971
rect 161293 15675 161757 15971
rect 162053 15675 162517 15971
rect 162813 15675 163277 15971
rect 163573 15675 164037 15971
rect 164333 15675 164797 15971
rect 165093 15675 165557 15971
rect 165853 15675 166317 15971
rect 166613 15675 167077 15971
rect 167373 15675 167837 15971
rect 168133 15675 168597 15971
rect 168893 15675 169357 15971
rect 169653 15675 170117 15971
rect 170413 15675 170877 15971
rect 171173 15675 171637 15971
rect 171933 15675 172397 15971
rect 172693 15675 173157 15971
rect 173453 15675 173917 15971
rect 174213 15675 174677 15971
rect 174973 15675 175437 15971
rect 175733 15675 176197 15971
rect 176493 15675 176825 15971
rect 157625 15211 176825 15675
rect 157625 14915 157957 15211
rect 158253 14915 158717 15211
rect 159013 14915 159477 15211
rect 159773 14915 160237 15211
rect 160533 14915 160997 15211
rect 161293 14915 161757 15211
rect 162053 14915 162517 15211
rect 162813 14915 163277 15211
rect 163573 14915 164037 15211
rect 164333 14915 164797 15211
rect 165093 14915 165557 15211
rect 165853 14915 166317 15211
rect 166613 14915 167077 15211
rect 167373 14915 167837 15211
rect 168133 14915 168597 15211
rect 168893 14915 169357 15211
rect 169653 14915 170117 15211
rect 170413 14915 170877 15211
rect 171173 14915 171637 15211
rect 171933 14915 172397 15211
rect 172693 14915 173157 15211
rect 173453 14915 173917 15211
rect 174213 14915 174677 15211
rect 174973 14915 175437 15211
rect 175733 14915 176197 15211
rect 176493 14915 176825 15211
rect 157625 14451 176825 14915
rect 157625 14155 157957 14451
rect 158253 14155 158717 14451
rect 159013 14155 159477 14451
rect 159773 14155 160237 14451
rect 160533 14155 160997 14451
rect 161293 14155 161757 14451
rect 162053 14155 162517 14451
rect 162813 14155 163277 14451
rect 163573 14155 164037 14451
rect 164333 14155 164797 14451
rect 165093 14155 165557 14451
rect 165853 14155 166317 14451
rect 166613 14155 167077 14451
rect 167373 14155 167837 14451
rect 168133 14155 168597 14451
rect 168893 14155 169357 14451
rect 169653 14155 170117 14451
rect 170413 14155 170877 14451
rect 171173 14155 171637 14451
rect 171933 14155 172397 14451
rect 172693 14155 173157 14451
rect 173453 14155 173917 14451
rect 174213 14155 174677 14451
rect 174973 14155 175437 14451
rect 175733 14155 176197 14451
rect 176493 14155 176825 14451
rect 157625 13691 176825 14155
rect 157625 13395 157957 13691
rect 158253 13395 158717 13691
rect 159013 13395 159477 13691
rect 159773 13395 160237 13691
rect 160533 13395 160997 13691
rect 161293 13395 161757 13691
rect 162053 13395 162517 13691
rect 162813 13395 163277 13691
rect 163573 13395 164037 13691
rect 164333 13395 164797 13691
rect 165093 13395 165557 13691
rect 165853 13395 166317 13691
rect 166613 13395 167077 13691
rect 167373 13395 167837 13691
rect 168133 13395 168597 13691
rect 168893 13395 169357 13691
rect 169653 13395 170117 13691
rect 170413 13395 170877 13691
rect 171173 13395 171637 13691
rect 171933 13395 172397 13691
rect 172693 13395 173157 13691
rect 173453 13395 173917 13691
rect 174213 13395 174677 13691
rect 174973 13395 175437 13691
rect 175733 13395 176197 13691
rect 176493 13395 176825 13691
rect 157625 12931 176825 13395
rect 157625 12635 157957 12931
rect 158253 12635 158717 12931
rect 159013 12635 159477 12931
rect 159773 12635 160237 12931
rect 160533 12635 160997 12931
rect 161293 12635 161757 12931
rect 162053 12635 162517 12931
rect 162813 12635 163277 12931
rect 163573 12635 164037 12931
rect 164333 12635 164797 12931
rect 165093 12635 165557 12931
rect 165853 12635 166317 12931
rect 166613 12635 167077 12931
rect 167373 12635 167837 12931
rect 168133 12635 168597 12931
rect 168893 12635 169357 12931
rect 169653 12635 170117 12931
rect 170413 12635 170877 12931
rect 171173 12635 171637 12931
rect 171933 12635 172397 12931
rect 172693 12635 173157 12931
rect 173453 12635 173917 12931
rect 174213 12635 174677 12931
rect 174973 12635 175437 12931
rect 175733 12635 176197 12931
rect 176493 12635 176825 12931
rect 157625 12171 176825 12635
rect 157625 11875 157957 12171
rect 158253 11875 158717 12171
rect 159013 11875 159477 12171
rect 159773 11875 160237 12171
rect 160533 11875 160997 12171
rect 161293 11875 161757 12171
rect 162053 11875 162517 12171
rect 162813 11875 163277 12171
rect 163573 11875 164037 12171
rect 164333 11875 164797 12171
rect 165093 11875 165557 12171
rect 165853 11875 166317 12171
rect 166613 11875 167077 12171
rect 167373 11875 167837 12171
rect 168133 11875 168597 12171
rect 168893 11875 169357 12171
rect 169653 11875 170117 12171
rect 170413 11875 170877 12171
rect 171173 11875 171637 12171
rect 171933 11875 172397 12171
rect 172693 11875 173157 12171
rect 173453 11875 173917 12171
rect 174213 11875 174677 12171
rect 174973 11875 175437 12171
rect 175733 11875 176197 12171
rect 176493 11875 176825 12171
rect 157625 11411 176825 11875
rect 157625 11115 157957 11411
rect 158253 11115 158717 11411
rect 159013 11115 159477 11411
rect 159773 11115 160237 11411
rect 160533 11115 160997 11411
rect 161293 11115 161757 11411
rect 162053 11115 162517 11411
rect 162813 11115 163277 11411
rect 163573 11115 164037 11411
rect 164333 11115 164797 11411
rect 165093 11115 165557 11411
rect 165853 11115 166317 11411
rect 166613 11115 167077 11411
rect 167373 11115 167837 11411
rect 168133 11115 168597 11411
rect 168893 11115 169357 11411
rect 169653 11115 170117 11411
rect 170413 11115 170877 11411
rect 171173 11115 171637 11411
rect 171933 11115 172397 11411
rect 172693 11115 173157 11411
rect 173453 11115 173917 11411
rect 174213 11115 174677 11411
rect 174973 11115 175437 11411
rect 175733 11115 176197 11411
rect 176493 11115 176825 11411
rect 157625 10651 176825 11115
rect 157625 10355 157957 10651
rect 158253 10355 158717 10651
rect 159013 10355 159477 10651
rect 159773 10355 160237 10651
rect 160533 10355 160997 10651
rect 161293 10355 161757 10651
rect 162053 10355 162517 10651
rect 162813 10355 163277 10651
rect 163573 10355 164037 10651
rect 164333 10355 164797 10651
rect 165093 10355 165557 10651
rect 165853 10355 166317 10651
rect 166613 10355 167077 10651
rect 167373 10355 167837 10651
rect 168133 10355 168597 10651
rect 168893 10355 169357 10651
rect 169653 10355 170117 10651
rect 170413 10355 170877 10651
rect 171173 10355 171637 10651
rect 171933 10355 172397 10651
rect 172693 10355 173157 10651
rect 173453 10355 173917 10651
rect 174213 10355 174677 10651
rect 174973 10355 175437 10651
rect 175733 10355 176197 10651
rect 176493 10355 176825 10651
rect 157625 9891 176825 10355
rect 186905 18344 211105 18713
rect 186905 18048 187077 18344
rect 187373 18048 187837 18344
rect 188133 18048 188597 18344
rect 188893 18048 189357 18344
rect 189653 18048 190117 18344
rect 190413 18048 190877 18344
rect 191173 18048 191637 18344
rect 191933 18048 192397 18344
rect 192693 18048 193157 18344
rect 193453 18048 193917 18344
rect 194213 18048 194677 18344
rect 194973 18048 195437 18344
rect 195733 18048 196197 18344
rect 196493 18048 196957 18344
rect 197253 18048 197717 18344
rect 198013 18048 198477 18344
rect 198773 18048 199237 18344
rect 199533 18048 199997 18344
rect 200293 18048 200757 18344
rect 201053 18048 201517 18344
rect 201813 18048 202277 18344
rect 202573 18048 203037 18344
rect 203333 18048 203797 18344
rect 204093 18048 204557 18344
rect 204853 18048 205317 18344
rect 205613 18048 206077 18344
rect 206373 18048 206837 18344
rect 207133 18048 207597 18344
rect 207893 18048 208357 18344
rect 208653 18048 209117 18344
rect 209413 18048 209877 18344
rect 210173 18048 210637 18344
rect 210933 18048 211105 18344
rect 186905 17584 211105 18048
rect 186905 17288 187077 17584
rect 187373 17288 187837 17584
rect 188133 17288 188597 17584
rect 188893 17288 189357 17584
rect 189653 17288 190117 17584
rect 190413 17288 190877 17584
rect 191173 17288 191637 17584
rect 191933 17288 192397 17584
rect 192693 17288 193157 17584
rect 193453 17288 193917 17584
rect 194213 17288 194677 17584
rect 194973 17288 195437 17584
rect 195733 17288 196197 17584
rect 196493 17288 196957 17584
rect 197253 17288 197717 17584
rect 198013 17288 198477 17584
rect 198773 17288 199237 17584
rect 199533 17288 199997 17584
rect 200293 17288 200757 17584
rect 201053 17288 201517 17584
rect 201813 17288 202277 17584
rect 202573 17288 203037 17584
rect 203333 17288 203797 17584
rect 204093 17288 204557 17584
rect 204853 17288 205317 17584
rect 205613 17288 206077 17584
rect 206373 17288 206837 17584
rect 207133 17288 207597 17584
rect 207893 17288 208357 17584
rect 208653 17288 209117 17584
rect 209413 17288 209877 17584
rect 210173 17288 210637 17584
rect 210933 17288 211105 17584
rect 186905 16824 211105 17288
rect 186905 16528 187077 16824
rect 187373 16528 187837 16824
rect 188133 16528 188597 16824
rect 188893 16528 189357 16824
rect 189653 16528 190117 16824
rect 190413 16528 190877 16824
rect 191173 16528 191637 16824
rect 191933 16528 192397 16824
rect 192693 16528 193157 16824
rect 193453 16528 193917 16824
rect 194213 16528 194677 16824
rect 194973 16528 195437 16824
rect 195733 16528 196197 16824
rect 196493 16528 196957 16824
rect 197253 16528 197717 16824
rect 198013 16528 198477 16824
rect 198773 16528 199237 16824
rect 199533 16528 199997 16824
rect 200293 16528 200757 16824
rect 201053 16528 201517 16824
rect 201813 16528 202277 16824
rect 202573 16528 203037 16824
rect 203333 16528 203797 16824
rect 204093 16528 204557 16824
rect 204853 16528 205317 16824
rect 205613 16528 206077 16824
rect 206373 16528 206837 16824
rect 207133 16528 207597 16824
rect 207893 16528 208357 16824
rect 208653 16528 209117 16824
rect 209413 16528 209877 16824
rect 210173 16528 210637 16824
rect 210933 16528 211105 16824
rect 186905 16064 211105 16528
rect 186905 15768 187077 16064
rect 187373 15768 187837 16064
rect 188133 15768 188597 16064
rect 188893 15768 189357 16064
rect 189653 15768 190117 16064
rect 190413 15768 190877 16064
rect 191173 15768 191637 16064
rect 191933 15768 192397 16064
rect 192693 15768 193157 16064
rect 193453 15768 193917 16064
rect 194213 15768 194677 16064
rect 194973 15768 195437 16064
rect 195733 15768 196197 16064
rect 196493 15768 196957 16064
rect 197253 15768 197717 16064
rect 198013 15768 198477 16064
rect 198773 15768 199237 16064
rect 199533 15768 199997 16064
rect 200293 15768 200757 16064
rect 201053 15768 201517 16064
rect 201813 15768 202277 16064
rect 202573 15768 203037 16064
rect 203333 15768 203797 16064
rect 204093 15768 204557 16064
rect 204853 15768 205317 16064
rect 205613 15768 206077 16064
rect 206373 15768 206837 16064
rect 207133 15768 207597 16064
rect 207893 15768 208357 16064
rect 208653 15768 209117 16064
rect 209413 15768 209877 16064
rect 210173 15768 210637 16064
rect 210933 15768 211105 16064
rect 186905 15304 211105 15768
rect 186905 15008 187077 15304
rect 187373 15008 187837 15304
rect 188133 15008 188597 15304
rect 188893 15008 189357 15304
rect 189653 15008 190117 15304
rect 190413 15008 190877 15304
rect 191173 15008 191637 15304
rect 191933 15008 192397 15304
rect 192693 15008 193157 15304
rect 193453 15008 193917 15304
rect 194213 15008 194677 15304
rect 194973 15008 195437 15304
rect 195733 15008 196197 15304
rect 196493 15008 196957 15304
rect 197253 15008 197717 15304
rect 198013 15008 198477 15304
rect 198773 15008 199237 15304
rect 199533 15008 199997 15304
rect 200293 15008 200757 15304
rect 201053 15008 201517 15304
rect 201813 15008 202277 15304
rect 202573 15008 203037 15304
rect 203333 15008 203797 15304
rect 204093 15008 204557 15304
rect 204853 15008 205317 15304
rect 205613 15008 206077 15304
rect 206373 15008 206837 15304
rect 207133 15008 207597 15304
rect 207893 15008 208357 15304
rect 208653 15008 209117 15304
rect 209413 15008 209877 15304
rect 210173 15008 210637 15304
rect 210933 15008 211105 15304
rect 186905 14544 211105 15008
rect 186905 14248 187077 14544
rect 187373 14248 187837 14544
rect 188133 14248 188597 14544
rect 188893 14248 189357 14544
rect 189653 14248 190117 14544
rect 190413 14248 190877 14544
rect 191173 14248 191637 14544
rect 191933 14248 192397 14544
rect 192693 14248 193157 14544
rect 193453 14248 193917 14544
rect 194213 14248 194677 14544
rect 194973 14248 195437 14544
rect 195733 14248 196197 14544
rect 196493 14248 196957 14544
rect 197253 14248 197717 14544
rect 198013 14248 198477 14544
rect 198773 14248 199237 14544
rect 199533 14248 199997 14544
rect 200293 14248 200757 14544
rect 201053 14248 201517 14544
rect 201813 14248 202277 14544
rect 202573 14248 203037 14544
rect 203333 14248 203797 14544
rect 204093 14248 204557 14544
rect 204853 14248 205317 14544
rect 205613 14248 206077 14544
rect 206373 14248 206837 14544
rect 207133 14248 207597 14544
rect 207893 14248 208357 14544
rect 208653 14248 209117 14544
rect 209413 14248 209877 14544
rect 210173 14248 210637 14544
rect 210933 14248 211105 14544
rect 186905 13784 211105 14248
rect 186905 13488 187077 13784
rect 187373 13488 187837 13784
rect 188133 13488 188597 13784
rect 188893 13488 189357 13784
rect 189653 13488 190117 13784
rect 190413 13488 190877 13784
rect 191173 13488 191637 13784
rect 191933 13488 192397 13784
rect 192693 13488 193157 13784
rect 193453 13488 193917 13784
rect 194213 13488 194677 13784
rect 194973 13488 195437 13784
rect 195733 13488 196197 13784
rect 196493 13488 196957 13784
rect 197253 13488 197717 13784
rect 198013 13488 198477 13784
rect 198773 13488 199237 13784
rect 199533 13488 199997 13784
rect 200293 13488 200757 13784
rect 201053 13488 201517 13784
rect 201813 13488 202277 13784
rect 202573 13488 203037 13784
rect 203333 13488 203797 13784
rect 204093 13488 204557 13784
rect 204853 13488 205317 13784
rect 205613 13488 206077 13784
rect 206373 13488 206837 13784
rect 207133 13488 207597 13784
rect 207893 13488 208357 13784
rect 208653 13488 209117 13784
rect 209413 13488 209877 13784
rect 210173 13488 210637 13784
rect 210933 13488 211105 13784
rect 186905 13024 211105 13488
rect 186905 12728 187077 13024
rect 187373 12728 187837 13024
rect 188133 12728 188597 13024
rect 188893 12728 189357 13024
rect 189653 12728 190117 13024
rect 190413 12728 190877 13024
rect 191173 12728 191637 13024
rect 191933 12728 192397 13024
rect 192693 12728 193157 13024
rect 193453 12728 193917 13024
rect 194213 12728 194677 13024
rect 194973 12728 195437 13024
rect 195733 12728 196197 13024
rect 196493 12728 196957 13024
rect 197253 12728 197717 13024
rect 198013 12728 198477 13024
rect 198773 12728 199237 13024
rect 199533 12728 199997 13024
rect 200293 12728 200757 13024
rect 201053 12728 201517 13024
rect 201813 12728 202277 13024
rect 202573 12728 203037 13024
rect 203333 12728 203797 13024
rect 204093 12728 204557 13024
rect 204853 12728 205317 13024
rect 205613 12728 206077 13024
rect 206373 12728 206837 13024
rect 207133 12728 207597 13024
rect 207893 12728 208357 13024
rect 208653 12728 209117 13024
rect 209413 12728 209877 13024
rect 210173 12728 210637 13024
rect 210933 12728 211105 13024
rect 186905 12264 211105 12728
rect 186905 11968 187077 12264
rect 187373 11968 187837 12264
rect 188133 11968 188597 12264
rect 188893 11968 189357 12264
rect 189653 11968 190117 12264
rect 190413 11968 190877 12264
rect 191173 11968 191637 12264
rect 191933 11968 192397 12264
rect 192693 11968 193157 12264
rect 193453 11968 193917 12264
rect 194213 11968 194677 12264
rect 194973 11968 195437 12264
rect 195733 11968 196197 12264
rect 196493 11968 196957 12264
rect 197253 11968 197717 12264
rect 198013 11968 198477 12264
rect 198773 11968 199237 12264
rect 199533 11968 199997 12264
rect 200293 11968 200757 12264
rect 201053 11968 201517 12264
rect 201813 11968 202277 12264
rect 202573 11968 203037 12264
rect 203333 11968 203797 12264
rect 204093 11968 204557 12264
rect 204853 11968 205317 12264
rect 205613 11968 206077 12264
rect 206373 11968 206837 12264
rect 207133 11968 207597 12264
rect 207893 11968 208357 12264
rect 208653 11968 209117 12264
rect 209413 11968 209877 12264
rect 210173 11968 210637 12264
rect 210933 11968 211105 12264
rect 186905 11504 211105 11968
rect 186905 11208 187077 11504
rect 187373 11208 187837 11504
rect 188133 11208 188597 11504
rect 188893 11208 189357 11504
rect 189653 11208 190117 11504
rect 190413 11208 190877 11504
rect 191173 11208 191637 11504
rect 191933 11208 192397 11504
rect 192693 11208 193157 11504
rect 193453 11208 193917 11504
rect 194213 11208 194677 11504
rect 194973 11208 195437 11504
rect 195733 11208 196197 11504
rect 196493 11208 196957 11504
rect 197253 11208 197717 11504
rect 198013 11208 198477 11504
rect 198773 11208 199237 11504
rect 199533 11208 199997 11504
rect 200293 11208 200757 11504
rect 201053 11208 201517 11504
rect 201813 11208 202277 11504
rect 202573 11208 203037 11504
rect 203333 11208 203797 11504
rect 204093 11208 204557 11504
rect 204853 11208 205317 11504
rect 205613 11208 206077 11504
rect 206373 11208 206837 11504
rect 207133 11208 207597 11504
rect 207893 11208 208357 11504
rect 208653 11208 209117 11504
rect 209413 11208 209877 11504
rect 210173 11208 210637 11504
rect 210933 11208 211105 11504
rect 186905 10744 211105 11208
rect 186905 10448 187077 10744
rect 187373 10448 187837 10744
rect 188133 10448 188597 10744
rect 188893 10448 189357 10744
rect 189653 10448 190117 10744
rect 190413 10448 190877 10744
rect 191173 10448 191637 10744
rect 191933 10448 192397 10744
rect 192693 10448 193157 10744
rect 193453 10448 193917 10744
rect 194213 10448 194677 10744
rect 194973 10448 195437 10744
rect 195733 10448 196197 10744
rect 196493 10448 196957 10744
rect 197253 10448 197717 10744
rect 198013 10448 198477 10744
rect 198773 10448 199237 10744
rect 199533 10448 199997 10744
rect 200293 10448 200757 10744
rect 201053 10448 201517 10744
rect 201813 10448 202277 10744
rect 202573 10448 203037 10744
rect 203333 10448 203797 10744
rect 204093 10448 204557 10744
rect 204853 10448 205317 10744
rect 205613 10448 206077 10744
rect 206373 10448 206837 10744
rect 207133 10448 207597 10744
rect 207893 10448 208357 10744
rect 208653 10448 209117 10744
rect 209413 10448 209877 10744
rect 210173 10448 210637 10744
rect 210933 10448 211105 10744
rect 186905 10116 211105 10448
rect 212555 29208 212995 29464
rect 212555 28944 212643 29208
rect 212907 28944 212995 29208
rect 212555 28688 212995 28944
rect 212555 28424 212643 28688
rect 212907 28424 212995 28688
rect 212555 28168 212995 28424
rect 212555 27904 212643 28168
rect 212907 27904 212995 28168
rect 212555 27648 212995 27904
rect 212555 27384 212643 27648
rect 212907 27384 212995 27648
rect 212555 27128 212995 27384
rect 212555 26864 212643 27128
rect 212907 26864 212995 27128
rect 212555 26608 212995 26864
rect 212555 26344 212643 26608
rect 212907 26344 212995 26608
rect 212555 26088 212995 26344
rect 212555 25824 212643 26088
rect 212907 25824 212995 26088
rect 212555 25568 212995 25824
rect 212555 25304 212643 25568
rect 212907 25304 212995 25568
rect 212555 25048 212995 25304
rect 212555 24784 212643 25048
rect 212907 24784 212995 25048
rect 212555 24528 212995 24784
rect 212555 24264 212643 24528
rect 212907 24264 212995 24528
rect 212555 24008 212995 24264
rect 212555 23744 212643 24008
rect 212907 23744 212995 24008
rect 212555 23488 212995 23744
rect 212555 23224 212643 23488
rect 212907 23224 212995 23488
rect 212555 22968 212995 23224
rect 212555 22704 212643 22968
rect 212907 22704 212995 22968
rect 212555 22448 212995 22704
rect 212555 22184 212643 22448
rect 212907 22184 212995 22448
rect 212555 21928 212995 22184
rect 212555 21664 212643 21928
rect 212907 21664 212995 21928
rect 212555 21408 212995 21664
rect 212555 21144 212643 21408
rect 212907 21144 212995 21408
rect 212555 20888 212995 21144
rect 212555 20624 212643 20888
rect 212907 20624 212995 20888
rect 212555 20368 212995 20624
rect 212555 20104 212643 20368
rect 212907 20104 212995 20368
rect 212555 19848 212995 20104
rect 212555 19584 212643 19848
rect 212907 19584 212995 19848
rect 212555 19328 212995 19584
rect 212555 19064 212643 19328
rect 212907 19064 212995 19328
rect 212555 18808 212995 19064
rect 212555 18544 212643 18808
rect 212907 18544 212995 18808
rect 212555 18288 212995 18544
rect 212555 18024 212643 18288
rect 212907 18024 212995 18288
rect 212555 17768 212995 18024
rect 212555 17504 212643 17768
rect 212907 17504 212995 17768
rect 212555 17248 212995 17504
rect 212555 16984 212643 17248
rect 212907 16984 212995 17248
rect 212555 16728 212995 16984
rect 212555 16464 212643 16728
rect 212907 16464 212995 16728
rect 212555 16208 212995 16464
rect 212555 15944 212643 16208
rect 212907 15944 212995 16208
rect 212555 15688 212995 15944
rect 212555 15424 212643 15688
rect 212907 15424 212995 15688
rect 212555 15168 212995 15424
rect 212555 14904 212643 15168
rect 212907 14904 212995 15168
rect 212555 14648 212995 14904
rect 212555 14384 212643 14648
rect 212907 14384 212995 14648
rect 212555 14128 212995 14384
rect 212555 13864 212643 14128
rect 212907 13864 212995 14128
rect 212555 13608 212995 13864
rect 212555 13344 212643 13608
rect 212907 13344 212995 13608
rect 212555 13088 212995 13344
rect 212555 12824 212643 13088
rect 212907 12824 212995 13088
rect 212555 12568 212995 12824
rect 212555 12304 212643 12568
rect 212907 12304 212995 12568
rect 212555 12048 212995 12304
rect 212555 11784 212643 12048
rect 212907 11784 212995 12048
rect 212555 11528 212995 11784
rect 212555 11264 212643 11528
rect 212907 11264 212995 11528
rect 212555 11008 212995 11264
rect 212555 10744 212643 11008
rect 212907 10744 212995 11008
rect 212555 10488 212995 10744
rect 212555 10224 212643 10488
rect 212907 10224 212995 10488
rect 157625 9595 157957 9891
rect 158253 9595 158717 9891
rect 159013 9595 159477 9891
rect 159773 9595 160237 9891
rect 160533 9595 160997 9891
rect 161293 9595 161757 9891
rect 162053 9595 162517 9891
rect 162813 9595 163277 9891
rect 163573 9595 164037 9891
rect 164333 9595 164797 9891
rect 165093 9595 165557 9891
rect 165853 9595 166317 9891
rect 166613 9595 167077 9891
rect 167373 9595 167837 9891
rect 168133 9595 168597 9891
rect 168893 9595 169357 9891
rect 169653 9595 170117 9891
rect 170413 9595 170877 9891
rect 171173 9595 171637 9891
rect 171933 9595 172397 9891
rect 172693 9595 173157 9891
rect 173453 9595 173917 9891
rect 174213 9595 174677 9891
rect 174973 9595 175437 9891
rect 175733 9595 176197 9891
rect 176493 9595 176825 9891
rect 157625 9131 176825 9595
rect 212555 9968 212995 10224
rect 212555 9704 212643 9968
rect 212907 9704 212995 9968
rect 212555 9401 212995 9704
rect 157625 8835 157957 9131
rect 158253 8835 158717 9131
rect 159013 8835 159477 9131
rect 159773 8835 160237 9131
rect 160533 8835 160997 9131
rect 161293 8835 161757 9131
rect 162053 8835 162517 9131
rect 162813 8835 163277 9131
rect 163573 8835 164037 9131
rect 164333 8835 164797 9131
rect 165093 8835 165557 9131
rect 165853 8835 166317 9131
rect 166613 8835 167077 9131
rect 167373 8835 167837 9131
rect 168133 8835 168597 9131
rect 168893 8835 169357 9131
rect 169653 8835 170117 9131
rect 170413 8835 170877 9131
rect 171173 8835 171637 9131
rect 171933 8835 172397 9131
rect 172693 8835 173157 9131
rect 173453 8835 173917 9131
rect 174213 8835 174677 9131
rect 174973 8835 175437 9131
rect 175733 8835 176197 9131
rect 176493 8835 176825 9131
rect 157625 8371 176825 8835
rect 157625 8075 157957 8371
rect 158253 8075 158717 8371
rect 159013 8075 159477 8371
rect 159773 8075 160237 8371
rect 160533 8075 160997 8371
rect 161293 8075 161757 8371
rect 162053 8075 162517 8371
rect 162813 8075 163277 8371
rect 163573 8075 164037 8371
rect 164333 8075 164797 8371
rect 165093 8075 165557 8371
rect 165853 8075 166317 8371
rect 166613 8075 167077 8371
rect 167373 8075 167837 8371
rect 168133 8075 168597 8371
rect 168893 8075 169357 8371
rect 169653 8075 170117 8371
rect 170413 8075 170877 8371
rect 171173 8075 171637 8371
rect 171933 8075 172397 8371
rect 172693 8075 173157 8371
rect 173453 8075 173917 8371
rect 174213 8075 174677 8371
rect 174973 8075 175437 8371
rect 175733 8075 176197 8371
rect 176493 8075 176825 8371
rect 157625 7611 176825 8075
rect 157625 7315 157957 7611
rect 158253 7315 158717 7611
rect 159013 7315 159477 7611
rect 159773 7315 160237 7611
rect 160533 7315 160997 7611
rect 161293 7315 161757 7611
rect 162053 7315 162517 7611
rect 162813 7315 163277 7611
rect 163573 7315 164037 7611
rect 164333 7315 164797 7611
rect 165093 7315 165557 7611
rect 165853 7315 166317 7611
rect 166613 7315 167077 7611
rect 167373 7315 167837 7611
rect 168133 7315 168597 7611
rect 168893 7315 169357 7611
rect 169653 7315 170117 7611
rect 170413 7315 170877 7611
rect 171173 7315 171637 7611
rect 171933 7315 172397 7611
rect 172693 7315 173157 7611
rect 173453 7315 173917 7611
rect 174213 7315 174677 7611
rect 174973 7315 175437 7611
rect 175733 7315 176197 7611
rect 176493 7315 176825 7611
rect 157625 7143 176825 7315
rect 112725 5605 178125 6003
rect 112725 5341 113613 5605
rect 113877 5341 114133 5605
rect 114397 5341 114653 5605
rect 114917 5341 115173 5605
rect 115437 5341 115693 5605
rect 115957 5341 116213 5605
rect 116477 5341 116733 5605
rect 116997 5341 117253 5605
rect 117517 5341 117773 5605
rect 118037 5341 118293 5605
rect 118557 5341 118813 5605
rect 119077 5341 119333 5605
rect 119597 5341 119853 5605
rect 120117 5341 120373 5605
rect 120637 5341 120893 5605
rect 121157 5341 121413 5605
rect 121677 5341 121933 5605
rect 122197 5341 122453 5605
rect 122717 5341 122973 5605
rect 123237 5341 123493 5605
rect 123757 5341 124013 5605
rect 124277 5341 124533 5605
rect 124797 5341 125053 5605
rect 125317 5341 125573 5605
rect 125837 5341 126093 5605
rect 126357 5341 126613 5605
rect 126877 5341 127133 5605
rect 127397 5341 127653 5605
rect 127917 5341 128173 5605
rect 128437 5341 128693 5605
rect 128957 5341 129213 5605
rect 129477 5341 129733 5605
rect 129997 5341 130253 5605
rect 130517 5341 130773 5605
rect 131037 5341 131293 5605
rect 131557 5341 131813 5605
rect 132077 5341 132333 5605
rect 132597 5341 132853 5605
rect 133117 5341 133373 5605
rect 133637 5341 135413 5605
rect 135677 5341 135933 5605
rect 136197 5341 136453 5605
rect 136717 5341 136973 5605
rect 137237 5341 137493 5605
rect 137757 5341 138013 5605
rect 138277 5341 138533 5605
rect 138797 5341 139053 5605
rect 139317 5341 139573 5605
rect 139837 5341 140093 5605
rect 140357 5341 140613 5605
rect 140877 5341 141133 5605
rect 141397 5341 141653 5605
rect 141917 5341 142173 5605
rect 142437 5341 142693 5605
rect 142957 5341 143213 5605
rect 143477 5341 143733 5605
rect 143997 5341 144253 5605
rect 144517 5341 144773 5605
rect 145037 5341 145293 5605
rect 145557 5341 145813 5605
rect 146077 5341 146333 5605
rect 146597 5341 146853 5605
rect 147117 5341 147373 5605
rect 147637 5341 147893 5605
rect 148157 5341 148413 5605
rect 148677 5341 148933 5605
rect 149197 5341 149453 5605
rect 149717 5341 149973 5605
rect 150237 5341 150493 5605
rect 150757 5341 151013 5605
rect 151277 5341 151533 5605
rect 151797 5341 152053 5605
rect 152317 5341 152573 5605
rect 152837 5341 153093 5605
rect 153357 5341 153613 5605
rect 153877 5341 154133 5605
rect 154397 5341 154653 5605
rect 154917 5341 155173 5605
rect 155437 5341 157213 5605
rect 157477 5341 157733 5605
rect 157997 5341 158253 5605
rect 158517 5341 158773 5605
rect 159037 5341 159293 5605
rect 159557 5341 159813 5605
rect 160077 5341 160333 5605
rect 160597 5341 160853 5605
rect 161117 5341 161373 5605
rect 161637 5341 161893 5605
rect 162157 5341 162413 5605
rect 162677 5341 162933 5605
rect 163197 5341 163453 5605
rect 163717 5341 163973 5605
rect 164237 5341 164493 5605
rect 164757 5341 165013 5605
rect 165277 5341 165533 5605
rect 165797 5341 166053 5605
rect 166317 5341 166573 5605
rect 166837 5341 167093 5605
rect 167357 5341 167613 5605
rect 167877 5341 168133 5605
rect 168397 5341 168653 5605
rect 168917 5341 169173 5605
rect 169437 5341 169693 5605
rect 169957 5341 170213 5605
rect 170477 5341 170733 5605
rect 170997 5341 171253 5605
rect 171517 5341 171773 5605
rect 172037 5341 172293 5605
rect 172557 5341 172813 5605
rect 173077 5341 173333 5605
rect 173597 5341 173853 5605
rect 174117 5341 174373 5605
rect 174637 5341 174893 5605
rect 175157 5341 175413 5605
rect 175677 5341 175933 5605
rect 176197 5341 176453 5605
rect 176717 5341 176973 5605
rect 177237 5341 178125 5605
rect 112725 4943 178125 5341
use nfet$2  nfet$2_0
timestamp 1676577649
transform 1 0 -60096 0 1 -162352
box -152 -44 30474 20044
use nfet$2  nfet$2_1
timestamp 1676577649
transform 1 0 -26096 0 1 -162352
box -152 -44 30474 20044
use nfet$2  nfet$2_2
timestamp 1676577649
transform 1 0 7904 0 1 -162352
box -152 -44 30474 20044
use nfet$2  nfet$2_3
timestamp 1676577649
transform 1 0 41904 0 1 -162352
box -152 -44 30474 20044
use nfet$2  nfet$2_4
timestamp 1676577649
transform 1 0 75904 0 1 -162352
box -152 -44 30474 20044
use nfet$2  nfet$2_5
timestamp 1676577649
transform 1 0 109904 0 1 -162352
box -152 -44 30474 20044
use nfet$2  nfet$2_6
timestamp 1676577649
transform 1 0 143904 0 1 -162352
box -152 -44 30474 20044
use nfet$2  nfet$2_7
timestamp 1676577649
transform 1 0 146886 0 1 -103119
box -152 -44 30474 20044
use nfet$2  nfet$2_8
timestamp 1676577649
transform 1 0 114886 0 1 -103119
box -152 -44 30474 20044
use nfet$2  nfet$2_9
timestamp 1676577649
transform 1 0 82886 0 1 -103119
box -152 -44 30474 20044
use nfet$2  nfet$2_10
timestamp 1676577649
transform 1 0 50886 0 1 -103119
box -152 -44 30474 20044
use nfet$2  nfet$2_11
timestamp 1676577649
transform 1 0 18886 0 1 -103119
box -152 -44 30474 20044
use nfet$2  nfet$2_12
timestamp 1676577649
transform 1 0 -13114 0 1 -103119
box -152 -44 30474 20044
use nfet$2  nfet$2_13
timestamp 1676577649
transform 1 0 -45114 0 1 -103119
box -152 -44 30474 20044
use nfet$2  nfet$2_14
timestamp 1676577649
transform 1 0 -77114 0 1 -103119
box -152 -44 30474 20044
use nfet$2  nfet$2_15
timestamp 1676577649
transform 1 0 -109114 0 1 -103119
box -152 -44 30474 20044
use nfet$2  nfet$2_16
timestamp 1676577649
transform 1 0 146886 0 1 -129119
box -152 -44 30474 20044
use nfet$2  nfet$2_17
timestamp 1676577649
transform 1 0 114886 0 1 -129119
box -152 -44 30474 20044
use nfet$2  nfet$2_18
timestamp 1676577649
transform 1 0 82886 0 1 -129119
box -152 -44 30474 20044
use nfet$2  nfet$2_19
timestamp 1676577649
transform 1 0 50886 0 1 -129119
box -152 -44 30474 20044
use nfet$2  nfet$2_20
timestamp 1676577649
transform 1 0 18886 0 1 -129119
box -152 -44 30474 20044
use nfet$2  nfet$2_21
timestamp 1676577649
transform 1 0 -13114 0 1 -129119
box -152 -44 30474 20044
use nfet$2  nfet$2_22
timestamp 1676577649
transform 1 0 -45114 0 1 -129119
box -152 -44 30474 20044
use nfet$2  nfet$2_23
timestamp 1676577649
transform 1 0 -77114 0 1 -129119
box -152 -44 30474 20044
use nfet$2  nfet$2_24
timestamp 1676577649
transform 1 0 -109114 0 1 -129119
box -152 -44 30474 20044
use nfet$2  nfet$2_25
timestamp 1676577649
transform 1 0 146886 0 1 -48119
box -152 -44 30474 20044
use nfet$2  nfet$2_26
timestamp 1676577649
transform 1 0 114886 0 1 -48119
box -152 -44 30474 20044
use nfet$2  nfet$2_27
timestamp 1676577649
transform 1 0 82886 0 1 -48119
box -152 -44 30474 20044
use nfet$2  nfet$2_28
timestamp 1676577649
transform 1 0 50886 0 1 -48119
box -152 -44 30474 20044
use nfet$2  nfet$2_29
timestamp 1676577649
transform 1 0 18886 0 1 -48119
box -152 -44 30474 20044
use nfet$2  nfet$2_30
timestamp 1676577649
transform 1 0 -13114 0 1 -48119
box -152 -44 30474 20044
use nfet$2  nfet$2_31
timestamp 1676577649
transform 1 0 -45114 0 1 -48119
box -152 -44 30474 20044
use nfet$2  nfet$2_32
timestamp 1676577649
transform 1 0 -77114 0 1 -48119
box -152 -44 30474 20044
use nfet$2  nfet$2_33
timestamp 1676577649
transform 1 0 -109114 0 1 -48119
box -152 -44 30474 20044
use nfet$2  nfet$2_34
timestamp 1676577649
transform 1 0 146886 0 1 -74119
box -152 -44 30474 20044
use nfet$2  nfet$2_35
timestamp 1676577649
transform 1 0 114886 0 1 -74119
box -152 -44 30474 20044
use nfet$2  nfet$2_36
timestamp 1676577649
transform 1 0 82886 0 1 -74119
box -152 -44 30474 20044
use nfet$2  nfet$2_37
timestamp 1676577649
transform 1 0 50886 0 1 -74119
box -152 -44 30474 20044
use nfet$2  nfet$2_38
timestamp 1676577649
transform 1 0 18886 0 1 -74119
box -152 -44 30474 20044
use nfet$2  nfet$2_39
timestamp 1676577649
transform 1 0 -13114 0 1 -74119
box -152 -44 30474 20044
use nfet$2  nfet$2_40
timestamp 1676577649
transform 1 0 -45114 0 1 -74119
box -152 -44 30474 20044
use nfet$2  nfet$2_41
timestamp 1676577649
transform 1 0 -77114 0 1 -74119
box -152 -44 30474 20044
use nfet$2  nfet$2_42
timestamp 1676577649
transform 1 0 -109114 0 1 -74119
box -152 -44 30474 20044
use nfet$4  nfet$4_0
timestamp 1676577649
transform 1 0 -105662 0 1 -142783
box -152 -44 378 4044
use nfet  nfet_0
timestamp 1676577649
transform 1 0 -97974 0 1 -162683
box -152 -44 18314 12044
use pfet$2  pfet$2_0
timestamp 1676577649
transform 1 0 -6782 0 1 4066
box -176 -86 662 2086
use pfet$4  pfet$4_0
timestamp 1676577649
transform 1 0 85016 0 1 5307
box -176 -86 24558 20086
use pfet$4  pfet$4_1
timestamp 1676577649
transform 1 0 58016 0 1 5307
box -176 -86 24558 20086
use pfet$4  pfet$4_2
timestamp 1676577649
transform 1 0 85016 0 1 -19693
box -176 -86 24558 20086
use pfet$4  pfet$4_3
timestamp 1676577649
transform 1 0 58016 0 1 -19693
box -176 -86 24558 20086
use pfet  pfet_0
timestamp 1676577649
transform 1 0 27894 0 1 -46
box -176 -86 25358 10086
use pfet  pfet_1
timestamp 1676577649
transform 1 0 -106 0 1 -46
box -176 -86 25358 10086
<< labels >>
flabel metal1 s -128799 -36371 -128799 -36371 2 FreeSans 73 0 0 0 vin1
port 1 nsew
flabel metal1 s -29619 24412 -29619 24412 2 FreeSans 73 0 0 0 vp
port 2 nsew
flabel metal1 s 186234 -94324 186234 -94324 2 FreeSans 73 0 0 0 vin2
port 3 nsew
flabel metal1 s 175714 -18102 175714 -18102 2 FreeSans 73 0 0 0 vout
port 4 nsew
flabel metal1 s 3120 -173713 3120 -173713 2 FreeSans 73 0 0 0 vss
port 5 nsew
flabel metal1 s 12521 30597 12521 30597 2 FreeSans 73 0 0 0 vdd
port 6 nsew
flabel polysilicon s -94027 -145689 -94027 -145689 2 FreeSans 57 0 0 0 vbias_tail
flabel metal2 s 12340 -21248 12340 -21248 2 FreeSans 89 0 0 0 vx
port 7 nsew
flabel metal2 s -77010 -136039 -77010 -136039 2 FreeSans 89 0 0 0 vtail
port 8 nsew
<< properties >>
string FIXED_BBOX -14213 -14031 -5023 -6761
<< end >>
