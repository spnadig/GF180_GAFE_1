** sch_path: /usr/local/google/home/nigelcoburn/MixedSignal_ENV/GF180_GAFE_1/opamp_rewire.sch
.subckt OTA_2stage vdd vss vin1 vin2 vp vout
*.PININFO vdd:B vss:B vin1:I vin2:I vp:I vout:O
M1 vtail vin1 vx vss nfet_03v3 L=1u W=10000u nf=100 m=18
M2 vtail vin2 net1 vss nfet_03v3 L=1u W=10000u nf=100 m=18
M3 vdd vx vx vdd pfet_03v3 L=2u W=2500u nf=50 m=1
M4 vdd vx net1 vdd pfet_03v3 L=2u W=2500u nf=50 m=1
M5 vss vbias_tail vtail vss nfet_03v3 L=1u W=3600u nf=60 m=1
M6 vbias_tail vbias_tail vss vss nfet_03v3 L=1u W=20u nf=1 m=1
M7 vdd vp vbias_tail vdd pfet_03v3 L=2u W=10u nf=1 m=1
M8 vdd net1 vout vdd pfet_03v3 L=0.7u W=10000u nf=100 m=4
M9 vss vbias_tail vout vss nfet_03v3 L=1u W=10000u nf=100 m=7
C2 vout vss 1p m=1
C1 net2 vout 3p m=1
R1 net1 net2 200 m=1
.ends
.end
