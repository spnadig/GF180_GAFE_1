* Extracted by KLayout with GF180 LVS runset on : 08/02/2023 01:33

.SUBCKT TopLevel_oscillator
M$1 \$25 \$4 \$2 \$25 pfet_03v3_dn L=5U W=0.5U AS=0.22P AD=0.22P PS=1.88U
+ PD=1.88U
M$2 \$25 \$2 \$3 \$25 pfet_03v3_dn L=5U W=0.5U AS=0.22P AD=0.22P PS=1.88U
+ PD=1.88U
M$3 \$25 \$3 \$4 \$25 pfet_03v3_dn L=5U W=0.5U AS=0.22P AD=0.22P PS=1.88U
+ PD=1.88U
M$4 \$1 \$4 \$2 \$1 nfet_03v3_dn L=5U W=0.5U AS=0.22P AD=0.22P PS=1.88U PD=1.88U
M$5 \$1 \$2 \$3 \$1 nfet_03v3_dn L=5U W=0.5U AS=0.22P AD=0.22P PS=1.88U PD=1.88U
M$6 \$1 \$3 \$4 \$1 nfet_03v3_dn L=5U W=0.5U AS=0.22P AD=0.22P PS=1.88U PD=1.88U
.ENDS TopLevel_oscillator
