* NGSPICE file created from Inverter.ext - technology: gf180mcuC

.subckt Inverter VDD GND IN OUT
X0 OUT IN GND GND nmos_3p3 w=0.22u l=0.28u
X1 OUT IN VDD VDD pmos_3p3 w=0.22u l=0.28u
.ends
