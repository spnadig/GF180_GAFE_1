(*blackbox*)
module OTA_2stage_macro (
`ifdef USE_POWER_PINS
    inout vdd,
    inout vss,
`endif
);
endmodule // OTA_2stage
