VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OTA_2stage
  CLASS BLOCK ;
  FOREIGN OTA_2stage ;
  ORIGIN 71.065 70.155 ;
  SIZE 45.950 BY 36.350 ;
  PIN vin1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT -657.770 -190.455 -632.000 -176.505 ;
    END
  END vin1
  PIN vp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT -157.970 104.405 -118.000 135.960 ;
    END
  END vp
  PIN vin2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 917.630 -477.530 943.025 -460.295 ;
    END
  END vin2
  PIN vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 870.620 -104.375 890.710 -74.875 ;
    END
  END vout
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT -572.210 -882.355 408.135 -856.395 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT -0.540 53.390 125.840 161.245 ;
    END
  END vdd
  OBS
      LAYER Nwell ;
        RECT -34.790 19.900 -30.600 30.760 ;
        RECT -1.410 -0.660 126.260 50.200 ;
        RECT 138.590 -0.660 266.260 50.200 ;
        RECT 289.200 26.105 412.870 126.965 ;
        RECT 424.200 26.105 547.870 126.965 ;
        RECT -72.565 -71.655 -23.615 -32.305 ;
        RECT 289.200 -98.895 412.870 1.965 ;
        RECT 424.200 -98.895 547.870 1.965 ;
      LAYER Pwell ;
        RECT -548.990 -243.525 -390.280 -138.790 ;
        RECT -388.990 -243.525 -230.280 -138.790 ;
        RECT -228.990 -243.525 -70.280 -138.790 ;
        RECT -68.990 -243.525 89.720 -138.790 ;
        RECT 91.010 -243.525 249.720 -138.790 ;
        RECT 251.010 -243.525 409.720 -138.790 ;
        RECT 411.010 -243.525 569.720 -138.790 ;
        RECT 571.010 -243.525 729.720 -138.790 ;
        RECT 731.010 -243.525 889.720 -138.790 ;
        RECT -548.990 -373.525 -390.280 -268.790 ;
        RECT -388.990 -373.525 -230.280 -268.790 ;
        RECT -228.990 -373.525 -70.280 -268.790 ;
        RECT -68.990 -373.525 89.720 -268.790 ;
        RECT 91.010 -373.525 249.720 -268.790 ;
        RECT 251.010 -373.525 409.720 -268.790 ;
        RECT 411.010 -373.525 569.720 -268.790 ;
        RECT 571.010 -373.525 729.720 -268.790 ;
        RECT 731.010 -373.525 889.720 -268.790 ;
        RECT -548.990 -518.525 -390.280 -413.700 ;
        RECT -388.990 -518.525 -230.280 -413.700 ;
        RECT -228.990 -518.525 -70.280 -413.700 ;
        RECT -68.990 -518.525 89.720 -413.700 ;
        RECT 91.010 -518.525 249.720 -413.700 ;
        RECT 251.010 -518.525 409.720 -413.700 ;
        RECT 411.010 -518.525 569.720 -413.700 ;
        RECT 571.010 -518.525 729.720 -413.700 ;
        RECT 731.010 -518.525 889.720 -413.700 ;
        RECT -548.990 -648.525 -390.280 -543.750 ;
        RECT -388.990 -648.525 -230.280 -543.750 ;
        RECT -228.990 -648.525 -70.280 -543.750 ;
        RECT -68.990 -648.525 89.720 -543.750 ;
        RECT 91.010 -648.525 249.720 -543.750 ;
        RECT 251.010 -648.525 409.720 -543.750 ;
        RECT 411.010 -648.525 569.720 -543.750 ;
        RECT 571.010 -648.525 729.720 -543.750 ;
        RECT 731.010 -648.525 889.720 -543.750 ;
        RECT -531.730 -716.810 -523.500 -690.985 ;
        RECT -493.095 -815.165 -396.230 -751.120 ;
        RECT -303.900 -814.690 -145.190 -710.190 ;
        RECT -133.900 -814.690 24.810 -710.190 ;
        RECT 36.100 -814.690 194.810 -710.190 ;
        RECT 206.100 -814.690 364.810 -710.190 ;
        RECT 376.100 -814.690 534.810 -710.190 ;
        RECT 546.100 -814.690 704.810 -710.190 ;
        RECT 716.100 -814.690 874.810 -710.190 ;
      LAYER Metal1 ;
        RECT -67.740 145.550 -0.540 161.245 ;
        RECT 125.840 145.550 549.305 161.245 ;
        RECT -169.365 104.405 -157.970 135.960 ;
        RECT -150.690 13.275 -85.050 29.445 ;
        RECT -57.750 20.320 -33.540 145.550 ;
        RECT 139.460 53.390 265.840 145.550 ;
        RECT -0.540 49.770 -0.160 53.390 ;
        RECT -31.400 13.275 -26.845 30.340 ;
        RECT -150.690 4.390 -26.845 13.275 ;
        RECT -150.690 -1.315 -85.050 4.390 ;
        RECT -1.330 -0.240 -0.160 49.770 ;
        RECT 1.980 -3.850 2.360 49.780 ;
        RECT 4.500 -0.240 4.880 53.390 ;
        RECT 7.020 -3.850 7.400 49.780 ;
        RECT 9.540 -0.240 9.920 53.390 ;
        RECT 12.060 -3.850 12.440 49.780 ;
        RECT 14.580 -0.240 14.960 53.390 ;
        RECT 17.100 -3.850 17.480 49.780 ;
        RECT 19.620 -0.240 20.000 53.390 ;
        RECT 22.140 -3.850 22.520 49.780 ;
        RECT 24.660 -0.240 25.040 53.390 ;
        RECT 27.180 -3.850 27.560 49.780 ;
        RECT 29.700 -0.240 30.080 53.390 ;
        RECT 32.220 -3.850 32.600 49.780 ;
        RECT 34.740 -0.240 35.120 53.390 ;
        RECT 37.260 -3.850 37.640 49.780 ;
        RECT 39.780 -0.240 40.160 53.390 ;
        RECT 42.300 -3.850 42.680 49.780 ;
        RECT 44.820 -0.240 45.200 53.390 ;
        RECT 47.340 -3.850 47.720 49.780 ;
        RECT 49.860 -0.240 50.240 53.390 ;
        RECT 52.380 -3.850 52.760 49.780 ;
        RECT 54.900 -0.240 55.280 53.390 ;
        RECT 57.420 -3.850 57.800 49.780 ;
        RECT 59.940 -0.240 60.320 53.390 ;
        RECT 62.460 -3.850 62.840 49.780 ;
        RECT 64.980 -0.240 65.360 53.390 ;
        RECT 67.500 -3.850 67.880 49.780 ;
        RECT 70.020 -0.240 70.400 53.390 ;
        RECT 72.540 -3.850 72.920 49.780 ;
        RECT 75.060 -0.240 75.440 53.390 ;
        RECT 77.580 -3.850 77.960 49.780 ;
        RECT 80.100 -0.240 80.480 53.390 ;
        RECT 82.620 -3.850 83.000 49.780 ;
        RECT 85.140 -0.240 85.520 53.390 ;
        RECT 87.660 -3.850 88.040 49.780 ;
        RECT 90.180 -0.240 90.560 53.390 ;
        RECT 92.700 -3.850 93.080 49.780 ;
        RECT 95.220 -0.240 95.600 53.390 ;
        RECT 97.740 -3.850 98.120 49.780 ;
        RECT 100.260 -0.240 100.640 53.390 ;
        RECT 102.780 -3.850 103.160 49.780 ;
        RECT 105.300 -0.240 105.680 53.390 ;
        RECT 107.820 -3.850 108.200 49.780 ;
        RECT 110.340 -0.240 110.720 53.390 ;
        RECT 112.860 -3.850 113.240 49.780 ;
        RECT 115.380 -0.240 115.760 53.390 ;
        RECT 117.900 -3.850 118.280 49.780 ;
        RECT 120.420 -0.240 120.800 53.390 ;
        RECT 122.940 -3.850 123.320 49.780 ;
        RECT 125.460 -0.240 125.840 53.390 ;
        RECT 139.460 49.770 139.840 53.390 ;
        RECT 138.670 -0.240 139.840 49.770 ;
        RECT 141.980 -3.850 142.360 49.780 ;
        RECT 144.500 -0.240 144.880 53.390 ;
        RECT 147.020 -3.850 147.400 49.780 ;
        RECT 149.540 -0.240 149.920 53.390 ;
        RECT 152.060 -3.850 152.440 49.780 ;
        RECT 154.580 -0.240 154.960 53.390 ;
        RECT 157.100 -3.850 157.480 49.780 ;
        RECT 159.620 -0.240 160.000 53.390 ;
        RECT 162.140 -3.850 162.520 49.780 ;
        RECT 164.660 -0.240 165.040 53.390 ;
        RECT 167.180 -3.850 167.560 49.780 ;
        RECT 169.700 -0.240 170.080 53.390 ;
        RECT 172.220 -3.850 172.600 49.780 ;
        RECT 174.740 -0.240 175.120 53.390 ;
        RECT 177.260 -3.850 177.640 49.780 ;
        RECT 179.780 -0.240 180.160 53.390 ;
        RECT 182.300 -3.850 182.680 49.780 ;
        RECT 184.820 -0.240 185.200 53.390 ;
        RECT 187.340 -3.850 187.720 49.780 ;
        RECT 189.860 -0.240 190.240 53.390 ;
        RECT 192.380 -3.850 192.760 49.780 ;
        RECT 194.900 -0.240 195.280 53.390 ;
        RECT 197.420 -3.850 197.800 49.780 ;
        RECT 199.940 -0.240 200.320 53.390 ;
        RECT 202.460 -3.850 202.840 49.780 ;
        RECT 204.980 -0.240 205.360 53.390 ;
        RECT 207.500 -3.850 207.880 49.780 ;
        RECT 210.020 -0.240 210.400 53.390 ;
        RECT 212.540 -3.850 212.920 49.780 ;
        RECT 215.060 -0.240 215.440 53.390 ;
        RECT 217.580 -3.850 217.960 49.780 ;
        RECT 220.100 -0.240 220.480 53.390 ;
        RECT 222.620 -3.850 223.000 49.780 ;
        RECT 225.140 -0.240 225.520 53.390 ;
        RECT 227.660 -3.850 228.040 49.780 ;
        RECT 230.180 -0.240 230.560 53.390 ;
        RECT 232.700 -3.850 233.080 49.780 ;
        RECT 235.220 -0.240 235.600 53.390 ;
        RECT 237.740 -3.850 238.120 49.780 ;
        RECT 240.260 -0.240 240.640 53.390 ;
        RECT 242.780 -3.850 243.160 49.780 ;
        RECT 245.300 -0.240 245.680 53.390 ;
        RECT 247.820 -3.850 248.200 49.780 ;
        RECT 250.340 -0.240 250.720 53.390 ;
        RECT 252.860 -3.850 253.240 49.780 ;
        RECT 255.380 -0.240 255.760 53.390 ;
        RECT 257.900 -3.850 258.280 49.780 ;
        RECT 260.420 -0.240 260.800 53.390 ;
        RECT 262.940 -3.850 263.320 49.780 ;
        RECT 265.460 -0.240 265.840 53.390 ;
        RECT 282.460 128.970 547.450 145.550 ;
        RECT 268.360 -3.850 279.100 18.760 ;
        RECT -71.640 -70.730 -24.540 -33.230 ;
        RECT 1.980 -95.175 128.360 -3.850 ;
        RECT 141.980 -8.925 279.100 -3.850 ;
        RECT 282.460 7.445 290.450 128.970 ;
        RECT 291.290 24.100 291.670 126.545 ;
        RECT 292.510 26.525 292.890 128.970 ;
        RECT 293.730 24.100 294.110 126.545 ;
        RECT 294.950 26.525 295.330 128.970 ;
        RECT 296.170 24.100 296.550 126.545 ;
        RECT 297.390 26.525 297.770 128.970 ;
        RECT 298.610 24.100 298.990 126.545 ;
        RECT 299.830 26.525 300.210 128.970 ;
        RECT 301.050 24.100 301.430 126.545 ;
        RECT 302.270 26.525 302.650 128.970 ;
        RECT 303.490 24.100 303.870 126.545 ;
        RECT 304.710 26.525 305.090 128.970 ;
        RECT 305.930 24.100 306.310 126.545 ;
        RECT 307.150 26.525 307.530 128.970 ;
        RECT 308.370 24.100 308.750 126.545 ;
        RECT 309.590 26.525 309.970 128.970 ;
        RECT 310.810 24.100 311.190 126.545 ;
        RECT 312.030 26.525 312.410 128.970 ;
        RECT 313.250 24.100 313.630 126.545 ;
        RECT 314.470 26.525 314.850 128.970 ;
        RECT 315.690 24.100 316.070 126.545 ;
        RECT 316.910 26.525 317.290 128.970 ;
        RECT 318.130 24.100 318.510 126.545 ;
        RECT 319.350 26.525 319.730 128.970 ;
        RECT 320.570 24.100 320.950 126.545 ;
        RECT 321.790 26.525 322.170 128.970 ;
        RECT 323.010 24.100 323.390 126.545 ;
        RECT 324.230 26.525 324.610 128.970 ;
        RECT 325.450 24.100 325.830 126.545 ;
        RECT 326.670 26.525 327.050 128.970 ;
        RECT 327.890 24.100 328.270 126.545 ;
        RECT 329.110 26.525 329.490 128.970 ;
        RECT 330.330 24.100 330.710 126.545 ;
        RECT 331.550 26.525 331.930 128.970 ;
        RECT 332.770 24.100 333.150 126.545 ;
        RECT 333.990 26.525 334.370 128.970 ;
        RECT 335.210 24.100 335.590 126.545 ;
        RECT 336.430 26.525 336.810 128.970 ;
        RECT 337.650 24.100 338.030 126.545 ;
        RECT 338.870 26.525 339.250 128.970 ;
        RECT 340.090 24.100 340.470 126.545 ;
        RECT 341.310 26.525 341.690 128.970 ;
        RECT 342.530 24.100 342.910 126.545 ;
        RECT 343.750 26.525 344.130 128.970 ;
        RECT 344.970 24.100 345.350 126.545 ;
        RECT 346.190 26.525 346.570 128.970 ;
        RECT 347.410 24.100 347.790 126.545 ;
        RECT 348.630 26.525 349.010 128.970 ;
        RECT 349.850 24.100 350.230 126.545 ;
        RECT 351.070 26.525 351.450 128.970 ;
        RECT 352.290 24.100 352.670 126.545 ;
        RECT 353.510 26.525 353.890 128.970 ;
        RECT 354.730 24.100 355.110 126.545 ;
        RECT 355.950 26.525 356.330 128.970 ;
        RECT 357.170 24.100 357.550 126.545 ;
        RECT 358.390 26.525 358.770 128.970 ;
        RECT 359.610 24.100 359.990 126.545 ;
        RECT 360.830 26.525 361.210 128.970 ;
        RECT 362.050 24.100 362.430 126.545 ;
        RECT 363.270 26.525 363.650 128.970 ;
        RECT 364.490 24.100 364.870 126.545 ;
        RECT 365.710 26.525 366.090 128.970 ;
        RECT 366.930 24.100 367.310 126.545 ;
        RECT 368.150 26.525 368.530 128.970 ;
        RECT 369.370 24.100 369.750 126.545 ;
        RECT 370.590 26.525 370.970 128.970 ;
        RECT 371.810 24.100 372.190 126.545 ;
        RECT 373.030 26.525 373.410 128.970 ;
        RECT 374.250 24.100 374.630 126.545 ;
        RECT 375.470 26.525 375.850 128.970 ;
        RECT 376.690 24.100 377.070 126.545 ;
        RECT 377.910 26.525 378.290 128.970 ;
        RECT 379.130 24.100 379.510 126.545 ;
        RECT 380.350 26.525 380.730 128.970 ;
        RECT 381.570 24.100 381.950 126.545 ;
        RECT 382.790 26.525 383.170 128.970 ;
        RECT 384.010 24.100 384.390 126.545 ;
        RECT 385.230 26.525 385.610 128.970 ;
        RECT 386.450 24.100 386.830 126.545 ;
        RECT 387.670 26.525 388.050 128.970 ;
        RECT 388.890 24.100 389.270 126.545 ;
        RECT 390.110 26.525 390.490 128.970 ;
        RECT 391.330 24.100 391.710 126.545 ;
        RECT 392.550 26.525 392.930 128.970 ;
        RECT 393.770 24.100 394.150 126.545 ;
        RECT 394.990 26.525 395.370 128.970 ;
        RECT 396.210 24.100 396.590 126.545 ;
        RECT 397.430 26.525 397.810 128.970 ;
        RECT 398.650 24.100 399.030 126.545 ;
        RECT 399.870 26.525 400.250 128.970 ;
        RECT 401.090 24.100 401.470 126.545 ;
        RECT 402.310 26.525 402.690 128.970 ;
        RECT 403.530 24.100 403.910 126.545 ;
        RECT 404.750 26.525 405.130 128.970 ;
        RECT 405.970 24.100 406.350 126.545 ;
        RECT 407.190 26.525 407.570 128.970 ;
        RECT 408.410 24.100 408.790 126.545 ;
        RECT 409.630 26.525 410.010 128.970 ;
        RECT 410.850 24.100 411.230 126.545 ;
        RECT 412.070 26.525 412.450 128.970 ;
        RECT 425.070 126.535 425.450 128.970 ;
        RECT 424.280 26.525 425.450 126.535 ;
        RECT 426.290 24.100 426.670 126.545 ;
        RECT 427.510 26.525 427.890 128.970 ;
        RECT 428.730 24.100 429.110 126.545 ;
        RECT 429.950 26.525 430.330 128.970 ;
        RECT 431.170 24.100 431.550 126.545 ;
        RECT 432.390 26.525 432.770 128.970 ;
        RECT 433.610 24.100 433.990 126.545 ;
        RECT 434.830 26.525 435.210 128.970 ;
        RECT 436.050 24.100 436.430 126.545 ;
        RECT 437.270 26.525 437.650 128.970 ;
        RECT 438.490 24.100 438.870 126.545 ;
        RECT 439.710 26.525 440.090 128.970 ;
        RECT 440.930 24.100 441.310 126.545 ;
        RECT 442.150 26.525 442.530 128.970 ;
        RECT 443.370 24.100 443.750 126.545 ;
        RECT 444.590 26.525 444.970 128.970 ;
        RECT 445.810 24.100 446.190 126.545 ;
        RECT 447.030 26.525 447.410 128.970 ;
        RECT 448.250 24.100 448.630 126.545 ;
        RECT 449.470 26.525 449.850 128.970 ;
        RECT 450.690 24.100 451.070 126.545 ;
        RECT 451.910 26.525 452.290 128.970 ;
        RECT 453.130 24.100 453.510 126.545 ;
        RECT 454.350 26.525 454.730 128.970 ;
        RECT 455.570 24.100 455.950 126.545 ;
        RECT 456.790 26.525 457.170 128.970 ;
        RECT 458.010 24.100 458.390 126.545 ;
        RECT 459.230 26.525 459.610 128.970 ;
        RECT 460.450 24.100 460.830 126.545 ;
        RECT 461.670 26.525 462.050 128.970 ;
        RECT 462.890 24.100 463.270 126.545 ;
        RECT 464.110 26.525 464.490 128.970 ;
        RECT 465.330 24.100 465.710 126.545 ;
        RECT 466.550 26.525 466.930 128.970 ;
        RECT 467.770 24.100 468.150 126.545 ;
        RECT 468.990 26.525 469.370 128.970 ;
        RECT 470.210 24.100 470.590 126.545 ;
        RECT 471.430 26.525 471.810 128.970 ;
        RECT 472.650 24.100 473.030 126.545 ;
        RECT 473.870 26.525 474.250 128.970 ;
        RECT 475.090 24.100 475.470 126.545 ;
        RECT 476.310 26.525 476.690 128.970 ;
        RECT 477.530 24.100 477.910 126.545 ;
        RECT 478.750 26.525 479.130 128.970 ;
        RECT 479.970 24.100 480.350 126.545 ;
        RECT 481.190 26.525 481.570 128.970 ;
        RECT 482.410 24.100 482.790 126.545 ;
        RECT 483.630 26.525 484.010 128.970 ;
        RECT 484.850 24.100 485.230 126.545 ;
        RECT 486.070 26.525 486.450 128.970 ;
        RECT 487.290 24.100 487.670 126.545 ;
        RECT 488.510 26.525 488.890 128.970 ;
        RECT 489.730 24.100 490.110 126.545 ;
        RECT 490.950 26.525 491.330 128.970 ;
        RECT 492.170 24.100 492.550 126.545 ;
        RECT 493.390 26.525 493.770 128.970 ;
        RECT 494.610 24.100 494.990 126.545 ;
        RECT 495.830 26.525 496.210 128.970 ;
        RECT 497.050 24.100 497.430 126.545 ;
        RECT 498.270 26.525 498.650 128.970 ;
        RECT 499.490 24.100 499.870 126.545 ;
        RECT 500.710 26.525 501.090 128.970 ;
        RECT 501.930 24.100 502.310 126.545 ;
        RECT 503.150 26.525 503.530 128.970 ;
        RECT 504.370 24.100 504.750 126.545 ;
        RECT 505.590 26.525 505.970 128.970 ;
        RECT 506.810 24.100 507.190 126.545 ;
        RECT 508.030 26.525 508.410 128.970 ;
        RECT 509.250 24.100 509.630 126.545 ;
        RECT 510.470 26.525 510.850 128.970 ;
        RECT 511.690 24.100 512.070 126.545 ;
        RECT 512.910 26.525 513.290 128.970 ;
        RECT 514.130 24.100 514.510 126.545 ;
        RECT 515.350 26.525 515.730 128.970 ;
        RECT 516.570 24.100 516.950 126.545 ;
        RECT 517.790 26.525 518.170 128.970 ;
        RECT 519.010 24.100 519.390 126.545 ;
        RECT 520.230 26.525 520.610 128.970 ;
        RECT 521.450 24.100 521.830 126.545 ;
        RECT 522.670 26.525 523.050 128.970 ;
        RECT 523.890 24.100 524.270 126.545 ;
        RECT 525.110 26.525 525.490 128.970 ;
        RECT 526.330 24.100 526.710 126.545 ;
        RECT 527.550 26.525 527.930 128.970 ;
        RECT 528.770 24.100 529.150 126.545 ;
        RECT 529.990 26.525 530.370 128.970 ;
        RECT 531.210 24.100 531.590 126.545 ;
        RECT 532.430 26.525 532.810 128.970 ;
        RECT 533.650 24.100 534.030 126.545 ;
        RECT 534.870 26.525 535.250 128.970 ;
        RECT 536.090 24.100 536.470 126.545 ;
        RECT 537.310 26.525 537.690 128.970 ;
        RECT 538.530 24.100 538.910 126.545 ;
        RECT 539.750 26.525 540.130 128.970 ;
        RECT 540.970 24.100 541.350 126.545 ;
        RECT 542.190 26.525 542.570 128.970 ;
        RECT 543.410 24.100 543.790 126.545 ;
        RECT 544.630 26.525 545.010 128.970 ;
        RECT 545.850 24.100 546.230 126.545 ;
        RECT 547.070 26.525 547.450 128.970 ;
        RECT 291.290 20.625 558.230 24.100 ;
        RECT 282.460 3.970 547.450 7.445 ;
        RECT 171.035 -95.645 254.970 -8.925 ;
        RECT 282.460 -98.475 290.450 3.970 ;
        RECT 291.290 -100.900 291.670 1.545 ;
        RECT 292.510 -98.475 292.890 3.970 ;
        RECT 293.730 -100.900 294.110 1.545 ;
        RECT 294.950 -98.475 295.330 3.970 ;
        RECT 296.170 -100.900 296.550 1.545 ;
        RECT 297.390 -98.475 297.770 3.970 ;
        RECT 298.610 -100.900 298.990 1.545 ;
        RECT 299.830 -98.475 300.210 3.970 ;
        RECT 301.050 -100.900 301.430 1.545 ;
        RECT 302.270 -98.475 302.650 3.970 ;
        RECT 303.490 -100.900 303.870 1.545 ;
        RECT 304.710 -98.475 305.090 3.970 ;
        RECT 305.930 -100.900 306.310 1.545 ;
        RECT 307.150 -98.475 307.530 3.970 ;
        RECT 308.370 -100.900 308.750 1.545 ;
        RECT 309.590 -98.475 309.970 3.970 ;
        RECT 310.810 -100.900 311.190 1.545 ;
        RECT 312.030 -98.475 312.410 3.970 ;
        RECT 313.250 -100.900 313.630 1.545 ;
        RECT 314.470 -98.475 314.850 3.970 ;
        RECT 315.690 -100.900 316.070 1.545 ;
        RECT 316.910 -98.475 317.290 3.970 ;
        RECT 318.130 -100.900 318.510 1.545 ;
        RECT 319.350 -98.475 319.730 3.970 ;
        RECT 320.570 -100.900 320.950 1.545 ;
        RECT 321.790 -98.475 322.170 3.970 ;
        RECT 323.010 -100.900 323.390 1.545 ;
        RECT 324.230 -98.475 324.610 3.970 ;
        RECT 325.450 -100.900 325.830 1.545 ;
        RECT 326.670 -98.475 327.050 3.970 ;
        RECT 327.890 -100.900 328.270 1.545 ;
        RECT 329.110 -98.475 329.490 3.970 ;
        RECT 330.330 -100.900 330.710 1.545 ;
        RECT 331.550 -98.475 331.930 3.970 ;
        RECT 332.770 -100.900 333.150 1.545 ;
        RECT 333.990 -98.475 334.370 3.970 ;
        RECT 335.210 -100.900 335.590 1.545 ;
        RECT 336.430 -98.475 336.810 3.970 ;
        RECT 337.650 -100.900 338.030 1.545 ;
        RECT 338.870 -98.475 339.250 3.970 ;
        RECT 340.090 -100.900 340.470 1.545 ;
        RECT 341.310 -98.475 341.690 3.970 ;
        RECT 342.530 -100.900 342.910 1.545 ;
        RECT 343.750 -98.475 344.130 3.970 ;
        RECT 344.970 -100.900 345.350 1.545 ;
        RECT 346.190 -98.475 346.570 3.970 ;
        RECT 347.410 -100.900 347.790 1.545 ;
        RECT 348.630 -98.475 349.010 3.970 ;
        RECT 349.850 -100.900 350.230 1.545 ;
        RECT 351.070 -98.475 351.450 3.970 ;
        RECT 352.290 -100.900 352.670 1.545 ;
        RECT 353.510 -98.475 353.890 3.970 ;
        RECT 354.730 -100.900 355.110 1.545 ;
        RECT 355.950 -98.475 356.330 3.970 ;
        RECT 357.170 -100.900 357.550 1.545 ;
        RECT 358.390 -98.475 358.770 3.970 ;
        RECT 359.610 -100.900 359.990 1.545 ;
        RECT 360.830 -98.475 361.210 3.970 ;
        RECT 362.050 -100.900 362.430 1.545 ;
        RECT 363.270 -98.475 363.650 3.970 ;
        RECT 364.490 -100.900 364.870 1.545 ;
        RECT 365.710 -98.475 366.090 3.970 ;
        RECT 366.930 -100.900 367.310 1.545 ;
        RECT 368.150 -98.475 368.530 3.970 ;
        RECT 369.370 -100.900 369.750 1.545 ;
        RECT 370.590 -98.475 370.970 3.970 ;
        RECT 371.810 -100.900 372.190 1.545 ;
        RECT 373.030 -98.475 373.410 3.970 ;
        RECT 374.250 -100.900 374.630 1.545 ;
        RECT 375.470 -98.475 375.850 3.970 ;
        RECT 376.690 -100.900 377.070 1.545 ;
        RECT 377.910 -98.475 378.290 3.970 ;
        RECT 379.130 -100.900 379.510 1.545 ;
        RECT 380.350 -98.475 380.730 3.970 ;
        RECT 381.570 -100.900 381.950 1.545 ;
        RECT 382.790 -98.475 383.170 3.970 ;
        RECT 384.010 -100.900 384.390 1.545 ;
        RECT 385.230 -98.475 385.610 3.970 ;
        RECT 386.450 -100.900 386.830 1.545 ;
        RECT 387.670 -98.475 388.050 3.970 ;
        RECT 388.890 -100.900 389.270 1.545 ;
        RECT 390.110 -98.475 390.490 3.970 ;
        RECT 391.330 -100.900 391.710 1.545 ;
        RECT 392.550 -98.475 392.930 3.970 ;
        RECT 393.770 -100.900 394.150 1.545 ;
        RECT 394.990 -98.475 395.370 3.970 ;
        RECT 396.210 -100.900 396.590 1.545 ;
        RECT 397.430 -98.475 397.810 3.970 ;
        RECT 398.650 -100.900 399.030 1.545 ;
        RECT 399.870 -98.475 400.250 3.970 ;
        RECT 401.090 -100.900 401.470 1.545 ;
        RECT 402.310 -98.475 402.690 3.970 ;
        RECT 403.530 -100.900 403.910 1.545 ;
        RECT 404.750 -98.475 405.130 3.970 ;
        RECT 405.970 -100.900 406.350 1.545 ;
        RECT 407.190 -98.475 407.570 3.970 ;
        RECT 408.410 -100.900 408.790 1.545 ;
        RECT 409.630 -98.475 410.010 3.970 ;
        RECT 410.850 -100.900 411.230 1.545 ;
        RECT 412.070 -98.475 412.450 3.970 ;
        RECT 425.070 1.535 425.450 3.970 ;
        RECT 424.280 -98.475 425.450 1.535 ;
        RECT 426.290 -100.900 426.670 1.545 ;
        RECT 427.510 -98.475 427.890 3.970 ;
        RECT 428.730 -100.900 429.110 1.545 ;
        RECT 429.950 -98.475 430.330 3.970 ;
        RECT 431.170 -100.900 431.550 1.545 ;
        RECT 432.390 -98.475 432.770 3.970 ;
        RECT 433.610 -100.900 433.990 1.545 ;
        RECT 434.830 -98.475 435.210 3.970 ;
        RECT 436.050 -100.900 436.430 1.545 ;
        RECT 437.270 -98.475 437.650 3.970 ;
        RECT 438.490 -100.900 438.870 1.545 ;
        RECT 439.710 -98.475 440.090 3.970 ;
        RECT 440.930 -100.900 441.310 1.545 ;
        RECT 442.150 -98.475 442.530 3.970 ;
        RECT 443.370 -100.900 443.750 1.545 ;
        RECT 444.590 -98.475 444.970 3.970 ;
        RECT 445.810 -100.900 446.190 1.545 ;
        RECT 447.030 -98.475 447.410 3.970 ;
        RECT 448.250 -100.900 448.630 1.545 ;
        RECT 449.470 -98.475 449.850 3.970 ;
        RECT 450.690 -100.900 451.070 1.545 ;
        RECT 451.910 -98.475 452.290 3.970 ;
        RECT 453.130 -100.900 453.510 1.545 ;
        RECT 454.350 -98.475 454.730 3.970 ;
        RECT 455.570 -100.900 455.950 1.545 ;
        RECT 456.790 -98.475 457.170 3.970 ;
        RECT 458.010 -100.900 458.390 1.545 ;
        RECT 459.230 -98.475 459.610 3.970 ;
        RECT 460.450 -100.900 460.830 1.545 ;
        RECT 461.670 -98.475 462.050 3.970 ;
        RECT 462.890 -100.900 463.270 1.545 ;
        RECT 464.110 -98.475 464.490 3.970 ;
        RECT 465.330 -100.900 465.710 1.545 ;
        RECT 466.550 -98.475 466.930 3.970 ;
        RECT 467.770 -100.900 468.150 1.545 ;
        RECT 468.990 -98.475 469.370 3.970 ;
        RECT 470.210 -100.900 470.590 1.545 ;
        RECT 471.430 -98.475 471.810 3.970 ;
        RECT 472.650 -100.900 473.030 1.545 ;
        RECT 473.870 -98.475 474.250 3.970 ;
        RECT 475.090 -100.900 475.470 1.545 ;
        RECT 476.310 -98.475 476.690 3.970 ;
        RECT 477.530 -100.900 477.910 1.545 ;
        RECT 478.750 -98.475 479.130 3.970 ;
        RECT 479.970 -100.900 480.350 1.545 ;
        RECT 481.190 -98.475 481.570 3.970 ;
        RECT 482.410 -100.900 482.790 1.545 ;
        RECT 483.630 -98.475 484.010 3.970 ;
        RECT 484.850 -100.900 485.230 1.545 ;
        RECT 486.070 -98.475 486.450 3.970 ;
        RECT 487.290 -100.900 487.670 1.545 ;
        RECT 488.510 -98.475 488.890 3.970 ;
        RECT 489.730 -100.900 490.110 1.545 ;
        RECT 490.950 -98.475 491.330 3.970 ;
        RECT 492.170 -100.900 492.550 1.545 ;
        RECT 493.390 -98.475 493.770 3.970 ;
        RECT 494.610 -100.900 494.990 1.545 ;
        RECT 495.830 -98.475 496.210 3.970 ;
        RECT 497.050 -100.900 497.430 1.545 ;
        RECT 498.270 -98.475 498.650 3.970 ;
        RECT 499.490 -100.900 499.870 1.545 ;
        RECT 500.710 -98.475 501.090 3.970 ;
        RECT 501.930 -100.900 502.310 1.545 ;
        RECT 503.150 -98.475 503.530 3.970 ;
        RECT 504.370 -100.900 504.750 1.545 ;
        RECT 505.590 -98.475 505.970 3.970 ;
        RECT 506.810 -100.900 507.190 1.545 ;
        RECT 508.030 -98.475 508.410 3.970 ;
        RECT 509.250 -100.900 509.630 1.545 ;
        RECT 510.470 -98.475 510.850 3.970 ;
        RECT 511.690 -100.900 512.070 1.545 ;
        RECT 512.910 -98.475 513.290 3.970 ;
        RECT 514.130 -100.900 514.510 1.545 ;
        RECT 515.350 -98.475 515.730 3.970 ;
        RECT 516.570 -100.900 516.950 1.545 ;
        RECT 517.790 -98.475 518.170 3.970 ;
        RECT 519.010 -100.900 519.390 1.545 ;
        RECT 520.230 -98.475 520.610 3.970 ;
        RECT 521.450 -100.900 521.830 1.545 ;
        RECT 522.670 -98.475 523.050 3.970 ;
        RECT 523.890 -100.900 524.270 1.545 ;
        RECT 525.110 -98.475 525.490 3.970 ;
        RECT 526.330 -100.900 526.710 1.545 ;
        RECT 527.550 -98.475 527.930 3.970 ;
        RECT 528.770 -100.900 529.150 1.545 ;
        RECT 529.990 -98.475 530.370 3.970 ;
        RECT 531.210 -100.900 531.590 1.545 ;
        RECT 532.430 -98.475 532.810 3.970 ;
        RECT 533.650 -100.900 534.030 1.545 ;
        RECT 534.870 -98.475 535.250 3.970 ;
        RECT 536.090 -100.900 536.470 1.545 ;
        RECT 537.310 -98.475 537.690 3.970 ;
        RECT 538.530 -100.900 538.910 1.545 ;
        RECT 539.750 -98.475 540.130 3.970 ;
        RECT 540.970 -100.900 541.350 1.545 ;
        RECT 542.190 -98.475 542.570 3.970 ;
        RECT 543.410 -100.900 543.790 1.545 ;
        RECT 544.630 -98.475 545.010 3.970 ;
        RECT 545.850 -100.900 546.230 1.545 ;
        RECT 547.070 -98.475 547.450 3.970 ;
        RECT 548.670 -74.875 558.230 20.625 ;
        RECT 548.670 -100.900 870.620 -74.875 ;
        RECT 291.290 -104.375 870.620 -100.900 ;
        RECT -545.580 -136.015 886.800 -115.075 ;
        RECT -657.770 -176.505 -632.000 -160.025 ;
        RECT -572.210 -240.595 -545.890 -140.595 ;
        RECT -572.210 -270.595 -545.930 -240.595 ;
        RECT -545.580 -240.605 -545.200 -136.015 ;
        RECT -544.060 -245.175 -543.680 -140.585 ;
        RECT -542.540 -240.605 -542.160 -136.015 ;
        RECT -541.020 -245.175 -540.640 -140.585 ;
        RECT -539.500 -240.605 -539.120 -136.015 ;
        RECT -537.980 -245.175 -537.600 -140.585 ;
        RECT -536.460 -240.605 -536.080 -136.015 ;
        RECT -534.940 -245.175 -534.560 -140.585 ;
        RECT -533.420 -240.605 -533.040 -136.015 ;
        RECT -531.900 -245.175 -531.520 -140.585 ;
        RECT -530.380 -240.605 -530.000 -136.015 ;
        RECT -528.860 -245.175 -528.480 -140.585 ;
        RECT -527.340 -240.605 -526.960 -136.015 ;
        RECT -525.820 -245.175 -525.440 -140.585 ;
        RECT -524.300 -240.605 -523.920 -136.015 ;
        RECT -522.780 -245.175 -522.400 -140.585 ;
        RECT -521.260 -240.605 -520.880 -136.015 ;
        RECT -519.740 -245.175 -519.360 -140.585 ;
        RECT -518.220 -240.605 -517.840 -136.015 ;
        RECT -516.700 -245.175 -516.320 -140.585 ;
        RECT -515.180 -240.605 -514.800 -136.015 ;
        RECT -513.660 -245.175 -513.280 -140.585 ;
        RECT -512.140 -240.605 -511.760 -136.015 ;
        RECT -510.620 -245.175 -510.240 -140.585 ;
        RECT -509.100 -240.605 -508.720 -136.015 ;
        RECT -507.580 -245.175 -507.200 -140.585 ;
        RECT -506.060 -240.605 -505.680 -136.015 ;
        RECT -504.540 -245.175 -504.160 -140.585 ;
        RECT -503.020 -240.605 -502.640 -136.015 ;
        RECT -501.500 -245.175 -501.120 -140.585 ;
        RECT -499.980 -240.605 -499.600 -136.015 ;
        RECT -498.460 -245.175 -498.080 -140.585 ;
        RECT -496.940 -240.605 -496.560 -136.015 ;
        RECT -495.420 -245.175 -495.040 -140.585 ;
        RECT -493.900 -240.605 -493.520 -136.015 ;
        RECT -492.380 -245.175 -492.000 -140.585 ;
        RECT -490.860 -240.605 -490.480 -136.015 ;
        RECT -489.340 -245.175 -488.960 -140.585 ;
        RECT -487.820 -240.605 -487.440 -136.015 ;
        RECT -486.300 -245.175 -485.920 -140.585 ;
        RECT -484.780 -240.605 -484.400 -136.015 ;
        RECT -483.260 -245.175 -482.880 -140.585 ;
        RECT -481.740 -240.605 -481.360 -136.015 ;
        RECT -480.220 -245.175 -479.840 -140.585 ;
        RECT -478.700 -240.605 -478.320 -136.015 ;
        RECT -477.180 -245.175 -476.800 -140.585 ;
        RECT -475.660 -240.605 -475.280 -136.015 ;
        RECT -474.140 -245.175 -473.760 -140.585 ;
        RECT -472.620 -240.605 -472.240 -136.015 ;
        RECT -471.100 -245.175 -470.720 -140.585 ;
        RECT -469.580 -240.605 -469.200 -136.015 ;
        RECT -468.060 -245.175 -467.680 -140.585 ;
        RECT -466.540 -240.605 -466.160 -136.015 ;
        RECT -465.020 -245.175 -464.640 -140.585 ;
        RECT -463.500 -240.605 -463.120 -136.015 ;
        RECT -461.980 -245.175 -461.600 -140.585 ;
        RECT -460.460 -240.605 -460.080 -136.015 ;
        RECT -458.940 -245.175 -458.560 -140.585 ;
        RECT -457.420 -240.605 -457.040 -136.015 ;
        RECT -455.900 -245.175 -455.520 -140.585 ;
        RECT -454.380 -240.605 -454.000 -136.015 ;
        RECT -452.860 -245.175 -452.480 -140.585 ;
        RECT -451.340 -240.605 -450.960 -136.015 ;
        RECT -449.820 -245.175 -449.440 -140.585 ;
        RECT -448.300 -240.605 -447.920 -136.015 ;
        RECT -446.780 -245.175 -446.400 -140.585 ;
        RECT -445.260 -240.605 -444.880 -136.015 ;
        RECT -443.740 -245.175 -443.360 -140.585 ;
        RECT -442.220 -240.605 -441.840 -136.015 ;
        RECT -440.700 -245.175 -440.320 -140.585 ;
        RECT -439.180 -240.605 -438.800 -136.015 ;
        RECT -437.660 -245.175 -437.280 -140.585 ;
        RECT -436.140 -240.605 -435.760 -136.015 ;
        RECT -434.620 -245.175 -434.240 -140.585 ;
        RECT -433.100 -240.605 -432.720 -136.015 ;
        RECT -431.580 -245.175 -431.200 -140.585 ;
        RECT -430.060 -240.605 -429.680 -136.015 ;
        RECT -428.540 -245.175 -428.160 -140.585 ;
        RECT -427.020 -240.605 -426.640 -136.015 ;
        RECT -425.500 -245.175 -425.120 -140.585 ;
        RECT -423.980 -240.605 -423.600 -136.015 ;
        RECT -422.460 -245.175 -422.080 -140.585 ;
        RECT -420.940 -240.605 -420.560 -136.015 ;
        RECT -419.420 -245.175 -419.040 -140.585 ;
        RECT -417.900 -240.605 -417.520 -136.015 ;
        RECT -416.380 -245.175 -416.000 -140.585 ;
        RECT -414.860 -240.605 -414.480 -136.015 ;
        RECT -413.340 -245.175 -412.960 -140.585 ;
        RECT -411.820 -240.605 -411.440 -136.015 ;
        RECT -410.300 -245.175 -409.920 -140.585 ;
        RECT -408.780 -240.605 -408.400 -136.015 ;
        RECT -407.260 -245.175 -406.880 -140.585 ;
        RECT -405.740 -240.605 -405.360 -136.015 ;
        RECT -404.220 -245.175 -403.840 -140.585 ;
        RECT -402.700 -240.605 -402.320 -136.015 ;
        RECT -401.180 -245.175 -400.800 -140.585 ;
        RECT -399.660 -240.605 -399.280 -136.015 ;
        RECT -398.140 -245.175 -397.760 -140.585 ;
        RECT -396.620 -240.605 -396.240 -136.015 ;
        RECT -395.100 -245.175 -394.720 -140.585 ;
        RECT -393.580 -240.605 -393.200 -136.015 ;
        RECT -385.580 -140.595 -385.200 -136.015 ;
        RECT -386.370 -240.605 -385.200 -140.595 ;
        RECT -384.060 -245.175 -383.680 -140.585 ;
        RECT -382.540 -240.605 -382.160 -136.015 ;
        RECT -381.020 -245.175 -380.640 -140.585 ;
        RECT -379.500 -240.605 -379.120 -136.015 ;
        RECT -377.980 -245.175 -377.600 -140.585 ;
        RECT -376.460 -240.605 -376.080 -136.015 ;
        RECT -374.940 -245.175 -374.560 -140.585 ;
        RECT -373.420 -240.605 -373.040 -136.015 ;
        RECT -371.900 -245.175 -371.520 -140.585 ;
        RECT -370.380 -240.605 -370.000 -136.015 ;
        RECT -368.860 -245.175 -368.480 -140.585 ;
        RECT -367.340 -240.605 -366.960 -136.015 ;
        RECT -365.820 -245.175 -365.440 -140.585 ;
        RECT -364.300 -240.605 -363.920 -136.015 ;
        RECT -362.780 -245.175 -362.400 -140.585 ;
        RECT -361.260 -240.605 -360.880 -136.015 ;
        RECT -359.740 -245.175 -359.360 -140.585 ;
        RECT -358.220 -240.605 -357.840 -136.015 ;
        RECT -356.700 -245.175 -356.320 -140.585 ;
        RECT -355.180 -240.605 -354.800 -136.015 ;
        RECT -353.660 -245.175 -353.280 -140.585 ;
        RECT -352.140 -240.605 -351.760 -136.015 ;
        RECT -350.620 -245.175 -350.240 -140.585 ;
        RECT -349.100 -240.605 -348.720 -136.015 ;
        RECT -347.580 -245.175 -347.200 -140.585 ;
        RECT -346.060 -240.605 -345.680 -136.015 ;
        RECT -344.540 -245.175 -344.160 -140.585 ;
        RECT -343.020 -240.605 -342.640 -136.015 ;
        RECT -341.500 -245.175 -341.120 -140.585 ;
        RECT -339.980 -240.605 -339.600 -136.015 ;
        RECT -338.460 -245.175 -338.080 -140.585 ;
        RECT -336.940 -240.605 -336.560 -136.015 ;
        RECT -335.420 -245.175 -335.040 -140.585 ;
        RECT -333.900 -240.605 -333.520 -136.015 ;
        RECT -332.380 -245.175 -332.000 -140.585 ;
        RECT -330.860 -240.605 -330.480 -136.015 ;
        RECT -329.340 -245.175 -328.960 -140.585 ;
        RECT -327.820 -240.605 -327.440 -136.015 ;
        RECT -326.300 -245.175 -325.920 -140.585 ;
        RECT -324.780 -240.605 -324.400 -136.015 ;
        RECT -323.260 -245.175 -322.880 -140.585 ;
        RECT -321.740 -240.605 -321.360 -136.015 ;
        RECT -320.220 -245.175 -319.840 -140.585 ;
        RECT -318.700 -240.605 -318.320 -136.015 ;
        RECT -317.180 -245.175 -316.800 -140.585 ;
        RECT -315.660 -240.605 -315.280 -136.015 ;
        RECT -314.140 -245.175 -313.760 -140.585 ;
        RECT -312.620 -240.605 -312.240 -136.015 ;
        RECT -311.100 -245.175 -310.720 -140.585 ;
        RECT -309.580 -240.605 -309.200 -136.015 ;
        RECT -308.060 -245.175 -307.680 -140.585 ;
        RECT -306.540 -240.605 -306.160 -136.015 ;
        RECT -305.020 -245.175 -304.640 -140.585 ;
        RECT -303.500 -240.605 -303.120 -136.015 ;
        RECT -301.980 -245.175 -301.600 -140.585 ;
        RECT -300.460 -240.605 -300.080 -136.015 ;
        RECT -298.940 -245.175 -298.560 -140.585 ;
        RECT -297.420 -240.605 -297.040 -136.015 ;
        RECT -295.900 -245.175 -295.520 -140.585 ;
        RECT -294.380 -240.605 -294.000 -136.015 ;
        RECT -292.860 -245.175 -292.480 -140.585 ;
        RECT -291.340 -240.605 -290.960 -136.015 ;
        RECT -289.820 -245.175 -289.440 -140.585 ;
        RECT -288.300 -240.605 -287.920 -136.015 ;
        RECT -286.780 -245.175 -286.400 -140.585 ;
        RECT -285.260 -240.605 -284.880 -136.015 ;
        RECT -283.740 -245.175 -283.360 -140.585 ;
        RECT -282.220 -240.605 -281.840 -136.015 ;
        RECT -280.700 -245.175 -280.320 -140.585 ;
        RECT -279.180 -240.605 -278.800 -136.015 ;
        RECT -277.660 -245.175 -277.280 -140.585 ;
        RECT -276.140 -240.605 -275.760 -136.015 ;
        RECT -274.620 -245.175 -274.240 -140.585 ;
        RECT -273.100 -240.605 -272.720 -136.015 ;
        RECT -271.580 -245.175 -271.200 -140.585 ;
        RECT -270.060 -240.605 -269.680 -136.015 ;
        RECT -268.540 -245.175 -268.160 -140.585 ;
        RECT -267.020 -240.605 -266.640 -136.015 ;
        RECT -265.500 -245.175 -265.120 -140.585 ;
        RECT -263.980 -240.605 -263.600 -136.015 ;
        RECT -262.460 -245.175 -262.080 -140.585 ;
        RECT -260.940 -240.605 -260.560 -136.015 ;
        RECT -259.420 -245.175 -259.040 -140.585 ;
        RECT -257.900 -240.605 -257.520 -136.015 ;
        RECT -256.380 -245.175 -256.000 -140.585 ;
        RECT -254.860 -240.605 -254.480 -136.015 ;
        RECT -253.340 -245.175 -252.960 -140.585 ;
        RECT -251.820 -240.605 -251.440 -136.015 ;
        RECT -250.300 -245.175 -249.920 -140.585 ;
        RECT -248.780 -240.605 -248.400 -136.015 ;
        RECT -247.260 -245.175 -246.880 -140.585 ;
        RECT -245.740 -240.605 -245.360 -136.015 ;
        RECT -244.220 -245.175 -243.840 -140.585 ;
        RECT -242.700 -240.605 -242.320 -136.015 ;
        RECT -241.180 -245.175 -240.800 -140.585 ;
        RECT -239.660 -240.605 -239.280 -136.015 ;
        RECT -238.140 -245.175 -237.760 -140.585 ;
        RECT -236.620 -240.605 -236.240 -136.015 ;
        RECT -235.100 -245.175 -234.720 -140.585 ;
        RECT -233.580 -240.605 -233.200 -136.015 ;
        RECT -225.580 -140.595 -225.200 -136.015 ;
        RECT -226.370 -240.605 -225.200 -140.595 ;
        RECT -224.060 -245.175 -223.680 -140.585 ;
        RECT -222.540 -240.605 -222.160 -136.015 ;
        RECT -221.020 -245.175 -220.640 -140.585 ;
        RECT -219.500 -240.605 -219.120 -136.015 ;
        RECT -217.980 -245.175 -217.600 -140.585 ;
        RECT -216.460 -240.605 -216.080 -136.015 ;
        RECT -214.940 -245.175 -214.560 -140.585 ;
        RECT -213.420 -240.605 -213.040 -136.015 ;
        RECT -211.900 -245.175 -211.520 -140.585 ;
        RECT -210.380 -240.605 -210.000 -136.015 ;
        RECT -208.860 -245.175 -208.480 -140.585 ;
        RECT -207.340 -240.605 -206.960 -136.015 ;
        RECT -205.820 -245.175 -205.440 -140.585 ;
        RECT -204.300 -240.605 -203.920 -136.015 ;
        RECT -202.780 -245.175 -202.400 -140.585 ;
        RECT -201.260 -240.605 -200.880 -136.015 ;
        RECT -199.740 -245.175 -199.360 -140.585 ;
        RECT -198.220 -240.605 -197.840 -136.015 ;
        RECT -196.700 -245.175 -196.320 -140.585 ;
        RECT -195.180 -240.605 -194.800 -136.015 ;
        RECT -193.660 -245.175 -193.280 -140.585 ;
        RECT -192.140 -240.605 -191.760 -136.015 ;
        RECT -190.620 -245.175 -190.240 -140.585 ;
        RECT -189.100 -240.605 -188.720 -136.015 ;
        RECT -187.580 -245.175 -187.200 -140.585 ;
        RECT -186.060 -240.605 -185.680 -136.015 ;
        RECT -184.540 -245.175 -184.160 -140.585 ;
        RECT -183.020 -240.605 -182.640 -136.015 ;
        RECT -181.500 -245.175 -181.120 -140.585 ;
        RECT -179.980 -240.605 -179.600 -136.015 ;
        RECT -178.460 -245.175 -178.080 -140.585 ;
        RECT -176.940 -240.605 -176.560 -136.015 ;
        RECT -175.420 -245.175 -175.040 -140.585 ;
        RECT -173.900 -240.605 -173.520 -136.015 ;
        RECT -172.380 -245.175 -172.000 -140.585 ;
        RECT -170.860 -240.605 -170.480 -136.015 ;
        RECT -169.340 -245.175 -168.960 -140.585 ;
        RECT -167.820 -240.605 -167.440 -136.015 ;
        RECT -166.300 -245.175 -165.920 -140.585 ;
        RECT -164.780 -240.605 -164.400 -136.015 ;
        RECT -163.260 -245.175 -162.880 -140.585 ;
        RECT -161.740 -240.605 -161.360 -136.015 ;
        RECT -160.220 -245.175 -159.840 -140.585 ;
        RECT -158.700 -240.605 -158.320 -136.015 ;
        RECT -157.180 -245.175 -156.800 -140.585 ;
        RECT -155.660 -240.605 -155.280 -136.015 ;
        RECT -154.140 -245.175 -153.760 -140.585 ;
        RECT -152.620 -240.605 -152.240 -136.015 ;
        RECT -151.100 -245.175 -150.720 -140.585 ;
        RECT -149.580 -240.605 -149.200 -136.015 ;
        RECT -148.060 -245.175 -147.680 -140.585 ;
        RECT -146.540 -240.605 -146.160 -136.015 ;
        RECT -145.020 -245.175 -144.640 -140.585 ;
        RECT -143.500 -240.605 -143.120 -136.015 ;
        RECT -141.980 -245.175 -141.600 -140.585 ;
        RECT -140.460 -240.605 -140.080 -136.015 ;
        RECT -138.940 -245.175 -138.560 -140.585 ;
        RECT -137.420 -240.605 -137.040 -136.015 ;
        RECT -135.900 -245.175 -135.520 -140.585 ;
        RECT -134.380 -240.605 -134.000 -136.015 ;
        RECT -132.860 -245.175 -132.480 -140.585 ;
        RECT -131.340 -240.605 -130.960 -136.015 ;
        RECT -129.820 -245.175 -129.440 -140.585 ;
        RECT -128.300 -240.605 -127.920 -136.015 ;
        RECT -126.780 -245.175 -126.400 -140.585 ;
        RECT -125.260 -240.605 -124.880 -136.015 ;
        RECT -123.740 -245.175 -123.360 -140.585 ;
        RECT -122.220 -240.605 -121.840 -136.015 ;
        RECT -120.700 -245.175 -120.320 -140.585 ;
        RECT -119.180 -240.605 -118.800 -136.015 ;
        RECT -117.660 -245.175 -117.280 -140.585 ;
        RECT -116.140 -240.605 -115.760 -136.015 ;
        RECT -114.620 -245.175 -114.240 -140.585 ;
        RECT -113.100 -240.605 -112.720 -136.015 ;
        RECT -111.580 -245.175 -111.200 -140.585 ;
        RECT -110.060 -240.605 -109.680 -136.015 ;
        RECT -108.540 -245.175 -108.160 -140.585 ;
        RECT -107.020 -240.605 -106.640 -136.015 ;
        RECT -105.500 -245.175 -105.120 -140.585 ;
        RECT -103.980 -240.605 -103.600 -136.015 ;
        RECT -102.460 -245.175 -102.080 -140.585 ;
        RECT -100.940 -240.605 -100.560 -136.015 ;
        RECT -99.420 -245.175 -99.040 -140.585 ;
        RECT -97.900 -240.605 -97.520 -136.015 ;
        RECT -96.380 -245.175 -96.000 -140.585 ;
        RECT -94.860 -240.605 -94.480 -136.015 ;
        RECT -93.340 -245.175 -92.960 -140.585 ;
        RECT -91.820 -240.605 -91.440 -136.015 ;
        RECT -90.300 -245.175 -89.920 -140.585 ;
        RECT -88.780 -240.605 -88.400 -136.015 ;
        RECT -87.260 -245.175 -86.880 -140.585 ;
        RECT -85.740 -240.605 -85.360 -136.015 ;
        RECT -84.220 -245.175 -83.840 -140.585 ;
        RECT -82.700 -240.605 -82.320 -136.015 ;
        RECT -81.180 -245.175 -80.800 -140.585 ;
        RECT -79.660 -240.605 -79.280 -136.015 ;
        RECT -78.140 -245.175 -77.760 -140.585 ;
        RECT -76.620 -240.605 -76.240 -136.015 ;
        RECT -75.100 -245.175 -74.720 -140.585 ;
        RECT -73.580 -240.605 -73.200 -136.015 ;
        RECT -65.580 -140.595 -65.200 -136.015 ;
        RECT -66.370 -240.605 -65.200 -140.595 ;
        RECT -64.060 -245.175 -63.680 -140.585 ;
        RECT -62.540 -240.605 -62.160 -136.015 ;
        RECT -61.020 -245.175 -60.640 -140.585 ;
        RECT -59.500 -240.605 -59.120 -136.015 ;
        RECT -57.980 -245.175 -57.600 -140.585 ;
        RECT -56.460 -240.605 -56.080 -136.015 ;
        RECT -54.940 -245.175 -54.560 -140.585 ;
        RECT -53.420 -240.605 -53.040 -136.015 ;
        RECT -51.900 -245.175 -51.520 -140.585 ;
        RECT -50.380 -240.605 -50.000 -136.015 ;
        RECT -48.860 -245.175 -48.480 -140.585 ;
        RECT -47.340 -240.605 -46.960 -136.015 ;
        RECT -45.820 -245.175 -45.440 -140.585 ;
        RECT -44.300 -240.605 -43.920 -136.015 ;
        RECT -42.780 -245.175 -42.400 -140.585 ;
        RECT -41.260 -240.605 -40.880 -136.015 ;
        RECT -39.740 -245.175 -39.360 -140.585 ;
        RECT -38.220 -240.605 -37.840 -136.015 ;
        RECT -36.700 -245.175 -36.320 -140.585 ;
        RECT -35.180 -240.605 -34.800 -136.015 ;
        RECT -33.660 -245.175 -33.280 -140.585 ;
        RECT -32.140 -240.605 -31.760 -136.015 ;
        RECT -30.620 -245.175 -30.240 -140.585 ;
        RECT -29.100 -240.605 -28.720 -136.015 ;
        RECT -27.580 -245.175 -27.200 -140.585 ;
        RECT -26.060 -240.605 -25.680 -136.015 ;
        RECT -24.540 -245.175 -24.160 -140.585 ;
        RECT -23.020 -240.605 -22.640 -136.015 ;
        RECT -21.500 -245.175 -21.120 -140.585 ;
        RECT -19.980 -240.605 -19.600 -136.015 ;
        RECT -18.460 -245.175 -18.080 -140.585 ;
        RECT -16.940 -240.605 -16.560 -136.015 ;
        RECT -15.420 -245.175 -15.040 -140.585 ;
        RECT -13.900 -240.605 -13.520 -136.015 ;
        RECT -12.380 -245.175 -12.000 -140.585 ;
        RECT -10.860 -240.605 -10.480 -136.015 ;
        RECT -9.340 -245.175 -8.960 -140.585 ;
        RECT -7.820 -240.605 -7.440 -136.015 ;
        RECT -6.300 -245.175 -5.920 -140.585 ;
        RECT -4.780 -240.605 -4.400 -136.015 ;
        RECT -3.260 -245.175 -2.880 -140.585 ;
        RECT -1.740 -240.605 -1.360 -136.015 ;
        RECT -0.220 -245.175 0.160 -140.585 ;
        RECT 1.300 -240.605 1.680 -136.015 ;
        RECT 2.820 -245.175 3.200 -140.585 ;
        RECT 4.340 -240.605 4.720 -136.015 ;
        RECT 5.860 -245.175 6.240 -140.585 ;
        RECT 7.380 -240.605 7.760 -136.015 ;
        RECT 8.900 -245.175 9.280 -140.585 ;
        RECT 10.420 -240.605 10.800 -136.015 ;
        RECT 11.940 -245.175 12.320 -140.585 ;
        RECT 13.460 -240.605 13.840 -136.015 ;
        RECT 14.980 -245.175 15.360 -140.585 ;
        RECT 16.500 -240.605 16.880 -136.015 ;
        RECT 18.020 -245.175 18.400 -140.585 ;
        RECT 19.540 -240.605 19.920 -136.015 ;
        RECT 21.060 -245.175 21.440 -140.585 ;
        RECT 22.580 -240.605 22.960 -136.015 ;
        RECT 24.100 -245.175 24.480 -140.585 ;
        RECT 25.620 -240.605 26.000 -136.015 ;
        RECT 27.140 -245.175 27.520 -140.585 ;
        RECT 28.660 -240.605 29.040 -136.015 ;
        RECT 30.180 -245.175 30.560 -140.585 ;
        RECT 31.700 -240.605 32.080 -136.015 ;
        RECT 33.220 -245.175 33.600 -140.585 ;
        RECT 34.740 -240.605 35.120 -136.015 ;
        RECT 36.260 -245.175 36.640 -140.585 ;
        RECT 37.780 -240.605 38.160 -136.015 ;
        RECT 39.300 -245.175 39.680 -140.585 ;
        RECT 40.820 -240.605 41.200 -136.015 ;
        RECT 42.340 -245.175 42.720 -140.585 ;
        RECT 43.860 -240.605 44.240 -136.015 ;
        RECT 45.380 -245.175 45.760 -140.585 ;
        RECT 46.900 -240.605 47.280 -136.015 ;
        RECT 48.420 -245.175 48.800 -140.585 ;
        RECT 49.940 -240.605 50.320 -136.015 ;
        RECT 51.460 -245.175 51.840 -140.585 ;
        RECT 52.980 -240.605 53.360 -136.015 ;
        RECT 54.500 -245.175 54.880 -140.585 ;
        RECT 56.020 -240.605 56.400 -136.015 ;
        RECT 57.540 -245.175 57.920 -140.585 ;
        RECT 59.060 -240.605 59.440 -136.015 ;
        RECT 60.580 -245.175 60.960 -140.585 ;
        RECT 62.100 -240.605 62.480 -136.015 ;
        RECT 63.620 -245.175 64.000 -140.585 ;
        RECT 65.140 -240.605 65.520 -136.015 ;
        RECT 66.660 -245.175 67.040 -140.585 ;
        RECT 68.180 -240.605 68.560 -136.015 ;
        RECT 69.700 -245.175 70.080 -140.585 ;
        RECT 71.220 -240.605 71.600 -136.015 ;
        RECT 72.740 -245.175 73.120 -140.585 ;
        RECT 74.260 -240.605 74.640 -136.015 ;
        RECT 75.780 -245.175 76.160 -140.585 ;
        RECT 77.300 -240.605 77.680 -136.015 ;
        RECT 78.820 -245.175 79.200 -140.585 ;
        RECT 80.340 -240.605 80.720 -136.015 ;
        RECT 81.860 -245.175 82.240 -140.585 ;
        RECT 83.380 -240.605 83.760 -136.015 ;
        RECT 84.900 -245.175 85.280 -140.585 ;
        RECT 86.420 -240.605 86.800 -136.015 ;
        RECT 94.420 -140.595 94.800 -136.015 ;
        RECT 93.630 -240.605 94.800 -140.595 ;
        RECT 95.940 -245.175 96.320 -140.585 ;
        RECT 97.460 -240.605 97.840 -136.015 ;
        RECT 98.980 -245.175 99.360 -140.585 ;
        RECT 100.500 -240.605 100.880 -136.015 ;
        RECT 102.020 -245.175 102.400 -140.585 ;
        RECT 103.540 -240.605 103.920 -136.015 ;
        RECT 105.060 -245.175 105.440 -140.585 ;
        RECT 106.580 -240.605 106.960 -136.015 ;
        RECT 108.100 -245.175 108.480 -140.585 ;
        RECT 109.620 -240.605 110.000 -136.015 ;
        RECT 111.140 -245.175 111.520 -140.585 ;
        RECT 112.660 -240.605 113.040 -136.015 ;
        RECT 114.180 -245.175 114.560 -140.585 ;
        RECT 115.700 -240.605 116.080 -136.015 ;
        RECT 117.220 -245.175 117.600 -140.585 ;
        RECT 118.740 -240.605 119.120 -136.015 ;
        RECT 120.260 -245.175 120.640 -140.585 ;
        RECT 121.780 -240.605 122.160 -136.015 ;
        RECT 123.300 -245.175 123.680 -140.585 ;
        RECT 124.820 -240.605 125.200 -136.015 ;
        RECT 126.340 -245.175 126.720 -140.585 ;
        RECT 127.860 -240.605 128.240 -136.015 ;
        RECT 129.380 -245.175 129.760 -140.585 ;
        RECT 130.900 -240.605 131.280 -136.015 ;
        RECT 132.420 -245.175 132.800 -140.585 ;
        RECT 133.940 -240.605 134.320 -136.015 ;
        RECT 135.460 -245.175 135.840 -140.585 ;
        RECT 136.980 -240.605 137.360 -136.015 ;
        RECT 138.500 -245.175 138.880 -140.585 ;
        RECT 140.020 -240.605 140.400 -136.015 ;
        RECT 141.540 -245.175 141.920 -140.585 ;
        RECT 143.060 -240.605 143.440 -136.015 ;
        RECT 144.580 -245.175 144.960 -140.585 ;
        RECT 146.100 -240.605 146.480 -136.015 ;
        RECT 147.620 -245.175 148.000 -140.585 ;
        RECT 149.140 -240.605 149.520 -136.015 ;
        RECT 150.660 -245.175 151.040 -140.585 ;
        RECT 152.180 -240.605 152.560 -136.015 ;
        RECT 153.700 -245.175 154.080 -140.585 ;
        RECT 155.220 -240.605 155.600 -136.015 ;
        RECT 156.740 -245.175 157.120 -140.585 ;
        RECT 158.260 -240.605 158.640 -136.015 ;
        RECT 159.780 -245.175 160.160 -140.585 ;
        RECT 161.300 -240.605 161.680 -136.015 ;
        RECT 162.820 -245.175 163.200 -140.585 ;
        RECT 164.340 -240.605 164.720 -136.015 ;
        RECT 165.860 -245.175 166.240 -140.585 ;
        RECT 167.380 -240.605 167.760 -136.015 ;
        RECT 168.900 -245.175 169.280 -140.585 ;
        RECT 170.420 -240.605 170.800 -136.015 ;
        RECT 171.940 -245.175 172.320 -140.585 ;
        RECT 173.460 -240.605 173.840 -136.015 ;
        RECT 174.980 -245.175 175.360 -140.585 ;
        RECT 176.500 -240.605 176.880 -136.015 ;
        RECT 178.020 -245.175 178.400 -140.585 ;
        RECT 179.540 -240.605 179.920 -136.015 ;
        RECT 181.060 -245.175 181.440 -140.585 ;
        RECT 182.580 -240.605 182.960 -136.015 ;
        RECT 184.100 -245.175 184.480 -140.585 ;
        RECT 185.620 -240.605 186.000 -136.015 ;
        RECT 187.140 -245.175 187.520 -140.585 ;
        RECT 188.660 -240.605 189.040 -136.015 ;
        RECT 190.180 -245.175 190.560 -140.585 ;
        RECT 191.700 -240.605 192.080 -136.015 ;
        RECT 193.220 -245.175 193.600 -140.585 ;
        RECT 194.740 -240.605 195.120 -136.015 ;
        RECT 196.260 -245.175 196.640 -140.585 ;
        RECT 197.780 -240.605 198.160 -136.015 ;
        RECT 199.300 -245.175 199.680 -140.585 ;
        RECT 200.820 -240.605 201.200 -136.015 ;
        RECT 202.340 -245.175 202.720 -140.585 ;
        RECT 203.860 -240.605 204.240 -136.015 ;
        RECT 205.380 -245.175 205.760 -140.585 ;
        RECT 206.900 -240.605 207.280 -136.015 ;
        RECT 208.420 -245.175 208.800 -140.585 ;
        RECT 209.940 -240.605 210.320 -136.015 ;
        RECT 211.460 -245.175 211.840 -140.585 ;
        RECT 212.980 -240.605 213.360 -136.015 ;
        RECT 214.500 -245.175 214.880 -140.585 ;
        RECT 216.020 -240.605 216.400 -136.015 ;
        RECT 217.540 -245.175 217.920 -140.585 ;
        RECT 219.060 -240.605 219.440 -136.015 ;
        RECT 220.580 -245.175 220.960 -140.585 ;
        RECT 222.100 -240.605 222.480 -136.015 ;
        RECT 223.620 -245.175 224.000 -140.585 ;
        RECT 225.140 -240.605 225.520 -136.015 ;
        RECT 226.660 -245.175 227.040 -140.585 ;
        RECT 228.180 -240.605 228.560 -136.015 ;
        RECT 229.700 -245.175 230.080 -140.585 ;
        RECT 231.220 -240.605 231.600 -136.015 ;
        RECT 232.740 -245.175 233.120 -140.585 ;
        RECT 234.260 -240.605 234.640 -136.015 ;
        RECT 235.780 -245.175 236.160 -140.585 ;
        RECT 237.300 -240.605 237.680 -136.015 ;
        RECT 238.820 -245.175 239.200 -140.585 ;
        RECT 240.340 -240.605 240.720 -136.015 ;
        RECT 241.860 -245.175 242.240 -140.585 ;
        RECT 243.380 -240.605 243.760 -136.015 ;
        RECT 244.900 -245.175 245.280 -140.585 ;
        RECT 246.420 -240.605 246.800 -136.015 ;
        RECT 254.420 -140.595 254.800 -136.015 ;
        RECT 253.630 -240.605 254.800 -140.595 ;
        RECT 255.940 -245.175 256.320 -140.585 ;
        RECT 257.460 -240.605 257.840 -136.015 ;
        RECT 258.980 -245.175 259.360 -140.585 ;
        RECT 260.500 -240.605 260.880 -136.015 ;
        RECT 262.020 -245.175 262.400 -140.585 ;
        RECT 263.540 -240.605 263.920 -136.015 ;
        RECT 265.060 -245.175 265.440 -140.585 ;
        RECT 266.580 -240.605 266.960 -136.015 ;
        RECT 268.100 -245.175 268.480 -140.585 ;
        RECT 269.620 -240.605 270.000 -136.015 ;
        RECT 271.140 -245.175 271.520 -140.585 ;
        RECT 272.660 -240.605 273.040 -136.015 ;
        RECT 274.180 -245.175 274.560 -140.585 ;
        RECT 275.700 -240.605 276.080 -136.015 ;
        RECT 277.220 -245.175 277.600 -140.585 ;
        RECT 278.740 -240.605 279.120 -136.015 ;
        RECT 280.260 -245.175 280.640 -140.585 ;
        RECT 281.780 -240.605 282.160 -136.015 ;
        RECT 283.300 -245.175 283.680 -140.585 ;
        RECT 284.820 -240.605 285.200 -136.015 ;
        RECT 286.340 -245.175 286.720 -140.585 ;
        RECT 287.860 -240.605 288.240 -136.015 ;
        RECT 289.380 -245.175 289.760 -140.585 ;
        RECT 290.900 -240.605 291.280 -136.015 ;
        RECT 292.420 -245.175 292.800 -140.585 ;
        RECT 293.940 -240.605 294.320 -136.015 ;
        RECT 295.460 -245.175 295.840 -140.585 ;
        RECT 296.980 -240.605 297.360 -136.015 ;
        RECT 298.500 -245.175 298.880 -140.585 ;
        RECT 300.020 -240.605 300.400 -136.015 ;
        RECT 301.540 -245.175 301.920 -140.585 ;
        RECT 303.060 -240.605 303.440 -136.015 ;
        RECT 304.580 -245.175 304.960 -140.585 ;
        RECT 306.100 -240.605 306.480 -136.015 ;
        RECT 307.620 -245.175 308.000 -140.585 ;
        RECT 309.140 -240.605 309.520 -136.015 ;
        RECT 310.660 -245.175 311.040 -140.585 ;
        RECT 312.180 -240.605 312.560 -136.015 ;
        RECT 313.700 -245.175 314.080 -140.585 ;
        RECT 315.220 -240.605 315.600 -136.015 ;
        RECT 316.740 -245.175 317.120 -140.585 ;
        RECT 318.260 -240.605 318.640 -136.015 ;
        RECT 319.780 -245.175 320.160 -140.585 ;
        RECT 321.300 -240.605 321.680 -136.015 ;
        RECT 322.820 -245.175 323.200 -140.585 ;
        RECT 324.340 -240.605 324.720 -136.015 ;
        RECT 325.860 -245.175 326.240 -140.585 ;
        RECT 327.380 -240.605 327.760 -136.015 ;
        RECT 328.900 -245.175 329.280 -140.585 ;
        RECT 330.420 -240.605 330.800 -136.015 ;
        RECT 331.940 -245.175 332.320 -140.585 ;
        RECT 333.460 -240.605 333.840 -136.015 ;
        RECT 334.980 -245.175 335.360 -140.585 ;
        RECT 336.500 -240.605 336.880 -136.015 ;
        RECT 338.020 -245.175 338.400 -140.585 ;
        RECT 339.540 -240.605 339.920 -136.015 ;
        RECT 341.060 -245.175 341.440 -140.585 ;
        RECT 342.580 -240.605 342.960 -136.015 ;
        RECT 344.100 -245.175 344.480 -140.585 ;
        RECT 345.620 -240.605 346.000 -136.015 ;
        RECT 347.140 -245.175 347.520 -140.585 ;
        RECT 348.660 -240.605 349.040 -136.015 ;
        RECT 350.180 -245.175 350.560 -140.585 ;
        RECT 351.700 -240.605 352.080 -136.015 ;
        RECT 353.220 -245.175 353.600 -140.585 ;
        RECT 354.740 -240.605 355.120 -136.015 ;
        RECT 356.260 -245.175 356.640 -140.585 ;
        RECT 357.780 -240.605 358.160 -136.015 ;
        RECT 359.300 -245.175 359.680 -140.585 ;
        RECT 360.820 -240.605 361.200 -136.015 ;
        RECT 362.340 -245.175 362.720 -140.585 ;
        RECT 363.860 -240.605 364.240 -136.015 ;
        RECT 365.380 -245.175 365.760 -140.585 ;
        RECT 366.900 -240.605 367.280 -136.015 ;
        RECT 368.420 -245.175 368.800 -140.585 ;
        RECT 369.940 -240.605 370.320 -136.015 ;
        RECT 371.460 -245.175 371.840 -140.585 ;
        RECT 372.980 -240.605 373.360 -136.015 ;
        RECT 374.500 -245.175 374.880 -140.585 ;
        RECT 376.020 -240.605 376.400 -136.015 ;
        RECT 377.540 -245.175 377.920 -140.585 ;
        RECT 379.060 -240.605 379.440 -136.015 ;
        RECT 380.580 -245.175 380.960 -140.585 ;
        RECT 382.100 -240.605 382.480 -136.015 ;
        RECT 383.620 -245.175 384.000 -140.585 ;
        RECT 385.140 -240.605 385.520 -136.015 ;
        RECT 386.660 -245.175 387.040 -140.585 ;
        RECT 388.180 -240.605 388.560 -136.015 ;
        RECT 389.700 -245.175 390.080 -140.585 ;
        RECT 391.220 -240.605 391.600 -136.015 ;
        RECT 392.740 -245.175 393.120 -140.585 ;
        RECT 394.260 -240.605 394.640 -136.015 ;
        RECT 395.780 -245.175 396.160 -140.585 ;
        RECT 397.300 -240.605 397.680 -136.015 ;
        RECT 398.820 -245.175 399.200 -140.585 ;
        RECT 400.340 -240.605 400.720 -136.015 ;
        RECT 401.860 -245.175 402.240 -140.585 ;
        RECT 403.380 -240.605 403.760 -136.015 ;
        RECT 404.900 -245.175 405.280 -140.585 ;
        RECT 406.420 -240.605 406.800 -136.015 ;
        RECT 414.420 -140.595 414.800 -136.015 ;
        RECT 413.630 -240.605 414.800 -140.595 ;
        RECT 415.940 -245.175 416.320 -140.585 ;
        RECT 417.460 -240.605 417.840 -136.015 ;
        RECT 418.980 -245.175 419.360 -140.585 ;
        RECT 420.500 -240.605 420.880 -136.015 ;
        RECT 422.020 -245.175 422.400 -140.585 ;
        RECT 423.540 -240.605 423.920 -136.015 ;
        RECT 425.060 -245.175 425.440 -140.585 ;
        RECT 426.580 -240.605 426.960 -136.015 ;
        RECT 428.100 -245.175 428.480 -140.585 ;
        RECT 429.620 -240.605 430.000 -136.015 ;
        RECT 431.140 -245.175 431.520 -140.585 ;
        RECT 432.660 -240.605 433.040 -136.015 ;
        RECT 434.180 -245.175 434.560 -140.585 ;
        RECT 435.700 -240.605 436.080 -136.015 ;
        RECT 437.220 -245.175 437.600 -140.585 ;
        RECT 438.740 -240.605 439.120 -136.015 ;
        RECT 440.260 -245.175 440.640 -140.585 ;
        RECT 441.780 -240.605 442.160 -136.015 ;
        RECT 443.300 -245.175 443.680 -140.585 ;
        RECT 444.820 -240.605 445.200 -136.015 ;
        RECT 446.340 -245.175 446.720 -140.585 ;
        RECT 447.860 -240.605 448.240 -136.015 ;
        RECT 449.380 -245.175 449.760 -140.585 ;
        RECT 450.900 -240.605 451.280 -136.015 ;
        RECT 452.420 -245.175 452.800 -140.585 ;
        RECT 453.940 -240.605 454.320 -136.015 ;
        RECT 455.460 -245.175 455.840 -140.585 ;
        RECT 456.980 -240.605 457.360 -136.015 ;
        RECT 458.500 -245.175 458.880 -140.585 ;
        RECT 460.020 -240.605 460.400 -136.015 ;
        RECT 461.540 -245.175 461.920 -140.585 ;
        RECT 463.060 -240.605 463.440 -136.015 ;
        RECT 464.580 -245.175 464.960 -140.585 ;
        RECT 466.100 -240.605 466.480 -136.015 ;
        RECT 467.620 -245.175 468.000 -140.585 ;
        RECT 469.140 -240.605 469.520 -136.015 ;
        RECT 470.660 -245.175 471.040 -140.585 ;
        RECT 472.180 -240.605 472.560 -136.015 ;
        RECT 473.700 -245.175 474.080 -140.585 ;
        RECT 475.220 -240.605 475.600 -136.015 ;
        RECT 476.740 -245.175 477.120 -140.585 ;
        RECT 478.260 -240.605 478.640 -136.015 ;
        RECT 479.780 -245.175 480.160 -140.585 ;
        RECT 481.300 -240.605 481.680 -136.015 ;
        RECT 482.820 -245.175 483.200 -140.585 ;
        RECT 484.340 -240.605 484.720 -136.015 ;
        RECT 485.860 -245.175 486.240 -140.585 ;
        RECT 487.380 -240.605 487.760 -136.015 ;
        RECT 488.900 -245.175 489.280 -140.585 ;
        RECT 490.420 -240.605 490.800 -136.015 ;
        RECT 491.940 -245.175 492.320 -140.585 ;
        RECT 493.460 -240.605 493.840 -136.015 ;
        RECT 494.980 -245.175 495.360 -140.585 ;
        RECT 496.500 -240.605 496.880 -136.015 ;
        RECT 498.020 -245.175 498.400 -140.585 ;
        RECT 499.540 -240.605 499.920 -136.015 ;
        RECT 501.060 -245.175 501.440 -140.585 ;
        RECT 502.580 -240.605 502.960 -136.015 ;
        RECT 504.100 -245.175 504.480 -140.585 ;
        RECT 505.620 -240.605 506.000 -136.015 ;
        RECT 507.140 -245.175 507.520 -140.585 ;
        RECT 508.660 -240.605 509.040 -136.015 ;
        RECT 510.180 -245.175 510.560 -140.585 ;
        RECT 511.700 -240.605 512.080 -136.015 ;
        RECT 513.220 -245.175 513.600 -140.585 ;
        RECT 514.740 -240.605 515.120 -136.015 ;
        RECT 516.260 -245.175 516.640 -140.585 ;
        RECT 517.780 -240.605 518.160 -136.015 ;
        RECT 519.300 -245.175 519.680 -140.585 ;
        RECT 520.820 -240.605 521.200 -136.015 ;
        RECT 522.340 -245.175 522.720 -140.585 ;
        RECT 523.860 -240.605 524.240 -136.015 ;
        RECT 525.380 -245.175 525.760 -140.585 ;
        RECT 526.900 -240.605 527.280 -136.015 ;
        RECT 528.420 -245.175 528.800 -140.585 ;
        RECT 529.940 -240.605 530.320 -136.015 ;
        RECT 531.460 -245.175 531.840 -140.585 ;
        RECT 532.980 -240.605 533.360 -136.015 ;
        RECT 534.500 -245.175 534.880 -140.585 ;
        RECT 536.020 -240.605 536.400 -136.015 ;
        RECT 537.540 -245.175 537.920 -140.585 ;
        RECT 539.060 -240.605 539.440 -136.015 ;
        RECT 540.580 -245.175 540.960 -140.585 ;
        RECT 542.100 -240.605 542.480 -136.015 ;
        RECT 543.620 -245.175 544.000 -140.585 ;
        RECT 545.140 -240.605 545.520 -136.015 ;
        RECT 546.660 -245.175 547.040 -140.585 ;
        RECT 548.180 -240.605 548.560 -136.015 ;
        RECT 549.700 -245.175 550.080 -140.585 ;
        RECT 551.220 -240.605 551.600 -136.015 ;
        RECT 552.740 -245.175 553.120 -140.585 ;
        RECT 554.260 -240.605 554.640 -136.015 ;
        RECT 555.780 -245.175 556.160 -140.585 ;
        RECT 557.300 -240.605 557.680 -136.015 ;
        RECT 558.820 -245.175 559.200 -140.585 ;
        RECT 560.340 -240.605 560.720 -136.015 ;
        RECT 561.860 -245.175 562.240 -140.585 ;
        RECT 563.380 -240.605 563.760 -136.015 ;
        RECT 564.900 -245.175 565.280 -140.585 ;
        RECT 566.420 -240.605 566.800 -136.015 ;
        RECT 574.420 -140.595 574.800 -136.015 ;
        RECT 573.630 -240.605 574.800 -140.595 ;
        RECT 575.940 -245.175 576.320 -140.585 ;
        RECT 577.460 -240.605 577.840 -136.015 ;
        RECT 578.980 -245.175 579.360 -140.585 ;
        RECT 580.500 -240.605 580.880 -136.015 ;
        RECT 582.020 -245.175 582.400 -140.585 ;
        RECT 583.540 -240.605 583.920 -136.015 ;
        RECT 585.060 -245.175 585.440 -140.585 ;
        RECT 586.580 -240.605 586.960 -136.015 ;
        RECT 588.100 -245.175 588.480 -140.585 ;
        RECT 589.620 -240.605 590.000 -136.015 ;
        RECT 591.140 -245.175 591.520 -140.585 ;
        RECT 592.660 -240.605 593.040 -136.015 ;
        RECT 594.180 -245.175 594.560 -140.585 ;
        RECT 595.700 -240.605 596.080 -136.015 ;
        RECT 597.220 -245.175 597.600 -140.585 ;
        RECT 598.740 -240.605 599.120 -136.015 ;
        RECT 600.260 -245.175 600.640 -140.585 ;
        RECT 601.780 -240.605 602.160 -136.015 ;
        RECT 603.300 -245.175 603.680 -140.585 ;
        RECT 604.820 -240.605 605.200 -136.015 ;
        RECT 606.340 -245.175 606.720 -140.585 ;
        RECT 607.860 -240.605 608.240 -136.015 ;
        RECT 609.380 -245.175 609.760 -140.585 ;
        RECT 610.900 -240.605 611.280 -136.015 ;
        RECT 612.420 -245.175 612.800 -140.585 ;
        RECT 613.940 -240.605 614.320 -136.015 ;
        RECT 615.460 -245.175 615.840 -140.585 ;
        RECT 616.980 -240.605 617.360 -136.015 ;
        RECT 618.500 -245.175 618.880 -140.585 ;
        RECT 620.020 -240.605 620.400 -136.015 ;
        RECT 621.540 -245.175 621.920 -140.585 ;
        RECT 623.060 -240.605 623.440 -136.015 ;
        RECT 624.580 -245.175 624.960 -140.585 ;
        RECT 626.100 -240.605 626.480 -136.015 ;
        RECT 627.620 -245.175 628.000 -140.585 ;
        RECT 629.140 -240.605 629.520 -136.015 ;
        RECT 630.660 -245.175 631.040 -140.585 ;
        RECT 632.180 -240.605 632.560 -136.015 ;
        RECT 633.700 -245.175 634.080 -140.585 ;
        RECT 635.220 -240.605 635.600 -136.015 ;
        RECT 636.740 -245.175 637.120 -140.585 ;
        RECT 638.260 -240.605 638.640 -136.015 ;
        RECT 639.780 -245.175 640.160 -140.585 ;
        RECT 641.300 -240.605 641.680 -136.015 ;
        RECT 642.820 -245.175 643.200 -140.585 ;
        RECT 644.340 -240.605 644.720 -136.015 ;
        RECT 645.860 -245.175 646.240 -140.585 ;
        RECT 647.380 -240.605 647.760 -136.015 ;
        RECT 648.900 -245.175 649.280 -140.585 ;
        RECT 650.420 -240.605 650.800 -136.015 ;
        RECT 651.940 -245.175 652.320 -140.585 ;
        RECT 653.460 -240.605 653.840 -136.015 ;
        RECT 654.980 -245.175 655.360 -140.585 ;
        RECT 656.500 -240.605 656.880 -136.015 ;
        RECT 658.020 -245.175 658.400 -140.585 ;
        RECT 659.540 -240.605 659.920 -136.015 ;
        RECT 661.060 -245.175 661.440 -140.585 ;
        RECT 662.580 -240.605 662.960 -136.015 ;
        RECT 664.100 -245.175 664.480 -140.585 ;
        RECT 665.620 -240.605 666.000 -136.015 ;
        RECT 667.140 -245.175 667.520 -140.585 ;
        RECT 668.660 -240.605 669.040 -136.015 ;
        RECT 670.180 -245.175 670.560 -140.585 ;
        RECT 671.700 -240.605 672.080 -136.015 ;
        RECT 673.220 -245.175 673.600 -140.585 ;
        RECT 674.740 -240.605 675.120 -136.015 ;
        RECT 676.260 -245.175 676.640 -140.585 ;
        RECT 677.780 -240.605 678.160 -136.015 ;
        RECT 679.300 -245.175 679.680 -140.585 ;
        RECT 680.820 -240.605 681.200 -136.015 ;
        RECT 682.340 -245.175 682.720 -140.585 ;
        RECT 683.860 -240.605 684.240 -136.015 ;
        RECT 685.380 -245.175 685.760 -140.585 ;
        RECT 686.900 -240.605 687.280 -136.015 ;
        RECT 688.420 -245.175 688.800 -140.585 ;
        RECT 689.940 -240.605 690.320 -136.015 ;
        RECT 691.460 -245.175 691.840 -140.585 ;
        RECT 692.980 -240.605 693.360 -136.015 ;
        RECT 694.500 -245.175 694.880 -140.585 ;
        RECT 696.020 -240.605 696.400 -136.015 ;
        RECT 697.540 -245.175 697.920 -140.585 ;
        RECT 699.060 -240.605 699.440 -136.015 ;
        RECT 700.580 -245.175 700.960 -140.585 ;
        RECT 702.100 -240.605 702.480 -136.015 ;
        RECT 703.620 -245.175 704.000 -140.585 ;
        RECT 705.140 -240.605 705.520 -136.015 ;
        RECT 706.660 -245.175 707.040 -140.585 ;
        RECT 708.180 -240.605 708.560 -136.015 ;
        RECT 709.700 -245.175 710.080 -140.585 ;
        RECT 711.220 -240.605 711.600 -136.015 ;
        RECT 712.740 -245.175 713.120 -140.585 ;
        RECT 714.260 -240.605 714.640 -136.015 ;
        RECT 715.780 -245.175 716.160 -140.585 ;
        RECT 717.300 -240.605 717.680 -136.015 ;
        RECT 718.820 -245.175 719.200 -140.585 ;
        RECT 720.340 -240.605 720.720 -136.015 ;
        RECT 721.860 -245.175 722.240 -140.585 ;
        RECT 723.380 -240.605 723.760 -136.015 ;
        RECT 724.900 -245.175 725.280 -140.585 ;
        RECT 726.420 -240.605 726.800 -136.015 ;
        RECT 734.420 -140.595 734.800 -136.015 ;
        RECT 733.630 -240.605 734.800 -140.595 ;
        RECT 735.940 -245.175 736.320 -140.585 ;
        RECT 737.460 -240.605 737.840 -136.015 ;
        RECT 738.980 -245.175 739.360 -140.585 ;
        RECT 740.500 -240.605 740.880 -136.015 ;
        RECT 742.020 -245.175 742.400 -140.585 ;
        RECT 743.540 -240.605 743.920 -136.015 ;
        RECT 745.060 -245.175 745.440 -140.585 ;
        RECT 746.580 -240.605 746.960 -136.015 ;
        RECT 748.100 -245.175 748.480 -140.585 ;
        RECT 749.620 -240.605 750.000 -136.015 ;
        RECT 751.140 -245.175 751.520 -140.585 ;
        RECT 752.660 -240.605 753.040 -136.015 ;
        RECT 754.180 -245.175 754.560 -140.585 ;
        RECT 755.700 -240.605 756.080 -136.015 ;
        RECT 757.220 -245.175 757.600 -140.585 ;
        RECT 758.740 -240.605 759.120 -136.015 ;
        RECT 760.260 -245.175 760.640 -140.585 ;
        RECT 761.780 -240.605 762.160 -136.015 ;
        RECT 763.300 -245.175 763.680 -140.585 ;
        RECT 764.820 -240.605 765.200 -136.015 ;
        RECT 766.340 -245.175 766.720 -140.585 ;
        RECT 767.860 -240.605 768.240 -136.015 ;
        RECT 769.380 -245.175 769.760 -140.585 ;
        RECT 770.900 -240.605 771.280 -136.015 ;
        RECT 772.420 -245.175 772.800 -140.585 ;
        RECT 773.940 -240.605 774.320 -136.015 ;
        RECT 775.460 -245.175 775.840 -140.585 ;
        RECT 776.980 -240.605 777.360 -136.015 ;
        RECT 778.500 -245.175 778.880 -140.585 ;
        RECT 780.020 -240.605 780.400 -136.015 ;
        RECT 781.540 -245.175 781.920 -140.585 ;
        RECT 783.060 -240.605 783.440 -136.015 ;
        RECT 784.580 -245.175 784.960 -140.585 ;
        RECT 786.100 -240.605 786.480 -136.015 ;
        RECT 787.620 -245.175 788.000 -140.585 ;
        RECT 789.140 -240.605 789.520 -136.015 ;
        RECT 790.660 -245.175 791.040 -140.585 ;
        RECT 792.180 -240.605 792.560 -136.015 ;
        RECT 793.700 -245.175 794.080 -140.585 ;
        RECT 795.220 -240.605 795.600 -136.015 ;
        RECT 796.740 -245.175 797.120 -140.585 ;
        RECT 798.260 -240.605 798.640 -136.015 ;
        RECT 799.780 -245.175 800.160 -140.585 ;
        RECT 801.300 -240.605 801.680 -136.015 ;
        RECT 802.820 -245.175 803.200 -140.585 ;
        RECT 804.340 -240.605 804.720 -136.015 ;
        RECT 805.860 -245.175 806.240 -140.585 ;
        RECT 807.380 -240.605 807.760 -136.015 ;
        RECT 808.900 -245.175 809.280 -140.585 ;
        RECT 810.420 -240.605 810.800 -136.015 ;
        RECT 811.940 -245.175 812.320 -140.585 ;
        RECT 813.460 -240.605 813.840 -136.015 ;
        RECT 814.980 -245.175 815.360 -140.585 ;
        RECT 816.500 -240.605 816.880 -136.015 ;
        RECT 818.020 -245.175 818.400 -140.585 ;
        RECT 819.540 -240.605 819.920 -136.015 ;
        RECT 821.060 -245.175 821.440 -140.585 ;
        RECT 822.580 -240.605 822.960 -136.015 ;
        RECT 824.100 -245.175 824.480 -140.585 ;
        RECT 825.620 -240.605 826.000 -136.015 ;
        RECT 827.140 -245.175 827.520 -140.585 ;
        RECT 828.660 -240.605 829.040 -136.015 ;
        RECT 830.180 -245.175 830.560 -140.585 ;
        RECT 831.700 -240.605 832.080 -136.015 ;
        RECT 833.220 -245.175 833.600 -140.585 ;
        RECT 834.740 -240.605 835.120 -136.015 ;
        RECT 836.260 -245.175 836.640 -140.585 ;
        RECT 837.780 -240.605 838.160 -136.015 ;
        RECT 839.300 -245.175 839.680 -140.585 ;
        RECT 840.820 -240.605 841.200 -136.015 ;
        RECT 842.340 -245.175 842.720 -140.585 ;
        RECT 843.860 -240.605 844.240 -136.015 ;
        RECT 845.380 -245.175 845.760 -140.585 ;
        RECT 846.900 -240.605 847.280 -136.015 ;
        RECT 848.420 -245.175 848.800 -140.585 ;
        RECT 849.940 -240.605 850.320 -136.015 ;
        RECT 851.460 -245.175 851.840 -140.585 ;
        RECT 852.980 -240.605 853.360 -136.015 ;
        RECT 854.500 -245.175 854.880 -140.585 ;
        RECT 856.020 -240.605 856.400 -136.015 ;
        RECT 857.540 -245.175 857.920 -140.585 ;
        RECT 859.060 -240.605 859.440 -136.015 ;
        RECT 860.580 -245.175 860.960 -140.585 ;
        RECT 862.100 -240.605 862.480 -136.015 ;
        RECT 863.620 -245.175 864.000 -140.585 ;
        RECT 865.140 -240.605 865.520 -136.015 ;
        RECT 866.660 -245.175 867.040 -140.585 ;
        RECT 868.180 -240.605 868.560 -136.015 ;
        RECT 869.700 -245.175 870.080 -140.585 ;
        RECT 871.220 -240.605 871.600 -136.015 ;
        RECT 872.740 -245.175 873.120 -140.585 ;
        RECT 874.260 -240.605 874.640 -136.015 ;
        RECT 875.780 -245.175 876.160 -140.585 ;
        RECT 877.300 -240.605 877.680 -136.015 ;
        RECT 878.820 -245.175 879.200 -140.585 ;
        RECT 880.340 -240.605 880.720 -136.015 ;
        RECT 881.860 -245.175 882.240 -140.585 ;
        RECT 883.380 -240.605 883.760 -136.015 ;
        RECT 884.900 -245.175 885.280 -140.585 ;
        RECT 886.420 -240.605 886.800 -136.015 ;
        RECT -544.060 -248.010 891.540 -245.175 ;
        RECT 542.480 -263.180 585.980 -252.860 ;
        RECT -545.580 -266.015 886.800 -263.180 ;
        RECT -572.210 -370.595 -545.890 -270.595 ;
        RECT -572.210 -415.595 -545.930 -370.595 ;
        RECT -545.580 -370.605 -545.200 -266.015 ;
        RECT -544.060 -375.175 -543.680 -270.585 ;
        RECT -542.540 -370.605 -542.160 -266.015 ;
        RECT -541.020 -375.175 -540.640 -270.585 ;
        RECT -539.500 -370.605 -539.120 -266.015 ;
        RECT -537.980 -375.175 -537.600 -270.585 ;
        RECT -536.460 -370.605 -536.080 -266.015 ;
        RECT -534.940 -375.175 -534.560 -270.585 ;
        RECT -533.420 -370.605 -533.040 -266.015 ;
        RECT -531.900 -375.175 -531.520 -270.585 ;
        RECT -530.380 -370.605 -530.000 -266.015 ;
        RECT -528.860 -375.175 -528.480 -270.585 ;
        RECT -527.340 -370.605 -526.960 -266.015 ;
        RECT -525.820 -375.175 -525.440 -270.585 ;
        RECT -524.300 -370.605 -523.920 -266.015 ;
        RECT -522.780 -375.175 -522.400 -270.585 ;
        RECT -521.260 -370.605 -520.880 -266.015 ;
        RECT -519.740 -375.175 -519.360 -270.585 ;
        RECT -518.220 -370.605 -517.840 -266.015 ;
        RECT -516.700 -375.175 -516.320 -270.585 ;
        RECT -515.180 -370.605 -514.800 -266.015 ;
        RECT -513.660 -375.175 -513.280 -270.585 ;
        RECT -512.140 -370.605 -511.760 -266.015 ;
        RECT -510.620 -375.175 -510.240 -270.585 ;
        RECT -509.100 -370.605 -508.720 -266.015 ;
        RECT -507.580 -375.175 -507.200 -270.585 ;
        RECT -506.060 -370.605 -505.680 -266.015 ;
        RECT -504.540 -375.175 -504.160 -270.585 ;
        RECT -503.020 -370.605 -502.640 -266.015 ;
        RECT -501.500 -375.175 -501.120 -270.585 ;
        RECT -499.980 -370.605 -499.600 -266.015 ;
        RECT -498.460 -375.175 -498.080 -270.585 ;
        RECT -496.940 -370.605 -496.560 -266.015 ;
        RECT -495.420 -375.175 -495.040 -270.585 ;
        RECT -493.900 -370.605 -493.520 -266.015 ;
        RECT -492.380 -375.175 -492.000 -270.585 ;
        RECT -490.860 -370.605 -490.480 -266.015 ;
        RECT -489.340 -375.175 -488.960 -270.585 ;
        RECT -487.820 -370.605 -487.440 -266.015 ;
        RECT -486.300 -375.175 -485.920 -270.585 ;
        RECT -484.780 -370.605 -484.400 -266.015 ;
        RECT -483.260 -375.175 -482.880 -270.585 ;
        RECT -481.740 -370.605 -481.360 -266.015 ;
        RECT -480.220 -375.175 -479.840 -270.585 ;
        RECT -478.700 -370.605 -478.320 -266.015 ;
        RECT -477.180 -375.175 -476.800 -270.585 ;
        RECT -475.660 -370.605 -475.280 -266.015 ;
        RECT -474.140 -375.175 -473.760 -270.585 ;
        RECT -472.620 -370.605 -472.240 -266.015 ;
        RECT -471.100 -375.175 -470.720 -270.585 ;
        RECT -469.580 -370.605 -469.200 -266.015 ;
        RECT -468.060 -375.175 -467.680 -270.585 ;
        RECT -466.540 -370.605 -466.160 -266.015 ;
        RECT -465.020 -375.175 -464.640 -270.585 ;
        RECT -463.500 -370.605 -463.120 -266.015 ;
        RECT -461.980 -375.175 -461.600 -270.585 ;
        RECT -460.460 -370.605 -460.080 -266.015 ;
        RECT -458.940 -375.175 -458.560 -270.585 ;
        RECT -457.420 -370.605 -457.040 -266.015 ;
        RECT -455.900 -375.175 -455.520 -270.585 ;
        RECT -454.380 -370.605 -454.000 -266.015 ;
        RECT -452.860 -375.175 -452.480 -270.585 ;
        RECT -451.340 -370.605 -450.960 -266.015 ;
        RECT -449.820 -375.175 -449.440 -270.585 ;
        RECT -448.300 -370.605 -447.920 -266.015 ;
        RECT -446.780 -375.175 -446.400 -270.585 ;
        RECT -445.260 -370.605 -444.880 -266.015 ;
        RECT -443.740 -375.175 -443.360 -270.585 ;
        RECT -442.220 -370.605 -441.840 -266.015 ;
        RECT -440.700 -375.175 -440.320 -270.585 ;
        RECT -439.180 -370.605 -438.800 -266.015 ;
        RECT -437.660 -375.175 -437.280 -270.585 ;
        RECT -436.140 -370.605 -435.760 -266.015 ;
        RECT -434.620 -375.175 -434.240 -270.585 ;
        RECT -433.100 -370.605 -432.720 -266.015 ;
        RECT -431.580 -375.175 -431.200 -270.585 ;
        RECT -430.060 -370.605 -429.680 -266.015 ;
        RECT -428.540 -375.175 -428.160 -270.585 ;
        RECT -427.020 -370.605 -426.640 -266.015 ;
        RECT -425.500 -375.175 -425.120 -270.585 ;
        RECT -423.980 -370.605 -423.600 -266.015 ;
        RECT -422.460 -375.175 -422.080 -270.585 ;
        RECT -420.940 -370.605 -420.560 -266.015 ;
        RECT -419.420 -375.175 -419.040 -270.585 ;
        RECT -417.900 -370.605 -417.520 -266.015 ;
        RECT -416.380 -375.175 -416.000 -270.585 ;
        RECT -414.860 -370.605 -414.480 -266.015 ;
        RECT -413.340 -375.175 -412.960 -270.585 ;
        RECT -411.820 -370.605 -411.440 -266.015 ;
        RECT -410.300 -375.175 -409.920 -270.585 ;
        RECT -408.780 -370.605 -408.400 -266.015 ;
        RECT -407.260 -375.175 -406.880 -270.585 ;
        RECT -405.740 -370.605 -405.360 -266.015 ;
        RECT -404.220 -375.175 -403.840 -270.585 ;
        RECT -402.700 -370.605 -402.320 -266.015 ;
        RECT -401.180 -375.175 -400.800 -270.585 ;
        RECT -399.660 -370.605 -399.280 -266.015 ;
        RECT -398.140 -375.175 -397.760 -270.585 ;
        RECT -396.620 -370.605 -396.240 -266.015 ;
        RECT -395.100 -375.175 -394.720 -270.585 ;
        RECT -393.580 -370.605 -393.200 -266.015 ;
        RECT -385.580 -270.595 -385.200 -266.015 ;
        RECT -386.370 -370.605 -385.200 -270.595 ;
        RECT -384.060 -375.175 -383.680 -270.585 ;
        RECT -382.540 -370.605 -382.160 -266.015 ;
        RECT -381.020 -375.175 -380.640 -270.585 ;
        RECT -379.500 -370.605 -379.120 -266.015 ;
        RECT -377.980 -375.175 -377.600 -270.585 ;
        RECT -376.460 -370.605 -376.080 -266.015 ;
        RECT -374.940 -375.175 -374.560 -270.585 ;
        RECT -373.420 -370.605 -373.040 -266.015 ;
        RECT -371.900 -375.175 -371.520 -270.585 ;
        RECT -370.380 -370.605 -370.000 -266.015 ;
        RECT -368.860 -375.175 -368.480 -270.585 ;
        RECT -367.340 -370.605 -366.960 -266.015 ;
        RECT -365.820 -375.175 -365.440 -270.585 ;
        RECT -364.300 -370.605 -363.920 -266.015 ;
        RECT -362.780 -375.175 -362.400 -270.585 ;
        RECT -361.260 -370.605 -360.880 -266.015 ;
        RECT -359.740 -375.175 -359.360 -270.585 ;
        RECT -358.220 -370.605 -357.840 -266.015 ;
        RECT -356.700 -375.175 -356.320 -270.585 ;
        RECT -355.180 -370.605 -354.800 -266.015 ;
        RECT -353.660 -375.175 -353.280 -270.585 ;
        RECT -352.140 -370.605 -351.760 -266.015 ;
        RECT -350.620 -375.175 -350.240 -270.585 ;
        RECT -349.100 -370.605 -348.720 -266.015 ;
        RECT -347.580 -375.175 -347.200 -270.585 ;
        RECT -346.060 -370.605 -345.680 -266.015 ;
        RECT -344.540 -375.175 -344.160 -270.585 ;
        RECT -343.020 -370.605 -342.640 -266.015 ;
        RECT -341.500 -375.175 -341.120 -270.585 ;
        RECT -339.980 -370.605 -339.600 -266.015 ;
        RECT -338.460 -375.175 -338.080 -270.585 ;
        RECT -336.940 -370.605 -336.560 -266.015 ;
        RECT -335.420 -375.175 -335.040 -270.585 ;
        RECT -333.900 -370.605 -333.520 -266.015 ;
        RECT -332.380 -375.175 -332.000 -270.585 ;
        RECT -330.860 -370.605 -330.480 -266.015 ;
        RECT -329.340 -375.175 -328.960 -270.585 ;
        RECT -327.820 -370.605 -327.440 -266.015 ;
        RECT -326.300 -375.175 -325.920 -270.585 ;
        RECT -324.780 -370.605 -324.400 -266.015 ;
        RECT -323.260 -375.175 -322.880 -270.585 ;
        RECT -321.740 -370.605 -321.360 -266.015 ;
        RECT -320.220 -375.175 -319.840 -270.585 ;
        RECT -318.700 -370.605 -318.320 -266.015 ;
        RECT -317.180 -375.175 -316.800 -270.585 ;
        RECT -315.660 -370.605 -315.280 -266.015 ;
        RECT -314.140 -375.175 -313.760 -270.585 ;
        RECT -312.620 -370.605 -312.240 -266.015 ;
        RECT -311.100 -375.175 -310.720 -270.585 ;
        RECT -309.580 -370.605 -309.200 -266.015 ;
        RECT -308.060 -375.175 -307.680 -270.585 ;
        RECT -306.540 -370.605 -306.160 -266.015 ;
        RECT -305.020 -375.175 -304.640 -270.585 ;
        RECT -303.500 -370.605 -303.120 -266.015 ;
        RECT -301.980 -375.175 -301.600 -270.585 ;
        RECT -300.460 -370.605 -300.080 -266.015 ;
        RECT -298.940 -375.175 -298.560 -270.585 ;
        RECT -297.420 -370.605 -297.040 -266.015 ;
        RECT -295.900 -375.175 -295.520 -270.585 ;
        RECT -294.380 -370.605 -294.000 -266.015 ;
        RECT -292.860 -375.175 -292.480 -270.585 ;
        RECT -291.340 -370.605 -290.960 -266.015 ;
        RECT -289.820 -375.175 -289.440 -270.585 ;
        RECT -288.300 -370.605 -287.920 -266.015 ;
        RECT -286.780 -375.175 -286.400 -270.585 ;
        RECT -285.260 -370.605 -284.880 -266.015 ;
        RECT -283.740 -375.175 -283.360 -270.585 ;
        RECT -282.220 -370.605 -281.840 -266.015 ;
        RECT -280.700 -375.175 -280.320 -270.585 ;
        RECT -279.180 -370.605 -278.800 -266.015 ;
        RECT -277.660 -375.175 -277.280 -270.585 ;
        RECT -276.140 -370.605 -275.760 -266.015 ;
        RECT -274.620 -375.175 -274.240 -270.585 ;
        RECT -273.100 -370.605 -272.720 -266.015 ;
        RECT -271.580 -375.175 -271.200 -270.585 ;
        RECT -270.060 -370.605 -269.680 -266.015 ;
        RECT -268.540 -375.175 -268.160 -270.585 ;
        RECT -267.020 -370.605 -266.640 -266.015 ;
        RECT -265.500 -375.175 -265.120 -270.585 ;
        RECT -263.980 -370.605 -263.600 -266.015 ;
        RECT -262.460 -375.175 -262.080 -270.585 ;
        RECT -260.940 -370.605 -260.560 -266.015 ;
        RECT -259.420 -375.175 -259.040 -270.585 ;
        RECT -257.900 -370.605 -257.520 -266.015 ;
        RECT -256.380 -375.175 -256.000 -270.585 ;
        RECT -254.860 -370.605 -254.480 -266.015 ;
        RECT -253.340 -375.175 -252.960 -270.585 ;
        RECT -251.820 -370.605 -251.440 -266.015 ;
        RECT -250.300 -375.175 -249.920 -270.585 ;
        RECT -248.780 -370.605 -248.400 -266.015 ;
        RECT -247.260 -375.175 -246.880 -270.585 ;
        RECT -245.740 -370.605 -245.360 -266.015 ;
        RECT -244.220 -375.175 -243.840 -270.585 ;
        RECT -242.700 -370.605 -242.320 -266.015 ;
        RECT -241.180 -375.175 -240.800 -270.585 ;
        RECT -239.660 -370.605 -239.280 -266.015 ;
        RECT -238.140 -375.175 -237.760 -270.585 ;
        RECT -236.620 -370.605 -236.240 -266.015 ;
        RECT -235.100 -375.175 -234.720 -270.585 ;
        RECT -233.580 -370.605 -233.200 -266.015 ;
        RECT -225.580 -270.595 -225.200 -266.015 ;
        RECT -226.370 -370.605 -225.200 -270.595 ;
        RECT -224.060 -375.175 -223.680 -270.585 ;
        RECT -222.540 -370.605 -222.160 -266.015 ;
        RECT -221.020 -375.175 -220.640 -270.585 ;
        RECT -219.500 -370.605 -219.120 -266.015 ;
        RECT -217.980 -375.175 -217.600 -270.585 ;
        RECT -216.460 -370.605 -216.080 -266.015 ;
        RECT -214.940 -375.175 -214.560 -270.585 ;
        RECT -213.420 -370.605 -213.040 -266.015 ;
        RECT -211.900 -375.175 -211.520 -270.585 ;
        RECT -210.380 -370.605 -210.000 -266.015 ;
        RECT -208.860 -375.175 -208.480 -270.585 ;
        RECT -207.340 -370.605 -206.960 -266.015 ;
        RECT -205.820 -375.175 -205.440 -270.585 ;
        RECT -204.300 -370.605 -203.920 -266.015 ;
        RECT -202.780 -375.175 -202.400 -270.585 ;
        RECT -201.260 -370.605 -200.880 -266.015 ;
        RECT -199.740 -375.175 -199.360 -270.585 ;
        RECT -198.220 -370.605 -197.840 -266.015 ;
        RECT -196.700 -375.175 -196.320 -270.585 ;
        RECT -195.180 -370.605 -194.800 -266.015 ;
        RECT -193.660 -375.175 -193.280 -270.585 ;
        RECT -192.140 -370.605 -191.760 -266.015 ;
        RECT -190.620 -375.175 -190.240 -270.585 ;
        RECT -189.100 -370.605 -188.720 -266.015 ;
        RECT -187.580 -375.175 -187.200 -270.585 ;
        RECT -186.060 -370.605 -185.680 -266.015 ;
        RECT -184.540 -375.175 -184.160 -270.585 ;
        RECT -183.020 -370.605 -182.640 -266.015 ;
        RECT -181.500 -375.175 -181.120 -270.585 ;
        RECT -179.980 -370.605 -179.600 -266.015 ;
        RECT -178.460 -375.175 -178.080 -270.585 ;
        RECT -176.940 -370.605 -176.560 -266.015 ;
        RECT -175.420 -375.175 -175.040 -270.585 ;
        RECT -173.900 -370.605 -173.520 -266.015 ;
        RECT -172.380 -375.175 -172.000 -270.585 ;
        RECT -170.860 -370.605 -170.480 -266.015 ;
        RECT -169.340 -375.175 -168.960 -270.585 ;
        RECT -167.820 -370.605 -167.440 -266.015 ;
        RECT -166.300 -375.175 -165.920 -270.585 ;
        RECT -164.780 -370.605 -164.400 -266.015 ;
        RECT -163.260 -375.175 -162.880 -270.585 ;
        RECT -161.740 -370.605 -161.360 -266.015 ;
        RECT -160.220 -375.175 -159.840 -270.585 ;
        RECT -158.700 -370.605 -158.320 -266.015 ;
        RECT -157.180 -375.175 -156.800 -270.585 ;
        RECT -155.660 -370.605 -155.280 -266.015 ;
        RECT -154.140 -375.175 -153.760 -270.585 ;
        RECT -152.620 -370.605 -152.240 -266.015 ;
        RECT -151.100 -375.175 -150.720 -270.585 ;
        RECT -149.580 -370.605 -149.200 -266.015 ;
        RECT -148.060 -375.175 -147.680 -270.585 ;
        RECT -146.540 -370.605 -146.160 -266.015 ;
        RECT -145.020 -375.175 -144.640 -270.585 ;
        RECT -143.500 -370.605 -143.120 -266.015 ;
        RECT -141.980 -375.175 -141.600 -270.585 ;
        RECT -140.460 -370.605 -140.080 -266.015 ;
        RECT -138.940 -375.175 -138.560 -270.585 ;
        RECT -137.420 -370.605 -137.040 -266.015 ;
        RECT -135.900 -375.175 -135.520 -270.585 ;
        RECT -134.380 -370.605 -134.000 -266.015 ;
        RECT -132.860 -375.175 -132.480 -270.585 ;
        RECT -131.340 -370.605 -130.960 -266.015 ;
        RECT -129.820 -375.175 -129.440 -270.585 ;
        RECT -128.300 -370.605 -127.920 -266.015 ;
        RECT -126.780 -375.175 -126.400 -270.585 ;
        RECT -125.260 -370.605 -124.880 -266.015 ;
        RECT -123.740 -375.175 -123.360 -270.585 ;
        RECT -122.220 -370.605 -121.840 -266.015 ;
        RECT -120.700 -375.175 -120.320 -270.585 ;
        RECT -119.180 -370.605 -118.800 -266.015 ;
        RECT -117.660 -375.175 -117.280 -270.585 ;
        RECT -116.140 -370.605 -115.760 -266.015 ;
        RECT -114.620 -375.175 -114.240 -270.585 ;
        RECT -113.100 -370.605 -112.720 -266.015 ;
        RECT -111.580 -375.175 -111.200 -270.585 ;
        RECT -110.060 -370.605 -109.680 -266.015 ;
        RECT -108.540 -375.175 -108.160 -270.585 ;
        RECT -107.020 -370.605 -106.640 -266.015 ;
        RECT -105.500 -375.175 -105.120 -270.585 ;
        RECT -103.980 -370.605 -103.600 -266.015 ;
        RECT -102.460 -375.175 -102.080 -270.585 ;
        RECT -100.940 -370.605 -100.560 -266.015 ;
        RECT -99.420 -375.175 -99.040 -270.585 ;
        RECT -97.900 -370.605 -97.520 -266.015 ;
        RECT -96.380 -375.175 -96.000 -270.585 ;
        RECT -94.860 -370.605 -94.480 -266.015 ;
        RECT -93.340 -375.175 -92.960 -270.585 ;
        RECT -91.820 -370.605 -91.440 -266.015 ;
        RECT -90.300 -375.175 -89.920 -270.585 ;
        RECT -88.780 -370.605 -88.400 -266.015 ;
        RECT -87.260 -375.175 -86.880 -270.585 ;
        RECT -85.740 -370.605 -85.360 -266.015 ;
        RECT -84.220 -375.175 -83.840 -270.585 ;
        RECT -82.700 -370.605 -82.320 -266.015 ;
        RECT -81.180 -375.175 -80.800 -270.585 ;
        RECT -79.660 -370.605 -79.280 -266.015 ;
        RECT -78.140 -375.175 -77.760 -270.585 ;
        RECT -76.620 -370.605 -76.240 -266.015 ;
        RECT -75.100 -375.175 -74.720 -270.585 ;
        RECT -73.580 -370.605 -73.200 -266.015 ;
        RECT -65.580 -270.595 -65.200 -266.015 ;
        RECT -66.370 -370.605 -65.200 -270.595 ;
        RECT -64.060 -375.175 -63.680 -270.585 ;
        RECT -62.540 -370.605 -62.160 -266.015 ;
        RECT -61.020 -375.175 -60.640 -270.585 ;
        RECT -59.500 -370.605 -59.120 -266.015 ;
        RECT -57.980 -375.175 -57.600 -270.585 ;
        RECT -56.460 -370.605 -56.080 -266.015 ;
        RECT -54.940 -375.175 -54.560 -270.585 ;
        RECT -53.420 -370.605 -53.040 -266.015 ;
        RECT -51.900 -375.175 -51.520 -270.585 ;
        RECT -50.380 -370.605 -50.000 -266.015 ;
        RECT -48.860 -375.175 -48.480 -270.585 ;
        RECT -47.340 -370.605 -46.960 -266.015 ;
        RECT -45.820 -375.175 -45.440 -270.585 ;
        RECT -44.300 -370.605 -43.920 -266.015 ;
        RECT -42.780 -375.175 -42.400 -270.585 ;
        RECT -41.260 -370.605 -40.880 -266.015 ;
        RECT -39.740 -375.175 -39.360 -270.585 ;
        RECT -38.220 -370.605 -37.840 -266.015 ;
        RECT -36.700 -375.175 -36.320 -270.585 ;
        RECT -35.180 -370.605 -34.800 -266.015 ;
        RECT -33.660 -375.175 -33.280 -270.585 ;
        RECT -32.140 -370.605 -31.760 -266.015 ;
        RECT -30.620 -375.175 -30.240 -270.585 ;
        RECT -29.100 -370.605 -28.720 -266.015 ;
        RECT -27.580 -375.175 -27.200 -270.585 ;
        RECT -26.060 -370.605 -25.680 -266.015 ;
        RECT -24.540 -375.175 -24.160 -270.585 ;
        RECT -23.020 -370.605 -22.640 -266.015 ;
        RECT -21.500 -375.175 -21.120 -270.585 ;
        RECT -19.980 -370.605 -19.600 -266.015 ;
        RECT -18.460 -375.175 -18.080 -270.585 ;
        RECT -16.940 -370.605 -16.560 -266.015 ;
        RECT -15.420 -375.175 -15.040 -270.585 ;
        RECT -13.900 -370.605 -13.520 -266.015 ;
        RECT -12.380 -375.175 -12.000 -270.585 ;
        RECT -10.860 -370.605 -10.480 -266.015 ;
        RECT -9.340 -375.175 -8.960 -270.585 ;
        RECT -7.820 -370.605 -7.440 -266.015 ;
        RECT -6.300 -375.175 -5.920 -270.585 ;
        RECT -4.780 -370.605 -4.400 -266.015 ;
        RECT -3.260 -375.175 -2.880 -270.585 ;
        RECT -1.740 -370.605 -1.360 -266.015 ;
        RECT -0.220 -375.175 0.160 -270.585 ;
        RECT 1.300 -370.605 1.680 -266.015 ;
        RECT 2.820 -375.175 3.200 -270.585 ;
        RECT 4.340 -370.605 4.720 -266.015 ;
        RECT 5.860 -375.175 6.240 -270.585 ;
        RECT 7.380 -370.605 7.760 -266.015 ;
        RECT 8.900 -375.175 9.280 -270.585 ;
        RECT 10.420 -370.605 10.800 -266.015 ;
        RECT 11.940 -375.175 12.320 -270.585 ;
        RECT 13.460 -370.605 13.840 -266.015 ;
        RECT 14.980 -375.175 15.360 -270.585 ;
        RECT 16.500 -370.605 16.880 -266.015 ;
        RECT 18.020 -375.175 18.400 -270.585 ;
        RECT 19.540 -370.605 19.920 -266.015 ;
        RECT 21.060 -375.175 21.440 -270.585 ;
        RECT 22.580 -370.605 22.960 -266.015 ;
        RECT 24.100 -375.175 24.480 -270.585 ;
        RECT 25.620 -370.605 26.000 -266.015 ;
        RECT 27.140 -375.175 27.520 -270.585 ;
        RECT 28.660 -370.605 29.040 -266.015 ;
        RECT 30.180 -375.175 30.560 -270.585 ;
        RECT 31.700 -370.605 32.080 -266.015 ;
        RECT 33.220 -375.175 33.600 -270.585 ;
        RECT 34.740 -370.605 35.120 -266.015 ;
        RECT 36.260 -375.175 36.640 -270.585 ;
        RECT 37.780 -370.605 38.160 -266.015 ;
        RECT 39.300 -375.175 39.680 -270.585 ;
        RECT 40.820 -370.605 41.200 -266.015 ;
        RECT 42.340 -375.175 42.720 -270.585 ;
        RECT 43.860 -370.605 44.240 -266.015 ;
        RECT 45.380 -375.175 45.760 -270.585 ;
        RECT 46.900 -370.605 47.280 -266.015 ;
        RECT 48.420 -375.175 48.800 -270.585 ;
        RECT 49.940 -370.605 50.320 -266.015 ;
        RECT 51.460 -375.175 51.840 -270.585 ;
        RECT 52.980 -370.605 53.360 -266.015 ;
        RECT 54.500 -375.175 54.880 -270.585 ;
        RECT 56.020 -370.605 56.400 -266.015 ;
        RECT 57.540 -375.175 57.920 -270.585 ;
        RECT 59.060 -370.605 59.440 -266.015 ;
        RECT 60.580 -375.175 60.960 -270.585 ;
        RECT 62.100 -370.605 62.480 -266.015 ;
        RECT 63.620 -375.175 64.000 -270.585 ;
        RECT 65.140 -370.605 65.520 -266.015 ;
        RECT 66.660 -375.175 67.040 -270.585 ;
        RECT 68.180 -370.605 68.560 -266.015 ;
        RECT 69.700 -375.175 70.080 -270.585 ;
        RECT 71.220 -370.605 71.600 -266.015 ;
        RECT 72.740 -375.175 73.120 -270.585 ;
        RECT 74.260 -370.605 74.640 -266.015 ;
        RECT 75.780 -375.175 76.160 -270.585 ;
        RECT 77.300 -370.605 77.680 -266.015 ;
        RECT 78.820 -375.175 79.200 -270.585 ;
        RECT 80.340 -370.605 80.720 -266.015 ;
        RECT 81.860 -375.175 82.240 -270.585 ;
        RECT 83.380 -370.605 83.760 -266.015 ;
        RECT 84.900 -375.175 85.280 -270.585 ;
        RECT 86.420 -370.605 86.800 -266.015 ;
        RECT 94.420 -270.595 94.800 -266.015 ;
        RECT 93.630 -370.605 94.800 -270.595 ;
        RECT 95.940 -375.175 96.320 -270.585 ;
        RECT 97.460 -370.605 97.840 -266.015 ;
        RECT 98.980 -375.175 99.360 -270.585 ;
        RECT 100.500 -370.605 100.880 -266.015 ;
        RECT 102.020 -375.175 102.400 -270.585 ;
        RECT 103.540 -370.605 103.920 -266.015 ;
        RECT 105.060 -375.175 105.440 -270.585 ;
        RECT 106.580 -370.605 106.960 -266.015 ;
        RECT 108.100 -375.175 108.480 -270.585 ;
        RECT 109.620 -370.605 110.000 -266.015 ;
        RECT 111.140 -375.175 111.520 -270.585 ;
        RECT 112.660 -370.605 113.040 -266.015 ;
        RECT 114.180 -375.175 114.560 -270.585 ;
        RECT 115.700 -370.605 116.080 -266.015 ;
        RECT 117.220 -375.175 117.600 -270.585 ;
        RECT 118.740 -370.605 119.120 -266.015 ;
        RECT 120.260 -375.175 120.640 -270.585 ;
        RECT 121.780 -370.605 122.160 -266.015 ;
        RECT 123.300 -375.175 123.680 -270.585 ;
        RECT 124.820 -370.605 125.200 -266.015 ;
        RECT 126.340 -375.175 126.720 -270.585 ;
        RECT 127.860 -370.605 128.240 -266.015 ;
        RECT 129.380 -375.175 129.760 -270.585 ;
        RECT 130.900 -370.605 131.280 -266.015 ;
        RECT 132.420 -375.175 132.800 -270.585 ;
        RECT 133.940 -370.605 134.320 -266.015 ;
        RECT 135.460 -375.175 135.840 -270.585 ;
        RECT 136.980 -370.605 137.360 -266.015 ;
        RECT 138.500 -375.175 138.880 -270.585 ;
        RECT 140.020 -370.605 140.400 -266.015 ;
        RECT 141.540 -375.175 141.920 -270.585 ;
        RECT 143.060 -370.605 143.440 -266.015 ;
        RECT 144.580 -375.175 144.960 -270.585 ;
        RECT 146.100 -370.605 146.480 -266.015 ;
        RECT 147.620 -375.175 148.000 -270.585 ;
        RECT 149.140 -370.605 149.520 -266.015 ;
        RECT 150.660 -375.175 151.040 -270.585 ;
        RECT 152.180 -370.605 152.560 -266.015 ;
        RECT 153.700 -375.175 154.080 -270.585 ;
        RECT 155.220 -370.605 155.600 -266.015 ;
        RECT 156.740 -375.175 157.120 -270.585 ;
        RECT 158.260 -370.605 158.640 -266.015 ;
        RECT 159.780 -375.175 160.160 -270.585 ;
        RECT 161.300 -370.605 161.680 -266.015 ;
        RECT 162.820 -375.175 163.200 -270.585 ;
        RECT 164.340 -370.605 164.720 -266.015 ;
        RECT 165.860 -375.175 166.240 -270.585 ;
        RECT 167.380 -370.605 167.760 -266.015 ;
        RECT 168.900 -375.175 169.280 -270.585 ;
        RECT 170.420 -370.605 170.800 -266.015 ;
        RECT 171.940 -375.175 172.320 -270.585 ;
        RECT 173.460 -370.605 173.840 -266.015 ;
        RECT 174.980 -375.175 175.360 -270.585 ;
        RECT 176.500 -370.605 176.880 -266.015 ;
        RECT 178.020 -375.175 178.400 -270.585 ;
        RECT 179.540 -370.605 179.920 -266.015 ;
        RECT 181.060 -375.175 181.440 -270.585 ;
        RECT 182.580 -370.605 182.960 -266.015 ;
        RECT 184.100 -375.175 184.480 -270.585 ;
        RECT 185.620 -370.605 186.000 -266.015 ;
        RECT 187.140 -375.175 187.520 -270.585 ;
        RECT 188.660 -370.605 189.040 -266.015 ;
        RECT 190.180 -375.175 190.560 -270.585 ;
        RECT 191.700 -370.605 192.080 -266.015 ;
        RECT 193.220 -375.175 193.600 -270.585 ;
        RECT 194.740 -370.605 195.120 -266.015 ;
        RECT 196.260 -375.175 196.640 -270.585 ;
        RECT 197.780 -370.605 198.160 -266.015 ;
        RECT 199.300 -375.175 199.680 -270.585 ;
        RECT 200.820 -370.605 201.200 -266.015 ;
        RECT 202.340 -375.175 202.720 -270.585 ;
        RECT 203.860 -370.605 204.240 -266.015 ;
        RECT 205.380 -375.175 205.760 -270.585 ;
        RECT 206.900 -370.605 207.280 -266.015 ;
        RECT 208.420 -375.175 208.800 -270.585 ;
        RECT 209.940 -370.605 210.320 -266.015 ;
        RECT 211.460 -375.175 211.840 -270.585 ;
        RECT 212.980 -370.605 213.360 -266.015 ;
        RECT 214.500 -375.175 214.880 -270.585 ;
        RECT 216.020 -370.605 216.400 -266.015 ;
        RECT 217.540 -375.175 217.920 -270.585 ;
        RECT 219.060 -370.605 219.440 -266.015 ;
        RECT 220.580 -375.175 220.960 -270.585 ;
        RECT 222.100 -370.605 222.480 -266.015 ;
        RECT 223.620 -375.175 224.000 -270.585 ;
        RECT 225.140 -370.605 225.520 -266.015 ;
        RECT 226.660 -375.175 227.040 -270.585 ;
        RECT 228.180 -370.605 228.560 -266.015 ;
        RECT 229.700 -375.175 230.080 -270.585 ;
        RECT 231.220 -370.605 231.600 -266.015 ;
        RECT 232.740 -375.175 233.120 -270.585 ;
        RECT 234.260 -370.605 234.640 -266.015 ;
        RECT 235.780 -375.175 236.160 -270.585 ;
        RECT 237.300 -370.605 237.680 -266.015 ;
        RECT 238.820 -375.175 239.200 -270.585 ;
        RECT 240.340 -370.605 240.720 -266.015 ;
        RECT 241.860 -375.175 242.240 -270.585 ;
        RECT 243.380 -370.605 243.760 -266.015 ;
        RECT 244.900 -375.175 245.280 -270.585 ;
        RECT 246.420 -370.605 246.800 -266.015 ;
        RECT 254.420 -270.595 254.800 -266.015 ;
        RECT 253.630 -370.605 254.800 -270.595 ;
        RECT 255.940 -375.175 256.320 -270.585 ;
        RECT 257.460 -370.605 257.840 -266.015 ;
        RECT 258.980 -375.175 259.360 -270.585 ;
        RECT 260.500 -370.605 260.880 -266.015 ;
        RECT 262.020 -375.175 262.400 -270.585 ;
        RECT 263.540 -370.605 263.920 -266.015 ;
        RECT 265.060 -375.175 265.440 -270.585 ;
        RECT 266.580 -370.605 266.960 -266.015 ;
        RECT 268.100 -375.175 268.480 -270.585 ;
        RECT 269.620 -370.605 270.000 -266.015 ;
        RECT 271.140 -375.175 271.520 -270.585 ;
        RECT 272.660 -370.605 273.040 -266.015 ;
        RECT 274.180 -375.175 274.560 -270.585 ;
        RECT 275.700 -370.605 276.080 -266.015 ;
        RECT 277.220 -375.175 277.600 -270.585 ;
        RECT 278.740 -370.605 279.120 -266.015 ;
        RECT 280.260 -375.175 280.640 -270.585 ;
        RECT 281.780 -370.605 282.160 -266.015 ;
        RECT 283.300 -375.175 283.680 -270.585 ;
        RECT 284.820 -370.605 285.200 -266.015 ;
        RECT 286.340 -375.175 286.720 -270.585 ;
        RECT 287.860 -370.605 288.240 -266.015 ;
        RECT 289.380 -375.175 289.760 -270.585 ;
        RECT 290.900 -370.605 291.280 -266.015 ;
        RECT 292.420 -375.175 292.800 -270.585 ;
        RECT 293.940 -370.605 294.320 -266.015 ;
        RECT 295.460 -375.175 295.840 -270.585 ;
        RECT 296.980 -370.605 297.360 -266.015 ;
        RECT 298.500 -375.175 298.880 -270.585 ;
        RECT 300.020 -370.605 300.400 -266.015 ;
        RECT 301.540 -375.175 301.920 -270.585 ;
        RECT 303.060 -370.605 303.440 -266.015 ;
        RECT 304.580 -375.175 304.960 -270.585 ;
        RECT 306.100 -370.605 306.480 -266.015 ;
        RECT 307.620 -375.175 308.000 -270.585 ;
        RECT 309.140 -370.605 309.520 -266.015 ;
        RECT 310.660 -375.175 311.040 -270.585 ;
        RECT 312.180 -370.605 312.560 -266.015 ;
        RECT 313.700 -375.175 314.080 -270.585 ;
        RECT 315.220 -370.605 315.600 -266.015 ;
        RECT 316.740 -375.175 317.120 -270.585 ;
        RECT 318.260 -370.605 318.640 -266.015 ;
        RECT 319.780 -375.175 320.160 -270.585 ;
        RECT 321.300 -370.605 321.680 -266.015 ;
        RECT 322.820 -375.175 323.200 -270.585 ;
        RECT 324.340 -370.605 324.720 -266.015 ;
        RECT 325.860 -375.175 326.240 -270.585 ;
        RECT 327.380 -370.605 327.760 -266.015 ;
        RECT 328.900 -375.175 329.280 -270.585 ;
        RECT 330.420 -370.605 330.800 -266.015 ;
        RECT 331.940 -375.175 332.320 -270.585 ;
        RECT 333.460 -370.605 333.840 -266.015 ;
        RECT 334.980 -375.175 335.360 -270.585 ;
        RECT 336.500 -370.605 336.880 -266.015 ;
        RECT 338.020 -375.175 338.400 -270.585 ;
        RECT 339.540 -370.605 339.920 -266.015 ;
        RECT 341.060 -375.175 341.440 -270.585 ;
        RECT 342.580 -370.605 342.960 -266.015 ;
        RECT 344.100 -375.175 344.480 -270.585 ;
        RECT 345.620 -370.605 346.000 -266.015 ;
        RECT 347.140 -375.175 347.520 -270.585 ;
        RECT 348.660 -370.605 349.040 -266.015 ;
        RECT 350.180 -375.175 350.560 -270.585 ;
        RECT 351.700 -370.605 352.080 -266.015 ;
        RECT 353.220 -375.175 353.600 -270.585 ;
        RECT 354.740 -370.605 355.120 -266.015 ;
        RECT 356.260 -375.175 356.640 -270.585 ;
        RECT 357.780 -370.605 358.160 -266.015 ;
        RECT 359.300 -375.175 359.680 -270.585 ;
        RECT 360.820 -370.605 361.200 -266.015 ;
        RECT 362.340 -375.175 362.720 -270.585 ;
        RECT 363.860 -370.605 364.240 -266.015 ;
        RECT 365.380 -375.175 365.760 -270.585 ;
        RECT 366.900 -370.605 367.280 -266.015 ;
        RECT 368.420 -375.175 368.800 -270.585 ;
        RECT 369.940 -370.605 370.320 -266.015 ;
        RECT 371.460 -375.175 371.840 -270.585 ;
        RECT 372.980 -370.605 373.360 -266.015 ;
        RECT 374.500 -375.175 374.880 -270.585 ;
        RECT 376.020 -370.605 376.400 -266.015 ;
        RECT 377.540 -375.175 377.920 -270.585 ;
        RECT 379.060 -370.605 379.440 -266.015 ;
        RECT 380.580 -375.175 380.960 -270.585 ;
        RECT 382.100 -370.605 382.480 -266.015 ;
        RECT 383.620 -375.175 384.000 -270.585 ;
        RECT 385.140 -370.605 385.520 -266.015 ;
        RECT 386.660 -375.175 387.040 -270.585 ;
        RECT 388.180 -370.605 388.560 -266.015 ;
        RECT 389.700 -375.175 390.080 -270.585 ;
        RECT 391.220 -370.605 391.600 -266.015 ;
        RECT 392.740 -375.175 393.120 -270.585 ;
        RECT 394.260 -370.605 394.640 -266.015 ;
        RECT 395.780 -375.175 396.160 -270.585 ;
        RECT 397.300 -370.605 397.680 -266.015 ;
        RECT 398.820 -375.175 399.200 -270.585 ;
        RECT 400.340 -370.605 400.720 -266.015 ;
        RECT 401.860 -375.175 402.240 -270.585 ;
        RECT 403.380 -370.605 403.760 -266.015 ;
        RECT 404.900 -375.175 405.280 -270.585 ;
        RECT 406.420 -370.605 406.800 -266.015 ;
        RECT 414.420 -270.595 414.800 -266.015 ;
        RECT 413.630 -370.605 414.800 -270.595 ;
        RECT 415.940 -375.175 416.320 -270.585 ;
        RECT 417.460 -370.605 417.840 -266.015 ;
        RECT 418.980 -375.175 419.360 -270.585 ;
        RECT 420.500 -370.605 420.880 -266.015 ;
        RECT 422.020 -375.175 422.400 -270.585 ;
        RECT 423.540 -370.605 423.920 -266.015 ;
        RECT 425.060 -375.175 425.440 -270.585 ;
        RECT 426.580 -370.605 426.960 -266.015 ;
        RECT 428.100 -375.175 428.480 -270.585 ;
        RECT 429.620 -370.605 430.000 -266.015 ;
        RECT 431.140 -375.175 431.520 -270.585 ;
        RECT 432.660 -370.605 433.040 -266.015 ;
        RECT 434.180 -375.175 434.560 -270.585 ;
        RECT 435.700 -370.605 436.080 -266.015 ;
        RECT 437.220 -375.175 437.600 -270.585 ;
        RECT 438.740 -370.605 439.120 -266.015 ;
        RECT 440.260 -375.175 440.640 -270.585 ;
        RECT 441.780 -370.605 442.160 -266.015 ;
        RECT 443.300 -375.175 443.680 -270.585 ;
        RECT 444.820 -370.605 445.200 -266.015 ;
        RECT 446.340 -375.175 446.720 -270.585 ;
        RECT 447.860 -370.605 448.240 -266.015 ;
        RECT 449.380 -375.175 449.760 -270.585 ;
        RECT 450.900 -370.605 451.280 -266.015 ;
        RECT 452.420 -375.175 452.800 -270.585 ;
        RECT 453.940 -370.605 454.320 -266.015 ;
        RECT 455.460 -375.175 455.840 -270.585 ;
        RECT 456.980 -370.605 457.360 -266.015 ;
        RECT 458.500 -375.175 458.880 -270.585 ;
        RECT 460.020 -370.605 460.400 -266.015 ;
        RECT 461.540 -375.175 461.920 -270.585 ;
        RECT 463.060 -370.605 463.440 -266.015 ;
        RECT 464.580 -375.175 464.960 -270.585 ;
        RECT 466.100 -370.605 466.480 -266.015 ;
        RECT 467.620 -375.175 468.000 -270.585 ;
        RECT 469.140 -370.605 469.520 -266.015 ;
        RECT 470.660 -375.175 471.040 -270.585 ;
        RECT 472.180 -370.605 472.560 -266.015 ;
        RECT 473.700 -375.175 474.080 -270.585 ;
        RECT 475.220 -370.605 475.600 -266.015 ;
        RECT 476.740 -375.175 477.120 -270.585 ;
        RECT 478.260 -370.605 478.640 -266.015 ;
        RECT 479.780 -375.175 480.160 -270.585 ;
        RECT 481.300 -370.605 481.680 -266.015 ;
        RECT 482.820 -375.175 483.200 -270.585 ;
        RECT 484.340 -370.605 484.720 -266.015 ;
        RECT 485.860 -375.175 486.240 -270.585 ;
        RECT 487.380 -370.605 487.760 -266.015 ;
        RECT 488.900 -375.175 489.280 -270.585 ;
        RECT 490.420 -370.605 490.800 -266.015 ;
        RECT 491.940 -375.175 492.320 -270.585 ;
        RECT 493.460 -370.605 493.840 -266.015 ;
        RECT 494.980 -375.175 495.360 -270.585 ;
        RECT 496.500 -370.605 496.880 -266.015 ;
        RECT 498.020 -375.175 498.400 -270.585 ;
        RECT 499.540 -370.605 499.920 -266.015 ;
        RECT 501.060 -375.175 501.440 -270.585 ;
        RECT 502.580 -370.605 502.960 -266.015 ;
        RECT 504.100 -375.175 504.480 -270.585 ;
        RECT 505.620 -370.605 506.000 -266.015 ;
        RECT 507.140 -375.175 507.520 -270.585 ;
        RECT 508.660 -370.605 509.040 -266.015 ;
        RECT 510.180 -375.175 510.560 -270.585 ;
        RECT 511.700 -370.605 512.080 -266.015 ;
        RECT 513.220 -375.175 513.600 -270.585 ;
        RECT 514.740 -370.605 515.120 -266.015 ;
        RECT 516.260 -375.175 516.640 -270.585 ;
        RECT 517.780 -370.605 518.160 -266.015 ;
        RECT 519.300 -375.175 519.680 -270.585 ;
        RECT 520.820 -370.605 521.200 -266.015 ;
        RECT 522.340 -375.175 522.720 -270.585 ;
        RECT 523.860 -370.605 524.240 -266.015 ;
        RECT 525.380 -375.175 525.760 -270.585 ;
        RECT 526.900 -370.605 527.280 -266.015 ;
        RECT 528.420 -375.175 528.800 -270.585 ;
        RECT 529.940 -370.605 530.320 -266.015 ;
        RECT 531.460 -375.175 531.840 -270.585 ;
        RECT 532.980 -370.605 533.360 -266.015 ;
        RECT 534.500 -375.175 534.880 -270.585 ;
        RECT 536.020 -370.605 536.400 -266.015 ;
        RECT 537.540 -375.175 537.920 -270.585 ;
        RECT 539.060 -370.605 539.440 -266.015 ;
        RECT 540.580 -375.175 540.960 -270.585 ;
        RECT 542.100 -370.605 542.480 -266.015 ;
        RECT 543.620 -375.175 544.000 -270.585 ;
        RECT 545.140 -370.605 545.520 -266.015 ;
        RECT 546.660 -375.175 547.040 -270.585 ;
        RECT 548.180 -370.605 548.560 -266.015 ;
        RECT 549.700 -375.175 550.080 -270.585 ;
        RECT 551.220 -370.605 551.600 -266.015 ;
        RECT 552.740 -375.175 553.120 -270.585 ;
        RECT 554.260 -370.605 554.640 -266.015 ;
        RECT 555.780 -375.175 556.160 -270.585 ;
        RECT 557.300 -370.605 557.680 -266.015 ;
        RECT 558.820 -375.175 559.200 -270.585 ;
        RECT 560.340 -370.605 560.720 -266.015 ;
        RECT 561.860 -375.175 562.240 -270.585 ;
        RECT 563.380 -370.605 563.760 -266.015 ;
        RECT 564.900 -375.175 565.280 -270.585 ;
        RECT 566.420 -370.605 566.800 -266.015 ;
        RECT 574.420 -270.595 574.800 -266.015 ;
        RECT 573.630 -370.605 574.800 -270.595 ;
        RECT 575.940 -375.175 576.320 -270.585 ;
        RECT 577.460 -370.605 577.840 -266.015 ;
        RECT 578.980 -375.175 579.360 -270.585 ;
        RECT 580.500 -370.605 580.880 -266.015 ;
        RECT 582.020 -375.175 582.400 -270.585 ;
        RECT 583.540 -370.605 583.920 -266.015 ;
        RECT 585.060 -375.175 585.440 -270.585 ;
        RECT 586.580 -370.605 586.960 -266.015 ;
        RECT 588.100 -375.175 588.480 -270.585 ;
        RECT 589.620 -370.605 590.000 -266.015 ;
        RECT 591.140 -375.175 591.520 -270.585 ;
        RECT 592.660 -370.605 593.040 -266.015 ;
        RECT 594.180 -375.175 594.560 -270.585 ;
        RECT 595.700 -370.605 596.080 -266.015 ;
        RECT 597.220 -375.175 597.600 -270.585 ;
        RECT 598.740 -370.605 599.120 -266.015 ;
        RECT 600.260 -375.175 600.640 -270.585 ;
        RECT 601.780 -370.605 602.160 -266.015 ;
        RECT 603.300 -375.175 603.680 -270.585 ;
        RECT 604.820 -370.605 605.200 -266.015 ;
        RECT 606.340 -375.175 606.720 -270.585 ;
        RECT 607.860 -370.605 608.240 -266.015 ;
        RECT 609.380 -375.175 609.760 -270.585 ;
        RECT 610.900 -370.605 611.280 -266.015 ;
        RECT 612.420 -375.175 612.800 -270.585 ;
        RECT 613.940 -370.605 614.320 -266.015 ;
        RECT 615.460 -375.175 615.840 -270.585 ;
        RECT 616.980 -370.605 617.360 -266.015 ;
        RECT 618.500 -375.175 618.880 -270.585 ;
        RECT 620.020 -370.605 620.400 -266.015 ;
        RECT 621.540 -375.175 621.920 -270.585 ;
        RECT 623.060 -370.605 623.440 -266.015 ;
        RECT 624.580 -375.175 624.960 -270.585 ;
        RECT 626.100 -370.605 626.480 -266.015 ;
        RECT 627.620 -375.175 628.000 -270.585 ;
        RECT 629.140 -370.605 629.520 -266.015 ;
        RECT 630.660 -375.175 631.040 -270.585 ;
        RECT 632.180 -370.605 632.560 -266.015 ;
        RECT 633.700 -375.175 634.080 -270.585 ;
        RECT 635.220 -370.605 635.600 -266.015 ;
        RECT 636.740 -375.175 637.120 -270.585 ;
        RECT 638.260 -370.605 638.640 -266.015 ;
        RECT 639.780 -375.175 640.160 -270.585 ;
        RECT 641.300 -370.605 641.680 -266.015 ;
        RECT 642.820 -375.175 643.200 -270.585 ;
        RECT 644.340 -370.605 644.720 -266.015 ;
        RECT 645.860 -375.175 646.240 -270.585 ;
        RECT 647.380 -370.605 647.760 -266.015 ;
        RECT 648.900 -375.175 649.280 -270.585 ;
        RECT 650.420 -370.605 650.800 -266.015 ;
        RECT 651.940 -375.175 652.320 -270.585 ;
        RECT 653.460 -370.605 653.840 -266.015 ;
        RECT 654.980 -375.175 655.360 -270.585 ;
        RECT 656.500 -370.605 656.880 -266.015 ;
        RECT 658.020 -375.175 658.400 -270.585 ;
        RECT 659.540 -370.605 659.920 -266.015 ;
        RECT 661.060 -375.175 661.440 -270.585 ;
        RECT 662.580 -370.605 662.960 -266.015 ;
        RECT 664.100 -375.175 664.480 -270.585 ;
        RECT 665.620 -370.605 666.000 -266.015 ;
        RECT 667.140 -375.175 667.520 -270.585 ;
        RECT 668.660 -370.605 669.040 -266.015 ;
        RECT 670.180 -375.175 670.560 -270.585 ;
        RECT 671.700 -370.605 672.080 -266.015 ;
        RECT 673.220 -375.175 673.600 -270.585 ;
        RECT 674.740 -370.605 675.120 -266.015 ;
        RECT 676.260 -375.175 676.640 -270.585 ;
        RECT 677.780 -370.605 678.160 -266.015 ;
        RECT 679.300 -375.175 679.680 -270.585 ;
        RECT 680.820 -370.605 681.200 -266.015 ;
        RECT 682.340 -375.175 682.720 -270.585 ;
        RECT 683.860 -370.605 684.240 -266.015 ;
        RECT 685.380 -375.175 685.760 -270.585 ;
        RECT 686.900 -370.605 687.280 -266.015 ;
        RECT 688.420 -375.175 688.800 -270.585 ;
        RECT 689.940 -370.605 690.320 -266.015 ;
        RECT 691.460 -375.175 691.840 -270.585 ;
        RECT 692.980 -370.605 693.360 -266.015 ;
        RECT 694.500 -375.175 694.880 -270.585 ;
        RECT 696.020 -370.605 696.400 -266.015 ;
        RECT 697.540 -375.175 697.920 -270.585 ;
        RECT 699.060 -370.605 699.440 -266.015 ;
        RECT 700.580 -375.175 700.960 -270.585 ;
        RECT 702.100 -370.605 702.480 -266.015 ;
        RECT 703.620 -375.175 704.000 -270.585 ;
        RECT 705.140 -370.605 705.520 -266.015 ;
        RECT 706.660 -375.175 707.040 -270.585 ;
        RECT 708.180 -370.605 708.560 -266.015 ;
        RECT 709.700 -375.175 710.080 -270.585 ;
        RECT 711.220 -370.605 711.600 -266.015 ;
        RECT 712.740 -375.175 713.120 -270.585 ;
        RECT 714.260 -370.605 714.640 -266.015 ;
        RECT 715.780 -375.175 716.160 -270.585 ;
        RECT 717.300 -370.605 717.680 -266.015 ;
        RECT 718.820 -375.175 719.200 -270.585 ;
        RECT 720.340 -370.605 720.720 -266.015 ;
        RECT 721.860 -375.175 722.240 -270.585 ;
        RECT 723.380 -370.605 723.760 -266.015 ;
        RECT 724.900 -375.175 725.280 -270.585 ;
        RECT 726.420 -370.605 726.800 -266.015 ;
        RECT 734.420 -270.595 734.800 -266.015 ;
        RECT 733.630 -370.605 734.800 -270.595 ;
        RECT 735.940 -375.175 736.320 -270.585 ;
        RECT 737.460 -370.605 737.840 -266.015 ;
        RECT 738.980 -375.175 739.360 -270.585 ;
        RECT 740.500 -370.605 740.880 -266.015 ;
        RECT 742.020 -375.175 742.400 -270.585 ;
        RECT 743.540 -370.605 743.920 -266.015 ;
        RECT 745.060 -375.175 745.440 -270.585 ;
        RECT 746.580 -370.605 746.960 -266.015 ;
        RECT 748.100 -375.175 748.480 -270.585 ;
        RECT 749.620 -370.605 750.000 -266.015 ;
        RECT 751.140 -375.175 751.520 -270.585 ;
        RECT 752.660 -370.605 753.040 -266.015 ;
        RECT 754.180 -375.175 754.560 -270.585 ;
        RECT 755.700 -370.605 756.080 -266.015 ;
        RECT 757.220 -375.175 757.600 -270.585 ;
        RECT 758.740 -370.605 759.120 -266.015 ;
        RECT 760.260 -375.175 760.640 -270.585 ;
        RECT 761.780 -370.605 762.160 -266.015 ;
        RECT 763.300 -375.175 763.680 -270.585 ;
        RECT 764.820 -370.605 765.200 -266.015 ;
        RECT 766.340 -375.175 766.720 -270.585 ;
        RECT 767.860 -370.605 768.240 -266.015 ;
        RECT 769.380 -375.175 769.760 -270.585 ;
        RECT 770.900 -370.605 771.280 -266.015 ;
        RECT 772.420 -375.175 772.800 -270.585 ;
        RECT 773.940 -370.605 774.320 -266.015 ;
        RECT 775.460 -375.175 775.840 -270.585 ;
        RECT 776.980 -370.605 777.360 -266.015 ;
        RECT 778.500 -375.175 778.880 -270.585 ;
        RECT 780.020 -370.605 780.400 -266.015 ;
        RECT 781.540 -375.175 781.920 -270.585 ;
        RECT 783.060 -370.605 783.440 -266.015 ;
        RECT 784.580 -375.175 784.960 -270.585 ;
        RECT 786.100 -370.605 786.480 -266.015 ;
        RECT 787.620 -375.175 788.000 -270.585 ;
        RECT 789.140 -370.605 789.520 -266.015 ;
        RECT 790.660 -375.175 791.040 -270.585 ;
        RECT 792.180 -370.605 792.560 -266.015 ;
        RECT 793.700 -375.175 794.080 -270.585 ;
        RECT 795.220 -370.605 795.600 -266.015 ;
        RECT 796.740 -375.175 797.120 -270.585 ;
        RECT 798.260 -370.605 798.640 -266.015 ;
        RECT 799.780 -375.175 800.160 -270.585 ;
        RECT 801.300 -370.605 801.680 -266.015 ;
        RECT 802.820 -375.175 803.200 -270.585 ;
        RECT 804.340 -370.605 804.720 -266.015 ;
        RECT 805.860 -375.175 806.240 -270.585 ;
        RECT 807.380 -370.605 807.760 -266.015 ;
        RECT 808.900 -375.175 809.280 -270.585 ;
        RECT 810.420 -370.605 810.800 -266.015 ;
        RECT 811.940 -375.175 812.320 -270.585 ;
        RECT 813.460 -370.605 813.840 -266.015 ;
        RECT 814.980 -375.175 815.360 -270.585 ;
        RECT 816.500 -370.605 816.880 -266.015 ;
        RECT 818.020 -375.175 818.400 -270.585 ;
        RECT 819.540 -370.605 819.920 -266.015 ;
        RECT 821.060 -375.175 821.440 -270.585 ;
        RECT 822.580 -370.605 822.960 -266.015 ;
        RECT 824.100 -375.175 824.480 -270.585 ;
        RECT 825.620 -370.605 826.000 -266.015 ;
        RECT 827.140 -375.175 827.520 -270.585 ;
        RECT 828.660 -370.605 829.040 -266.015 ;
        RECT 830.180 -375.175 830.560 -270.585 ;
        RECT 831.700 -370.605 832.080 -266.015 ;
        RECT 833.220 -375.175 833.600 -270.585 ;
        RECT 834.740 -370.605 835.120 -266.015 ;
        RECT 836.260 -375.175 836.640 -270.585 ;
        RECT 837.780 -370.605 838.160 -266.015 ;
        RECT 839.300 -375.175 839.680 -270.585 ;
        RECT 840.820 -370.605 841.200 -266.015 ;
        RECT 842.340 -375.175 842.720 -270.585 ;
        RECT 843.860 -370.605 844.240 -266.015 ;
        RECT 845.380 -375.175 845.760 -270.585 ;
        RECT 846.900 -370.605 847.280 -266.015 ;
        RECT 848.420 -375.175 848.800 -270.585 ;
        RECT 849.940 -370.605 850.320 -266.015 ;
        RECT 851.460 -375.175 851.840 -270.585 ;
        RECT 852.980 -370.605 853.360 -266.015 ;
        RECT 854.500 -375.175 854.880 -270.585 ;
        RECT 856.020 -370.605 856.400 -266.015 ;
        RECT 857.540 -375.175 857.920 -270.585 ;
        RECT 859.060 -370.605 859.440 -266.015 ;
        RECT 860.580 -375.175 860.960 -270.585 ;
        RECT 862.100 -370.605 862.480 -266.015 ;
        RECT 863.620 -375.175 864.000 -270.585 ;
        RECT 865.140 -370.605 865.520 -266.015 ;
        RECT 866.660 -375.175 867.040 -270.585 ;
        RECT 868.180 -370.605 868.560 -266.015 ;
        RECT 869.700 -375.175 870.080 -270.585 ;
        RECT 871.220 -370.605 871.600 -266.015 ;
        RECT 872.740 -375.175 873.120 -270.585 ;
        RECT 874.260 -370.605 874.640 -266.015 ;
        RECT 875.780 -375.175 876.160 -270.585 ;
        RECT 877.300 -370.605 877.680 -266.015 ;
        RECT 878.820 -375.175 879.200 -270.585 ;
        RECT 880.340 -370.605 880.720 -266.015 ;
        RECT 881.860 -375.175 882.240 -270.585 ;
        RECT 883.380 -370.605 883.760 -266.015 ;
        RECT 884.900 -375.175 885.280 -270.585 ;
        RECT 886.420 -370.605 886.800 -266.015 ;
        RECT 888.320 -375.175 891.540 -248.010 ;
        RECT -544.060 -378.010 891.540 -375.175 ;
        RECT -544.060 -384.605 888.320 -378.010 ;
        RECT -545.580 -411.015 886.800 -401.350 ;
        RECT -572.210 -515.595 -545.890 -415.595 ;
        RECT -572.210 -545.595 -545.930 -515.595 ;
        RECT -545.580 -515.605 -545.200 -411.015 ;
        RECT -544.060 -520.175 -543.680 -415.585 ;
        RECT -542.540 -515.605 -542.160 -411.015 ;
        RECT -541.020 -520.175 -540.640 -415.585 ;
        RECT -539.500 -515.605 -539.120 -411.015 ;
        RECT -537.980 -520.175 -537.600 -415.585 ;
        RECT -536.460 -515.605 -536.080 -411.015 ;
        RECT -534.940 -520.175 -534.560 -415.585 ;
        RECT -533.420 -515.605 -533.040 -411.015 ;
        RECT -531.900 -520.175 -531.520 -415.585 ;
        RECT -530.380 -515.605 -530.000 -411.015 ;
        RECT -528.860 -520.175 -528.480 -415.585 ;
        RECT -527.340 -515.605 -526.960 -411.015 ;
        RECT -525.820 -520.175 -525.440 -415.585 ;
        RECT -524.300 -515.605 -523.920 -411.015 ;
        RECT -522.780 -520.175 -522.400 -415.585 ;
        RECT -521.260 -515.605 -520.880 -411.015 ;
        RECT -519.740 -520.175 -519.360 -415.585 ;
        RECT -518.220 -515.605 -517.840 -411.015 ;
        RECT -516.700 -520.175 -516.320 -415.585 ;
        RECT -515.180 -515.605 -514.800 -411.015 ;
        RECT -513.660 -520.175 -513.280 -415.585 ;
        RECT -512.140 -515.605 -511.760 -411.015 ;
        RECT -510.620 -520.175 -510.240 -415.585 ;
        RECT -509.100 -515.605 -508.720 -411.015 ;
        RECT -507.580 -520.175 -507.200 -415.585 ;
        RECT -506.060 -515.605 -505.680 -411.015 ;
        RECT -504.540 -520.175 -504.160 -415.585 ;
        RECT -503.020 -515.605 -502.640 -411.015 ;
        RECT -501.500 -520.175 -501.120 -415.585 ;
        RECT -499.980 -515.605 -499.600 -411.015 ;
        RECT -498.460 -520.175 -498.080 -415.585 ;
        RECT -496.940 -515.605 -496.560 -411.015 ;
        RECT -495.420 -520.175 -495.040 -415.585 ;
        RECT -493.900 -515.605 -493.520 -411.015 ;
        RECT -492.380 -520.175 -492.000 -415.585 ;
        RECT -490.860 -515.605 -490.480 -411.015 ;
        RECT -489.340 -520.175 -488.960 -415.585 ;
        RECT -487.820 -515.605 -487.440 -411.015 ;
        RECT -486.300 -520.175 -485.920 -415.585 ;
        RECT -484.780 -515.605 -484.400 -411.015 ;
        RECT -483.260 -520.175 -482.880 -415.585 ;
        RECT -481.740 -515.605 -481.360 -411.015 ;
        RECT -480.220 -520.175 -479.840 -415.585 ;
        RECT -478.700 -515.605 -478.320 -411.015 ;
        RECT -477.180 -520.175 -476.800 -415.585 ;
        RECT -475.660 -515.605 -475.280 -411.015 ;
        RECT -474.140 -520.175 -473.760 -415.585 ;
        RECT -472.620 -515.605 -472.240 -411.015 ;
        RECT -471.100 -520.175 -470.720 -415.585 ;
        RECT -469.580 -515.605 -469.200 -411.015 ;
        RECT -468.060 -520.175 -467.680 -415.585 ;
        RECT -466.540 -515.605 -466.160 -411.015 ;
        RECT -465.020 -520.175 -464.640 -415.585 ;
        RECT -463.500 -515.605 -463.120 -411.015 ;
        RECT -461.980 -520.175 -461.600 -415.585 ;
        RECT -460.460 -515.605 -460.080 -411.015 ;
        RECT -458.940 -520.175 -458.560 -415.585 ;
        RECT -457.420 -515.605 -457.040 -411.015 ;
        RECT -455.900 -520.175 -455.520 -415.585 ;
        RECT -454.380 -515.605 -454.000 -411.015 ;
        RECT -452.860 -520.175 -452.480 -415.585 ;
        RECT -451.340 -515.605 -450.960 -411.015 ;
        RECT -449.820 -520.175 -449.440 -415.585 ;
        RECT -448.300 -515.605 -447.920 -411.015 ;
        RECT -446.780 -520.175 -446.400 -415.585 ;
        RECT -445.260 -515.605 -444.880 -411.015 ;
        RECT -443.740 -520.175 -443.360 -415.585 ;
        RECT -442.220 -515.605 -441.840 -411.015 ;
        RECT -440.700 -520.175 -440.320 -415.585 ;
        RECT -439.180 -515.605 -438.800 -411.015 ;
        RECT -437.660 -520.175 -437.280 -415.585 ;
        RECT -436.140 -515.605 -435.760 -411.015 ;
        RECT -434.620 -520.175 -434.240 -415.585 ;
        RECT -433.100 -515.605 -432.720 -411.015 ;
        RECT -431.580 -520.175 -431.200 -415.585 ;
        RECT -430.060 -515.605 -429.680 -411.015 ;
        RECT -428.540 -520.175 -428.160 -415.585 ;
        RECT -427.020 -515.605 -426.640 -411.015 ;
        RECT -425.500 -520.175 -425.120 -415.585 ;
        RECT -423.980 -515.605 -423.600 -411.015 ;
        RECT -422.460 -520.175 -422.080 -415.585 ;
        RECT -420.940 -515.605 -420.560 -411.015 ;
        RECT -419.420 -520.175 -419.040 -415.585 ;
        RECT -417.900 -515.605 -417.520 -411.015 ;
        RECT -416.380 -520.175 -416.000 -415.585 ;
        RECT -414.860 -515.605 -414.480 -411.015 ;
        RECT -413.340 -520.175 -412.960 -415.585 ;
        RECT -411.820 -515.605 -411.440 -411.015 ;
        RECT -410.300 -520.175 -409.920 -415.585 ;
        RECT -408.780 -515.605 -408.400 -411.015 ;
        RECT -407.260 -520.175 -406.880 -415.585 ;
        RECT -405.740 -515.605 -405.360 -411.015 ;
        RECT -404.220 -520.175 -403.840 -415.585 ;
        RECT -402.700 -515.605 -402.320 -411.015 ;
        RECT -401.180 -520.175 -400.800 -415.585 ;
        RECT -399.660 -515.605 -399.280 -411.015 ;
        RECT -398.140 -520.175 -397.760 -415.585 ;
        RECT -396.620 -515.605 -396.240 -411.015 ;
        RECT -395.100 -520.175 -394.720 -415.585 ;
        RECT -393.580 -515.605 -393.200 -411.015 ;
        RECT -385.580 -415.595 -385.200 -411.015 ;
        RECT -386.370 -515.605 -385.200 -415.595 ;
        RECT -384.060 -520.175 -383.680 -415.585 ;
        RECT -382.540 -515.605 -382.160 -411.015 ;
        RECT -381.020 -520.175 -380.640 -415.585 ;
        RECT -379.500 -515.605 -379.120 -411.015 ;
        RECT -377.980 -520.175 -377.600 -415.585 ;
        RECT -376.460 -515.605 -376.080 -411.015 ;
        RECT -374.940 -520.175 -374.560 -415.585 ;
        RECT -373.420 -515.605 -373.040 -411.015 ;
        RECT -371.900 -520.175 -371.520 -415.585 ;
        RECT -370.380 -515.605 -370.000 -411.015 ;
        RECT -368.860 -520.175 -368.480 -415.585 ;
        RECT -367.340 -515.605 -366.960 -411.015 ;
        RECT -365.820 -520.175 -365.440 -415.585 ;
        RECT -364.300 -515.605 -363.920 -411.015 ;
        RECT -362.780 -520.175 -362.400 -415.585 ;
        RECT -361.260 -515.605 -360.880 -411.015 ;
        RECT -359.740 -520.175 -359.360 -415.585 ;
        RECT -358.220 -515.605 -357.840 -411.015 ;
        RECT -356.700 -520.175 -356.320 -415.585 ;
        RECT -355.180 -515.605 -354.800 -411.015 ;
        RECT -353.660 -520.175 -353.280 -415.585 ;
        RECT -352.140 -515.605 -351.760 -411.015 ;
        RECT -350.620 -520.175 -350.240 -415.585 ;
        RECT -349.100 -515.605 -348.720 -411.015 ;
        RECT -347.580 -520.175 -347.200 -415.585 ;
        RECT -346.060 -515.605 -345.680 -411.015 ;
        RECT -344.540 -520.175 -344.160 -415.585 ;
        RECT -343.020 -515.605 -342.640 -411.015 ;
        RECT -341.500 -520.175 -341.120 -415.585 ;
        RECT -339.980 -515.605 -339.600 -411.015 ;
        RECT -338.460 -520.175 -338.080 -415.585 ;
        RECT -336.940 -515.605 -336.560 -411.015 ;
        RECT -335.420 -520.175 -335.040 -415.585 ;
        RECT -333.900 -515.605 -333.520 -411.015 ;
        RECT -332.380 -520.175 -332.000 -415.585 ;
        RECT -330.860 -515.605 -330.480 -411.015 ;
        RECT -329.340 -520.175 -328.960 -415.585 ;
        RECT -327.820 -515.605 -327.440 -411.015 ;
        RECT -326.300 -520.175 -325.920 -415.585 ;
        RECT -324.780 -515.605 -324.400 -411.015 ;
        RECT -323.260 -520.175 -322.880 -415.585 ;
        RECT -321.740 -515.605 -321.360 -411.015 ;
        RECT -320.220 -520.175 -319.840 -415.585 ;
        RECT -318.700 -515.605 -318.320 -411.015 ;
        RECT -317.180 -520.175 -316.800 -415.585 ;
        RECT -315.660 -515.605 -315.280 -411.015 ;
        RECT -314.140 -520.175 -313.760 -415.585 ;
        RECT -312.620 -515.605 -312.240 -411.015 ;
        RECT -311.100 -520.175 -310.720 -415.585 ;
        RECT -309.580 -515.605 -309.200 -411.015 ;
        RECT -308.060 -520.175 -307.680 -415.585 ;
        RECT -306.540 -515.605 -306.160 -411.015 ;
        RECT -305.020 -520.175 -304.640 -415.585 ;
        RECT -303.500 -515.605 -303.120 -411.015 ;
        RECT -301.980 -520.175 -301.600 -415.585 ;
        RECT -300.460 -515.605 -300.080 -411.015 ;
        RECT -298.940 -520.175 -298.560 -415.585 ;
        RECT -297.420 -515.605 -297.040 -411.015 ;
        RECT -295.900 -520.175 -295.520 -415.585 ;
        RECT -294.380 -515.605 -294.000 -411.015 ;
        RECT -292.860 -520.175 -292.480 -415.585 ;
        RECT -291.340 -515.605 -290.960 -411.015 ;
        RECT -289.820 -520.175 -289.440 -415.585 ;
        RECT -288.300 -515.605 -287.920 -411.015 ;
        RECT -286.780 -520.175 -286.400 -415.585 ;
        RECT -285.260 -515.605 -284.880 -411.015 ;
        RECT -283.740 -520.175 -283.360 -415.585 ;
        RECT -282.220 -515.605 -281.840 -411.015 ;
        RECT -280.700 -520.175 -280.320 -415.585 ;
        RECT -279.180 -515.605 -278.800 -411.015 ;
        RECT -277.660 -520.175 -277.280 -415.585 ;
        RECT -276.140 -515.605 -275.760 -411.015 ;
        RECT -274.620 -520.175 -274.240 -415.585 ;
        RECT -273.100 -515.605 -272.720 -411.015 ;
        RECT -271.580 -520.175 -271.200 -415.585 ;
        RECT -270.060 -515.605 -269.680 -411.015 ;
        RECT -268.540 -520.175 -268.160 -415.585 ;
        RECT -267.020 -515.605 -266.640 -411.015 ;
        RECT -265.500 -520.175 -265.120 -415.585 ;
        RECT -263.980 -515.605 -263.600 -411.015 ;
        RECT -262.460 -520.175 -262.080 -415.585 ;
        RECT -260.940 -515.605 -260.560 -411.015 ;
        RECT -259.420 -520.175 -259.040 -415.585 ;
        RECT -257.900 -515.605 -257.520 -411.015 ;
        RECT -256.380 -520.175 -256.000 -415.585 ;
        RECT -254.860 -515.605 -254.480 -411.015 ;
        RECT -253.340 -520.175 -252.960 -415.585 ;
        RECT -251.820 -515.605 -251.440 -411.015 ;
        RECT -250.300 -520.175 -249.920 -415.585 ;
        RECT -248.780 -515.605 -248.400 -411.015 ;
        RECT -247.260 -520.175 -246.880 -415.585 ;
        RECT -245.740 -515.605 -245.360 -411.015 ;
        RECT -244.220 -520.175 -243.840 -415.585 ;
        RECT -242.700 -515.605 -242.320 -411.015 ;
        RECT -241.180 -520.175 -240.800 -415.585 ;
        RECT -239.660 -515.605 -239.280 -411.015 ;
        RECT -238.140 -520.175 -237.760 -415.585 ;
        RECT -236.620 -515.605 -236.240 -411.015 ;
        RECT -235.100 -520.175 -234.720 -415.585 ;
        RECT -233.580 -515.605 -233.200 -411.015 ;
        RECT -225.580 -415.595 -225.200 -411.015 ;
        RECT -226.370 -515.605 -225.200 -415.595 ;
        RECT -224.060 -520.175 -223.680 -415.585 ;
        RECT -222.540 -515.605 -222.160 -411.015 ;
        RECT -221.020 -520.175 -220.640 -415.585 ;
        RECT -219.500 -515.605 -219.120 -411.015 ;
        RECT -217.980 -520.175 -217.600 -415.585 ;
        RECT -216.460 -515.605 -216.080 -411.015 ;
        RECT -214.940 -520.175 -214.560 -415.585 ;
        RECT -213.420 -515.605 -213.040 -411.015 ;
        RECT -211.900 -520.175 -211.520 -415.585 ;
        RECT -210.380 -515.605 -210.000 -411.015 ;
        RECT -208.860 -520.175 -208.480 -415.585 ;
        RECT -207.340 -515.605 -206.960 -411.015 ;
        RECT -205.820 -520.175 -205.440 -415.585 ;
        RECT -204.300 -515.605 -203.920 -411.015 ;
        RECT -202.780 -520.175 -202.400 -415.585 ;
        RECT -201.260 -515.605 -200.880 -411.015 ;
        RECT -199.740 -520.175 -199.360 -415.585 ;
        RECT -198.220 -515.605 -197.840 -411.015 ;
        RECT -196.700 -520.175 -196.320 -415.585 ;
        RECT -195.180 -515.605 -194.800 -411.015 ;
        RECT -193.660 -520.175 -193.280 -415.585 ;
        RECT -192.140 -515.605 -191.760 -411.015 ;
        RECT -190.620 -520.175 -190.240 -415.585 ;
        RECT -189.100 -515.605 -188.720 -411.015 ;
        RECT -187.580 -520.175 -187.200 -415.585 ;
        RECT -186.060 -515.605 -185.680 -411.015 ;
        RECT -184.540 -520.175 -184.160 -415.585 ;
        RECT -183.020 -515.605 -182.640 -411.015 ;
        RECT -181.500 -520.175 -181.120 -415.585 ;
        RECT -179.980 -515.605 -179.600 -411.015 ;
        RECT -178.460 -520.175 -178.080 -415.585 ;
        RECT -176.940 -515.605 -176.560 -411.015 ;
        RECT -175.420 -520.175 -175.040 -415.585 ;
        RECT -173.900 -515.605 -173.520 -411.015 ;
        RECT -172.380 -520.175 -172.000 -415.585 ;
        RECT -170.860 -515.605 -170.480 -411.015 ;
        RECT -169.340 -520.175 -168.960 -415.585 ;
        RECT -167.820 -515.605 -167.440 -411.015 ;
        RECT -166.300 -520.175 -165.920 -415.585 ;
        RECT -164.780 -515.605 -164.400 -411.015 ;
        RECT -163.260 -520.175 -162.880 -415.585 ;
        RECT -161.740 -515.605 -161.360 -411.015 ;
        RECT -160.220 -520.175 -159.840 -415.585 ;
        RECT -158.700 -515.605 -158.320 -411.015 ;
        RECT -157.180 -520.175 -156.800 -415.585 ;
        RECT -155.660 -515.605 -155.280 -411.015 ;
        RECT -154.140 -520.175 -153.760 -415.585 ;
        RECT -152.620 -515.605 -152.240 -411.015 ;
        RECT -151.100 -520.175 -150.720 -415.585 ;
        RECT -149.580 -515.605 -149.200 -411.015 ;
        RECT -148.060 -520.175 -147.680 -415.585 ;
        RECT -146.540 -515.605 -146.160 -411.015 ;
        RECT -145.020 -520.175 -144.640 -415.585 ;
        RECT -143.500 -515.605 -143.120 -411.015 ;
        RECT -141.980 -520.175 -141.600 -415.585 ;
        RECT -140.460 -515.605 -140.080 -411.015 ;
        RECT -138.940 -520.175 -138.560 -415.585 ;
        RECT -137.420 -515.605 -137.040 -411.015 ;
        RECT -135.900 -520.175 -135.520 -415.585 ;
        RECT -134.380 -515.605 -134.000 -411.015 ;
        RECT -132.860 -520.175 -132.480 -415.585 ;
        RECT -131.340 -515.605 -130.960 -411.015 ;
        RECT -129.820 -520.175 -129.440 -415.585 ;
        RECT -128.300 -515.605 -127.920 -411.015 ;
        RECT -126.780 -520.175 -126.400 -415.585 ;
        RECT -125.260 -515.605 -124.880 -411.015 ;
        RECT -123.740 -520.175 -123.360 -415.585 ;
        RECT -122.220 -515.605 -121.840 -411.015 ;
        RECT -120.700 -520.175 -120.320 -415.585 ;
        RECT -119.180 -515.605 -118.800 -411.015 ;
        RECT -117.660 -520.175 -117.280 -415.585 ;
        RECT -116.140 -515.605 -115.760 -411.015 ;
        RECT -114.620 -520.175 -114.240 -415.585 ;
        RECT -113.100 -515.605 -112.720 -411.015 ;
        RECT -111.580 -520.175 -111.200 -415.585 ;
        RECT -110.060 -515.605 -109.680 -411.015 ;
        RECT -108.540 -520.175 -108.160 -415.585 ;
        RECT -107.020 -515.605 -106.640 -411.015 ;
        RECT -105.500 -520.175 -105.120 -415.585 ;
        RECT -103.980 -515.605 -103.600 -411.015 ;
        RECT -102.460 -520.175 -102.080 -415.585 ;
        RECT -100.940 -515.605 -100.560 -411.015 ;
        RECT -99.420 -520.175 -99.040 -415.585 ;
        RECT -97.900 -515.605 -97.520 -411.015 ;
        RECT -96.380 -520.175 -96.000 -415.585 ;
        RECT -94.860 -515.605 -94.480 -411.015 ;
        RECT -93.340 -520.175 -92.960 -415.585 ;
        RECT -91.820 -515.605 -91.440 -411.015 ;
        RECT -90.300 -520.175 -89.920 -415.585 ;
        RECT -88.780 -515.605 -88.400 -411.015 ;
        RECT -87.260 -520.175 -86.880 -415.585 ;
        RECT -85.740 -515.605 -85.360 -411.015 ;
        RECT -84.220 -520.175 -83.840 -415.585 ;
        RECT -82.700 -515.605 -82.320 -411.015 ;
        RECT -81.180 -520.175 -80.800 -415.585 ;
        RECT -79.660 -515.605 -79.280 -411.015 ;
        RECT -78.140 -520.175 -77.760 -415.585 ;
        RECT -76.620 -515.605 -76.240 -411.015 ;
        RECT -75.100 -520.175 -74.720 -415.585 ;
        RECT -73.580 -515.605 -73.200 -411.015 ;
        RECT -65.580 -415.595 -65.200 -411.015 ;
        RECT -66.370 -515.605 -65.200 -415.595 ;
        RECT -64.060 -520.175 -63.680 -415.585 ;
        RECT -62.540 -515.605 -62.160 -411.015 ;
        RECT -61.020 -520.175 -60.640 -415.585 ;
        RECT -59.500 -515.605 -59.120 -411.015 ;
        RECT -57.980 -520.175 -57.600 -415.585 ;
        RECT -56.460 -515.605 -56.080 -411.015 ;
        RECT -54.940 -520.175 -54.560 -415.585 ;
        RECT -53.420 -515.605 -53.040 -411.015 ;
        RECT -51.900 -520.175 -51.520 -415.585 ;
        RECT -50.380 -515.605 -50.000 -411.015 ;
        RECT -48.860 -520.175 -48.480 -415.585 ;
        RECT -47.340 -515.605 -46.960 -411.015 ;
        RECT -45.820 -520.175 -45.440 -415.585 ;
        RECT -44.300 -515.605 -43.920 -411.015 ;
        RECT -42.780 -520.175 -42.400 -415.585 ;
        RECT -41.260 -515.605 -40.880 -411.015 ;
        RECT -39.740 -520.175 -39.360 -415.585 ;
        RECT -38.220 -515.605 -37.840 -411.015 ;
        RECT -36.700 -520.175 -36.320 -415.585 ;
        RECT -35.180 -515.605 -34.800 -411.015 ;
        RECT -33.660 -520.175 -33.280 -415.585 ;
        RECT -32.140 -515.605 -31.760 -411.015 ;
        RECT -30.620 -520.175 -30.240 -415.585 ;
        RECT -29.100 -515.605 -28.720 -411.015 ;
        RECT -27.580 -520.175 -27.200 -415.585 ;
        RECT -26.060 -515.605 -25.680 -411.015 ;
        RECT -24.540 -520.175 -24.160 -415.585 ;
        RECT -23.020 -515.605 -22.640 -411.015 ;
        RECT -21.500 -520.175 -21.120 -415.585 ;
        RECT -19.980 -515.605 -19.600 -411.015 ;
        RECT -18.460 -520.175 -18.080 -415.585 ;
        RECT -16.940 -515.605 -16.560 -411.015 ;
        RECT -15.420 -520.175 -15.040 -415.585 ;
        RECT -13.900 -515.605 -13.520 -411.015 ;
        RECT -12.380 -520.175 -12.000 -415.585 ;
        RECT -10.860 -515.605 -10.480 -411.015 ;
        RECT -9.340 -520.175 -8.960 -415.585 ;
        RECT -7.820 -515.605 -7.440 -411.015 ;
        RECT -6.300 -520.175 -5.920 -415.585 ;
        RECT -4.780 -515.605 -4.400 -411.015 ;
        RECT -3.260 -520.175 -2.880 -415.585 ;
        RECT -1.740 -515.605 -1.360 -411.015 ;
        RECT -0.220 -520.175 0.160 -415.585 ;
        RECT 1.300 -515.605 1.680 -411.015 ;
        RECT 2.820 -520.175 3.200 -415.585 ;
        RECT 4.340 -515.605 4.720 -411.015 ;
        RECT 5.860 -520.175 6.240 -415.585 ;
        RECT 7.380 -515.605 7.760 -411.015 ;
        RECT 8.900 -520.175 9.280 -415.585 ;
        RECT 10.420 -515.605 10.800 -411.015 ;
        RECT 11.940 -520.175 12.320 -415.585 ;
        RECT 13.460 -515.605 13.840 -411.015 ;
        RECT 14.980 -520.175 15.360 -415.585 ;
        RECT 16.500 -515.605 16.880 -411.015 ;
        RECT 18.020 -520.175 18.400 -415.585 ;
        RECT 19.540 -515.605 19.920 -411.015 ;
        RECT 21.060 -520.175 21.440 -415.585 ;
        RECT 22.580 -515.605 22.960 -411.015 ;
        RECT 24.100 -520.175 24.480 -415.585 ;
        RECT 25.620 -515.605 26.000 -411.015 ;
        RECT 27.140 -520.175 27.520 -415.585 ;
        RECT 28.660 -515.605 29.040 -411.015 ;
        RECT 30.180 -520.175 30.560 -415.585 ;
        RECT 31.700 -515.605 32.080 -411.015 ;
        RECT 33.220 -520.175 33.600 -415.585 ;
        RECT 34.740 -515.605 35.120 -411.015 ;
        RECT 36.260 -520.175 36.640 -415.585 ;
        RECT 37.780 -515.605 38.160 -411.015 ;
        RECT 39.300 -520.175 39.680 -415.585 ;
        RECT 40.820 -515.605 41.200 -411.015 ;
        RECT 42.340 -520.175 42.720 -415.585 ;
        RECT 43.860 -515.605 44.240 -411.015 ;
        RECT 45.380 -520.175 45.760 -415.585 ;
        RECT 46.900 -515.605 47.280 -411.015 ;
        RECT 48.420 -520.175 48.800 -415.585 ;
        RECT 49.940 -515.605 50.320 -411.015 ;
        RECT 51.460 -520.175 51.840 -415.585 ;
        RECT 52.980 -515.605 53.360 -411.015 ;
        RECT 54.500 -520.175 54.880 -415.585 ;
        RECT 56.020 -515.605 56.400 -411.015 ;
        RECT 57.540 -520.175 57.920 -415.585 ;
        RECT 59.060 -515.605 59.440 -411.015 ;
        RECT 60.580 -520.175 60.960 -415.585 ;
        RECT 62.100 -515.605 62.480 -411.015 ;
        RECT 63.620 -520.175 64.000 -415.585 ;
        RECT 65.140 -515.605 65.520 -411.015 ;
        RECT 66.660 -520.175 67.040 -415.585 ;
        RECT 68.180 -515.605 68.560 -411.015 ;
        RECT 69.700 -520.175 70.080 -415.585 ;
        RECT 71.220 -515.605 71.600 -411.015 ;
        RECT 72.740 -520.175 73.120 -415.585 ;
        RECT 74.260 -515.605 74.640 -411.015 ;
        RECT 75.780 -520.175 76.160 -415.585 ;
        RECT 77.300 -515.605 77.680 -411.015 ;
        RECT 78.820 -520.175 79.200 -415.585 ;
        RECT 80.340 -515.605 80.720 -411.015 ;
        RECT 81.860 -520.175 82.240 -415.585 ;
        RECT 83.380 -515.605 83.760 -411.015 ;
        RECT 84.900 -520.175 85.280 -415.585 ;
        RECT 86.420 -515.605 86.800 -411.015 ;
        RECT 94.420 -415.595 94.800 -411.015 ;
        RECT 93.630 -515.605 94.800 -415.595 ;
        RECT 95.940 -520.175 96.320 -415.585 ;
        RECT 97.460 -515.605 97.840 -411.015 ;
        RECT 98.980 -520.175 99.360 -415.585 ;
        RECT 100.500 -515.605 100.880 -411.015 ;
        RECT 102.020 -520.175 102.400 -415.585 ;
        RECT 103.540 -515.605 103.920 -411.015 ;
        RECT 105.060 -520.175 105.440 -415.585 ;
        RECT 106.580 -515.605 106.960 -411.015 ;
        RECT 108.100 -520.175 108.480 -415.585 ;
        RECT 109.620 -515.605 110.000 -411.015 ;
        RECT 111.140 -520.175 111.520 -415.585 ;
        RECT 112.660 -515.605 113.040 -411.015 ;
        RECT 114.180 -520.175 114.560 -415.585 ;
        RECT 115.700 -515.605 116.080 -411.015 ;
        RECT 117.220 -520.175 117.600 -415.585 ;
        RECT 118.740 -515.605 119.120 -411.015 ;
        RECT 120.260 -520.175 120.640 -415.585 ;
        RECT 121.780 -515.605 122.160 -411.015 ;
        RECT 123.300 -520.175 123.680 -415.585 ;
        RECT 124.820 -515.605 125.200 -411.015 ;
        RECT 126.340 -520.175 126.720 -415.585 ;
        RECT 127.860 -515.605 128.240 -411.015 ;
        RECT 129.380 -520.175 129.760 -415.585 ;
        RECT 130.900 -515.605 131.280 -411.015 ;
        RECT 132.420 -520.175 132.800 -415.585 ;
        RECT 133.940 -515.605 134.320 -411.015 ;
        RECT 135.460 -520.175 135.840 -415.585 ;
        RECT 136.980 -515.605 137.360 -411.015 ;
        RECT 138.500 -520.175 138.880 -415.585 ;
        RECT 140.020 -515.605 140.400 -411.015 ;
        RECT 141.540 -520.175 141.920 -415.585 ;
        RECT 143.060 -515.605 143.440 -411.015 ;
        RECT 144.580 -520.175 144.960 -415.585 ;
        RECT 146.100 -515.605 146.480 -411.015 ;
        RECT 147.620 -520.175 148.000 -415.585 ;
        RECT 149.140 -515.605 149.520 -411.015 ;
        RECT 150.660 -520.175 151.040 -415.585 ;
        RECT 152.180 -515.605 152.560 -411.015 ;
        RECT 153.700 -520.175 154.080 -415.585 ;
        RECT 155.220 -515.605 155.600 -411.015 ;
        RECT 156.740 -520.175 157.120 -415.585 ;
        RECT 158.260 -515.605 158.640 -411.015 ;
        RECT 159.780 -520.175 160.160 -415.585 ;
        RECT 161.300 -515.605 161.680 -411.015 ;
        RECT 162.820 -520.175 163.200 -415.585 ;
        RECT 164.340 -515.605 164.720 -411.015 ;
        RECT 165.860 -520.175 166.240 -415.585 ;
        RECT 167.380 -515.605 167.760 -411.015 ;
        RECT 168.900 -520.175 169.280 -415.585 ;
        RECT 170.420 -515.605 170.800 -411.015 ;
        RECT 171.940 -520.175 172.320 -415.585 ;
        RECT 173.460 -515.605 173.840 -411.015 ;
        RECT 174.980 -520.175 175.360 -415.585 ;
        RECT 176.500 -515.605 176.880 -411.015 ;
        RECT 178.020 -520.175 178.400 -415.585 ;
        RECT 179.540 -515.605 179.920 -411.015 ;
        RECT 181.060 -520.175 181.440 -415.585 ;
        RECT 182.580 -515.605 182.960 -411.015 ;
        RECT 184.100 -520.175 184.480 -415.585 ;
        RECT 185.620 -515.605 186.000 -411.015 ;
        RECT 187.140 -520.175 187.520 -415.585 ;
        RECT 188.660 -515.605 189.040 -411.015 ;
        RECT 190.180 -520.175 190.560 -415.585 ;
        RECT 191.700 -515.605 192.080 -411.015 ;
        RECT 193.220 -520.175 193.600 -415.585 ;
        RECT 194.740 -515.605 195.120 -411.015 ;
        RECT 196.260 -520.175 196.640 -415.585 ;
        RECT 197.780 -515.605 198.160 -411.015 ;
        RECT 199.300 -520.175 199.680 -415.585 ;
        RECT 200.820 -515.605 201.200 -411.015 ;
        RECT 202.340 -520.175 202.720 -415.585 ;
        RECT 203.860 -515.605 204.240 -411.015 ;
        RECT 205.380 -520.175 205.760 -415.585 ;
        RECT 206.900 -515.605 207.280 -411.015 ;
        RECT 208.420 -520.175 208.800 -415.585 ;
        RECT 209.940 -515.605 210.320 -411.015 ;
        RECT 211.460 -520.175 211.840 -415.585 ;
        RECT 212.980 -515.605 213.360 -411.015 ;
        RECT 214.500 -520.175 214.880 -415.585 ;
        RECT 216.020 -515.605 216.400 -411.015 ;
        RECT 217.540 -520.175 217.920 -415.585 ;
        RECT 219.060 -515.605 219.440 -411.015 ;
        RECT 220.580 -520.175 220.960 -415.585 ;
        RECT 222.100 -515.605 222.480 -411.015 ;
        RECT 223.620 -520.175 224.000 -415.585 ;
        RECT 225.140 -515.605 225.520 -411.015 ;
        RECT 226.660 -520.175 227.040 -415.585 ;
        RECT 228.180 -515.605 228.560 -411.015 ;
        RECT 229.700 -520.175 230.080 -415.585 ;
        RECT 231.220 -515.605 231.600 -411.015 ;
        RECT 232.740 -520.175 233.120 -415.585 ;
        RECT 234.260 -515.605 234.640 -411.015 ;
        RECT 235.780 -520.175 236.160 -415.585 ;
        RECT 237.300 -515.605 237.680 -411.015 ;
        RECT 238.820 -520.175 239.200 -415.585 ;
        RECT 240.340 -515.605 240.720 -411.015 ;
        RECT 241.860 -520.175 242.240 -415.585 ;
        RECT 243.380 -515.605 243.760 -411.015 ;
        RECT 244.900 -520.175 245.280 -415.585 ;
        RECT 246.420 -515.605 246.800 -411.015 ;
        RECT 254.420 -415.595 254.800 -411.015 ;
        RECT 253.630 -515.605 254.800 -415.595 ;
        RECT 255.940 -520.175 256.320 -415.585 ;
        RECT 257.460 -515.605 257.840 -411.015 ;
        RECT 258.980 -520.175 259.360 -415.585 ;
        RECT 260.500 -515.605 260.880 -411.015 ;
        RECT 262.020 -520.175 262.400 -415.585 ;
        RECT 263.540 -515.605 263.920 -411.015 ;
        RECT 265.060 -520.175 265.440 -415.585 ;
        RECT 266.580 -515.605 266.960 -411.015 ;
        RECT 268.100 -520.175 268.480 -415.585 ;
        RECT 269.620 -515.605 270.000 -411.015 ;
        RECT 271.140 -520.175 271.520 -415.585 ;
        RECT 272.660 -515.605 273.040 -411.015 ;
        RECT 274.180 -520.175 274.560 -415.585 ;
        RECT 275.700 -515.605 276.080 -411.015 ;
        RECT 277.220 -520.175 277.600 -415.585 ;
        RECT 278.740 -515.605 279.120 -411.015 ;
        RECT 280.260 -520.175 280.640 -415.585 ;
        RECT 281.780 -515.605 282.160 -411.015 ;
        RECT 283.300 -520.175 283.680 -415.585 ;
        RECT 284.820 -515.605 285.200 -411.015 ;
        RECT 286.340 -520.175 286.720 -415.585 ;
        RECT 287.860 -515.605 288.240 -411.015 ;
        RECT 289.380 -520.175 289.760 -415.585 ;
        RECT 290.900 -515.605 291.280 -411.015 ;
        RECT 292.420 -520.175 292.800 -415.585 ;
        RECT 293.940 -515.605 294.320 -411.015 ;
        RECT 295.460 -520.175 295.840 -415.585 ;
        RECT 296.980 -515.605 297.360 -411.015 ;
        RECT 298.500 -520.175 298.880 -415.585 ;
        RECT 300.020 -515.605 300.400 -411.015 ;
        RECT 301.540 -520.175 301.920 -415.585 ;
        RECT 303.060 -515.605 303.440 -411.015 ;
        RECT 304.580 -520.175 304.960 -415.585 ;
        RECT 306.100 -515.605 306.480 -411.015 ;
        RECT 307.620 -520.175 308.000 -415.585 ;
        RECT 309.140 -515.605 309.520 -411.015 ;
        RECT 310.660 -520.175 311.040 -415.585 ;
        RECT 312.180 -515.605 312.560 -411.015 ;
        RECT 313.700 -520.175 314.080 -415.585 ;
        RECT 315.220 -515.605 315.600 -411.015 ;
        RECT 316.740 -520.175 317.120 -415.585 ;
        RECT 318.260 -515.605 318.640 -411.015 ;
        RECT 319.780 -520.175 320.160 -415.585 ;
        RECT 321.300 -515.605 321.680 -411.015 ;
        RECT 322.820 -520.175 323.200 -415.585 ;
        RECT 324.340 -515.605 324.720 -411.015 ;
        RECT 325.860 -520.175 326.240 -415.585 ;
        RECT 327.380 -515.605 327.760 -411.015 ;
        RECT 328.900 -520.175 329.280 -415.585 ;
        RECT 330.420 -515.605 330.800 -411.015 ;
        RECT 331.940 -520.175 332.320 -415.585 ;
        RECT 333.460 -515.605 333.840 -411.015 ;
        RECT 334.980 -520.175 335.360 -415.585 ;
        RECT 336.500 -515.605 336.880 -411.015 ;
        RECT 338.020 -520.175 338.400 -415.585 ;
        RECT 339.540 -515.605 339.920 -411.015 ;
        RECT 341.060 -520.175 341.440 -415.585 ;
        RECT 342.580 -515.605 342.960 -411.015 ;
        RECT 344.100 -520.175 344.480 -415.585 ;
        RECT 345.620 -515.605 346.000 -411.015 ;
        RECT 347.140 -520.175 347.520 -415.585 ;
        RECT 348.660 -515.605 349.040 -411.015 ;
        RECT 350.180 -520.175 350.560 -415.585 ;
        RECT 351.700 -515.605 352.080 -411.015 ;
        RECT 353.220 -520.175 353.600 -415.585 ;
        RECT 354.740 -515.605 355.120 -411.015 ;
        RECT 356.260 -520.175 356.640 -415.585 ;
        RECT 357.780 -515.605 358.160 -411.015 ;
        RECT 359.300 -520.175 359.680 -415.585 ;
        RECT 360.820 -515.605 361.200 -411.015 ;
        RECT 362.340 -520.175 362.720 -415.585 ;
        RECT 363.860 -515.605 364.240 -411.015 ;
        RECT 365.380 -520.175 365.760 -415.585 ;
        RECT 366.900 -515.605 367.280 -411.015 ;
        RECT 368.420 -520.175 368.800 -415.585 ;
        RECT 369.940 -515.605 370.320 -411.015 ;
        RECT 371.460 -520.175 371.840 -415.585 ;
        RECT 372.980 -515.605 373.360 -411.015 ;
        RECT 374.500 -520.175 374.880 -415.585 ;
        RECT 376.020 -515.605 376.400 -411.015 ;
        RECT 377.540 -520.175 377.920 -415.585 ;
        RECT 379.060 -515.605 379.440 -411.015 ;
        RECT 380.580 -520.175 380.960 -415.585 ;
        RECT 382.100 -515.605 382.480 -411.015 ;
        RECT 383.620 -520.175 384.000 -415.585 ;
        RECT 385.140 -515.605 385.520 -411.015 ;
        RECT 386.660 -520.175 387.040 -415.585 ;
        RECT 388.180 -515.605 388.560 -411.015 ;
        RECT 389.700 -520.175 390.080 -415.585 ;
        RECT 391.220 -515.605 391.600 -411.015 ;
        RECT 392.740 -520.175 393.120 -415.585 ;
        RECT 394.260 -515.605 394.640 -411.015 ;
        RECT 395.780 -520.175 396.160 -415.585 ;
        RECT 397.300 -515.605 397.680 -411.015 ;
        RECT 398.820 -520.175 399.200 -415.585 ;
        RECT 400.340 -515.605 400.720 -411.015 ;
        RECT 401.860 -520.175 402.240 -415.585 ;
        RECT 403.380 -515.605 403.760 -411.015 ;
        RECT 404.900 -520.175 405.280 -415.585 ;
        RECT 406.420 -515.605 406.800 -411.015 ;
        RECT 414.420 -415.595 414.800 -411.015 ;
        RECT 413.630 -515.605 414.800 -415.595 ;
        RECT 415.940 -520.175 416.320 -415.585 ;
        RECT 417.460 -515.605 417.840 -411.015 ;
        RECT 418.980 -520.175 419.360 -415.585 ;
        RECT 420.500 -515.605 420.880 -411.015 ;
        RECT 422.020 -520.175 422.400 -415.585 ;
        RECT 423.540 -515.605 423.920 -411.015 ;
        RECT 425.060 -520.175 425.440 -415.585 ;
        RECT 426.580 -515.605 426.960 -411.015 ;
        RECT 428.100 -520.175 428.480 -415.585 ;
        RECT 429.620 -515.605 430.000 -411.015 ;
        RECT 431.140 -520.175 431.520 -415.585 ;
        RECT 432.660 -515.605 433.040 -411.015 ;
        RECT 434.180 -520.175 434.560 -415.585 ;
        RECT 435.700 -515.605 436.080 -411.015 ;
        RECT 437.220 -520.175 437.600 -415.585 ;
        RECT 438.740 -515.605 439.120 -411.015 ;
        RECT 440.260 -520.175 440.640 -415.585 ;
        RECT 441.780 -515.605 442.160 -411.015 ;
        RECT 443.300 -520.175 443.680 -415.585 ;
        RECT 444.820 -515.605 445.200 -411.015 ;
        RECT 446.340 -520.175 446.720 -415.585 ;
        RECT 447.860 -515.605 448.240 -411.015 ;
        RECT 449.380 -520.175 449.760 -415.585 ;
        RECT 450.900 -515.605 451.280 -411.015 ;
        RECT 452.420 -520.175 452.800 -415.585 ;
        RECT 453.940 -515.605 454.320 -411.015 ;
        RECT 455.460 -520.175 455.840 -415.585 ;
        RECT 456.980 -515.605 457.360 -411.015 ;
        RECT 458.500 -520.175 458.880 -415.585 ;
        RECT 460.020 -515.605 460.400 -411.015 ;
        RECT 461.540 -520.175 461.920 -415.585 ;
        RECT 463.060 -515.605 463.440 -411.015 ;
        RECT 464.580 -520.175 464.960 -415.585 ;
        RECT 466.100 -515.605 466.480 -411.015 ;
        RECT 467.620 -520.175 468.000 -415.585 ;
        RECT 469.140 -515.605 469.520 -411.015 ;
        RECT 470.660 -520.175 471.040 -415.585 ;
        RECT 472.180 -515.605 472.560 -411.015 ;
        RECT 473.700 -520.175 474.080 -415.585 ;
        RECT 475.220 -515.605 475.600 -411.015 ;
        RECT 476.740 -520.175 477.120 -415.585 ;
        RECT 478.260 -515.605 478.640 -411.015 ;
        RECT 479.780 -520.175 480.160 -415.585 ;
        RECT 481.300 -515.605 481.680 -411.015 ;
        RECT 482.820 -520.175 483.200 -415.585 ;
        RECT 484.340 -515.605 484.720 -411.015 ;
        RECT 485.860 -520.175 486.240 -415.585 ;
        RECT 487.380 -515.605 487.760 -411.015 ;
        RECT 488.900 -520.175 489.280 -415.585 ;
        RECT 490.420 -515.605 490.800 -411.015 ;
        RECT 491.940 -520.175 492.320 -415.585 ;
        RECT 493.460 -515.605 493.840 -411.015 ;
        RECT 494.980 -520.175 495.360 -415.585 ;
        RECT 496.500 -515.605 496.880 -411.015 ;
        RECT 498.020 -520.175 498.400 -415.585 ;
        RECT 499.540 -515.605 499.920 -411.015 ;
        RECT 501.060 -520.175 501.440 -415.585 ;
        RECT 502.580 -515.605 502.960 -411.015 ;
        RECT 504.100 -520.175 504.480 -415.585 ;
        RECT 505.620 -515.605 506.000 -411.015 ;
        RECT 507.140 -520.175 507.520 -415.585 ;
        RECT 508.660 -515.605 509.040 -411.015 ;
        RECT 510.180 -520.175 510.560 -415.585 ;
        RECT 511.700 -515.605 512.080 -411.015 ;
        RECT 513.220 -520.175 513.600 -415.585 ;
        RECT 514.740 -515.605 515.120 -411.015 ;
        RECT 516.260 -520.175 516.640 -415.585 ;
        RECT 517.780 -515.605 518.160 -411.015 ;
        RECT 519.300 -520.175 519.680 -415.585 ;
        RECT 520.820 -515.605 521.200 -411.015 ;
        RECT 522.340 -520.175 522.720 -415.585 ;
        RECT 523.860 -515.605 524.240 -411.015 ;
        RECT 525.380 -520.175 525.760 -415.585 ;
        RECT 526.900 -515.605 527.280 -411.015 ;
        RECT 528.420 -520.175 528.800 -415.585 ;
        RECT 529.940 -515.605 530.320 -411.015 ;
        RECT 531.460 -520.175 531.840 -415.585 ;
        RECT 532.980 -515.605 533.360 -411.015 ;
        RECT 534.500 -520.175 534.880 -415.585 ;
        RECT 536.020 -515.605 536.400 -411.015 ;
        RECT 537.540 -520.175 537.920 -415.585 ;
        RECT 539.060 -515.605 539.440 -411.015 ;
        RECT 540.580 -520.175 540.960 -415.585 ;
        RECT 542.100 -515.605 542.480 -411.015 ;
        RECT 543.620 -520.175 544.000 -415.585 ;
        RECT 545.140 -515.605 545.520 -411.015 ;
        RECT 546.660 -520.175 547.040 -415.585 ;
        RECT 548.180 -515.605 548.560 -411.015 ;
        RECT 549.700 -520.175 550.080 -415.585 ;
        RECT 551.220 -515.605 551.600 -411.015 ;
        RECT 552.740 -520.175 553.120 -415.585 ;
        RECT 554.260 -515.605 554.640 -411.015 ;
        RECT 555.780 -520.175 556.160 -415.585 ;
        RECT 557.300 -515.605 557.680 -411.015 ;
        RECT 558.820 -520.175 559.200 -415.585 ;
        RECT 560.340 -515.605 560.720 -411.015 ;
        RECT 561.860 -520.175 562.240 -415.585 ;
        RECT 563.380 -515.605 563.760 -411.015 ;
        RECT 564.900 -520.175 565.280 -415.585 ;
        RECT 566.420 -515.605 566.800 -411.015 ;
        RECT 574.420 -415.595 574.800 -411.015 ;
        RECT 573.630 -515.605 574.800 -415.595 ;
        RECT 575.940 -520.175 576.320 -415.585 ;
        RECT 577.460 -515.605 577.840 -411.015 ;
        RECT 578.980 -520.175 579.360 -415.585 ;
        RECT 580.500 -515.605 580.880 -411.015 ;
        RECT 582.020 -520.175 582.400 -415.585 ;
        RECT 583.540 -515.605 583.920 -411.015 ;
        RECT 585.060 -520.175 585.440 -415.585 ;
        RECT 586.580 -515.605 586.960 -411.015 ;
        RECT 588.100 -520.175 588.480 -415.585 ;
        RECT 589.620 -515.605 590.000 -411.015 ;
        RECT 591.140 -520.175 591.520 -415.585 ;
        RECT 592.660 -515.605 593.040 -411.015 ;
        RECT 594.180 -520.175 594.560 -415.585 ;
        RECT 595.700 -515.605 596.080 -411.015 ;
        RECT 597.220 -520.175 597.600 -415.585 ;
        RECT 598.740 -515.605 599.120 -411.015 ;
        RECT 600.260 -520.175 600.640 -415.585 ;
        RECT 601.780 -515.605 602.160 -411.015 ;
        RECT 603.300 -520.175 603.680 -415.585 ;
        RECT 604.820 -515.605 605.200 -411.015 ;
        RECT 606.340 -520.175 606.720 -415.585 ;
        RECT 607.860 -515.605 608.240 -411.015 ;
        RECT 609.380 -520.175 609.760 -415.585 ;
        RECT 610.900 -515.605 611.280 -411.015 ;
        RECT 612.420 -520.175 612.800 -415.585 ;
        RECT 613.940 -515.605 614.320 -411.015 ;
        RECT 615.460 -520.175 615.840 -415.585 ;
        RECT 616.980 -515.605 617.360 -411.015 ;
        RECT 618.500 -520.175 618.880 -415.585 ;
        RECT 620.020 -515.605 620.400 -411.015 ;
        RECT 621.540 -520.175 621.920 -415.585 ;
        RECT 623.060 -515.605 623.440 -411.015 ;
        RECT 624.580 -520.175 624.960 -415.585 ;
        RECT 626.100 -515.605 626.480 -411.015 ;
        RECT 627.620 -520.175 628.000 -415.585 ;
        RECT 629.140 -515.605 629.520 -411.015 ;
        RECT 630.660 -520.175 631.040 -415.585 ;
        RECT 632.180 -515.605 632.560 -411.015 ;
        RECT 633.700 -520.175 634.080 -415.585 ;
        RECT 635.220 -515.605 635.600 -411.015 ;
        RECT 636.740 -520.175 637.120 -415.585 ;
        RECT 638.260 -515.605 638.640 -411.015 ;
        RECT 639.780 -520.175 640.160 -415.585 ;
        RECT 641.300 -515.605 641.680 -411.015 ;
        RECT 642.820 -520.175 643.200 -415.585 ;
        RECT 644.340 -515.605 644.720 -411.015 ;
        RECT 645.860 -520.175 646.240 -415.585 ;
        RECT 647.380 -515.605 647.760 -411.015 ;
        RECT 648.900 -520.175 649.280 -415.585 ;
        RECT 650.420 -515.605 650.800 -411.015 ;
        RECT 651.940 -520.175 652.320 -415.585 ;
        RECT 653.460 -515.605 653.840 -411.015 ;
        RECT 654.980 -520.175 655.360 -415.585 ;
        RECT 656.500 -515.605 656.880 -411.015 ;
        RECT 658.020 -520.175 658.400 -415.585 ;
        RECT 659.540 -515.605 659.920 -411.015 ;
        RECT 661.060 -520.175 661.440 -415.585 ;
        RECT 662.580 -515.605 662.960 -411.015 ;
        RECT 664.100 -520.175 664.480 -415.585 ;
        RECT 665.620 -515.605 666.000 -411.015 ;
        RECT 667.140 -520.175 667.520 -415.585 ;
        RECT 668.660 -515.605 669.040 -411.015 ;
        RECT 670.180 -520.175 670.560 -415.585 ;
        RECT 671.700 -515.605 672.080 -411.015 ;
        RECT 673.220 -520.175 673.600 -415.585 ;
        RECT 674.740 -515.605 675.120 -411.015 ;
        RECT 676.260 -520.175 676.640 -415.585 ;
        RECT 677.780 -515.605 678.160 -411.015 ;
        RECT 679.300 -520.175 679.680 -415.585 ;
        RECT 680.820 -515.605 681.200 -411.015 ;
        RECT 682.340 -520.175 682.720 -415.585 ;
        RECT 683.860 -515.605 684.240 -411.015 ;
        RECT 685.380 -520.175 685.760 -415.585 ;
        RECT 686.900 -515.605 687.280 -411.015 ;
        RECT 688.420 -520.175 688.800 -415.585 ;
        RECT 689.940 -515.605 690.320 -411.015 ;
        RECT 691.460 -520.175 691.840 -415.585 ;
        RECT 692.980 -515.605 693.360 -411.015 ;
        RECT 694.500 -520.175 694.880 -415.585 ;
        RECT 696.020 -515.605 696.400 -411.015 ;
        RECT 697.540 -520.175 697.920 -415.585 ;
        RECT 699.060 -515.605 699.440 -411.015 ;
        RECT 700.580 -520.175 700.960 -415.585 ;
        RECT 702.100 -515.605 702.480 -411.015 ;
        RECT 703.620 -520.175 704.000 -415.585 ;
        RECT 705.140 -515.605 705.520 -411.015 ;
        RECT 706.660 -520.175 707.040 -415.585 ;
        RECT 708.180 -515.605 708.560 -411.015 ;
        RECT 709.700 -520.175 710.080 -415.585 ;
        RECT 711.220 -515.605 711.600 -411.015 ;
        RECT 712.740 -520.175 713.120 -415.585 ;
        RECT 714.260 -515.605 714.640 -411.015 ;
        RECT 715.780 -520.175 716.160 -415.585 ;
        RECT 717.300 -515.605 717.680 -411.015 ;
        RECT 718.820 -520.175 719.200 -415.585 ;
        RECT 720.340 -515.605 720.720 -411.015 ;
        RECT 721.860 -520.175 722.240 -415.585 ;
        RECT 723.380 -515.605 723.760 -411.015 ;
        RECT 724.900 -520.175 725.280 -415.585 ;
        RECT 726.420 -515.605 726.800 -411.015 ;
        RECT 734.420 -415.595 734.800 -411.015 ;
        RECT 733.630 -515.605 734.800 -415.595 ;
        RECT 735.940 -520.175 736.320 -415.585 ;
        RECT 737.460 -515.605 737.840 -411.015 ;
        RECT 738.980 -520.175 739.360 -415.585 ;
        RECT 740.500 -515.605 740.880 -411.015 ;
        RECT 742.020 -520.175 742.400 -415.585 ;
        RECT 743.540 -515.605 743.920 -411.015 ;
        RECT 745.060 -520.175 745.440 -415.585 ;
        RECT 746.580 -515.605 746.960 -411.015 ;
        RECT 748.100 -520.175 748.480 -415.585 ;
        RECT 749.620 -515.605 750.000 -411.015 ;
        RECT 751.140 -520.175 751.520 -415.585 ;
        RECT 752.660 -515.605 753.040 -411.015 ;
        RECT 754.180 -520.175 754.560 -415.585 ;
        RECT 755.700 -515.605 756.080 -411.015 ;
        RECT 757.220 -520.175 757.600 -415.585 ;
        RECT 758.740 -515.605 759.120 -411.015 ;
        RECT 760.260 -520.175 760.640 -415.585 ;
        RECT 761.780 -515.605 762.160 -411.015 ;
        RECT 763.300 -520.175 763.680 -415.585 ;
        RECT 764.820 -515.605 765.200 -411.015 ;
        RECT 766.340 -520.175 766.720 -415.585 ;
        RECT 767.860 -515.605 768.240 -411.015 ;
        RECT 769.380 -520.175 769.760 -415.585 ;
        RECT 770.900 -515.605 771.280 -411.015 ;
        RECT 772.420 -520.175 772.800 -415.585 ;
        RECT 773.940 -515.605 774.320 -411.015 ;
        RECT 775.460 -520.175 775.840 -415.585 ;
        RECT 776.980 -515.605 777.360 -411.015 ;
        RECT 778.500 -520.175 778.880 -415.585 ;
        RECT 780.020 -515.605 780.400 -411.015 ;
        RECT 781.540 -520.175 781.920 -415.585 ;
        RECT 783.060 -515.605 783.440 -411.015 ;
        RECT 784.580 -520.175 784.960 -415.585 ;
        RECT 786.100 -515.605 786.480 -411.015 ;
        RECT 787.620 -520.175 788.000 -415.585 ;
        RECT 789.140 -515.605 789.520 -411.015 ;
        RECT 790.660 -520.175 791.040 -415.585 ;
        RECT 792.180 -515.605 792.560 -411.015 ;
        RECT 793.700 -520.175 794.080 -415.585 ;
        RECT 795.220 -515.605 795.600 -411.015 ;
        RECT 796.740 -520.175 797.120 -415.585 ;
        RECT 798.260 -515.605 798.640 -411.015 ;
        RECT 799.780 -520.175 800.160 -415.585 ;
        RECT 801.300 -515.605 801.680 -411.015 ;
        RECT 802.820 -520.175 803.200 -415.585 ;
        RECT 804.340 -515.605 804.720 -411.015 ;
        RECT 805.860 -520.175 806.240 -415.585 ;
        RECT 807.380 -515.605 807.760 -411.015 ;
        RECT 808.900 -520.175 809.280 -415.585 ;
        RECT 810.420 -515.605 810.800 -411.015 ;
        RECT 811.940 -520.175 812.320 -415.585 ;
        RECT 813.460 -515.605 813.840 -411.015 ;
        RECT 814.980 -520.175 815.360 -415.585 ;
        RECT 816.500 -515.605 816.880 -411.015 ;
        RECT 818.020 -520.175 818.400 -415.585 ;
        RECT 819.540 -515.605 819.920 -411.015 ;
        RECT 821.060 -520.175 821.440 -415.585 ;
        RECT 822.580 -515.605 822.960 -411.015 ;
        RECT 824.100 -520.175 824.480 -415.585 ;
        RECT 825.620 -515.605 826.000 -411.015 ;
        RECT 827.140 -520.175 827.520 -415.585 ;
        RECT 828.660 -515.605 829.040 -411.015 ;
        RECT 830.180 -520.175 830.560 -415.585 ;
        RECT 831.700 -515.605 832.080 -411.015 ;
        RECT 833.220 -520.175 833.600 -415.585 ;
        RECT 834.740 -515.605 835.120 -411.015 ;
        RECT 836.260 -520.175 836.640 -415.585 ;
        RECT 837.780 -515.605 838.160 -411.015 ;
        RECT 839.300 -520.175 839.680 -415.585 ;
        RECT 840.820 -515.605 841.200 -411.015 ;
        RECT 842.340 -520.175 842.720 -415.585 ;
        RECT 843.860 -515.605 844.240 -411.015 ;
        RECT 845.380 -520.175 845.760 -415.585 ;
        RECT 846.900 -515.605 847.280 -411.015 ;
        RECT 848.420 -520.175 848.800 -415.585 ;
        RECT 849.940 -515.605 850.320 -411.015 ;
        RECT 851.460 -520.175 851.840 -415.585 ;
        RECT 852.980 -515.605 853.360 -411.015 ;
        RECT 854.500 -520.175 854.880 -415.585 ;
        RECT 856.020 -515.605 856.400 -411.015 ;
        RECT 857.540 -520.175 857.920 -415.585 ;
        RECT 859.060 -515.605 859.440 -411.015 ;
        RECT 860.580 -520.175 860.960 -415.585 ;
        RECT 862.100 -515.605 862.480 -411.015 ;
        RECT 863.620 -520.175 864.000 -415.585 ;
        RECT 865.140 -515.605 865.520 -411.015 ;
        RECT 866.660 -520.175 867.040 -415.585 ;
        RECT 868.180 -515.605 868.560 -411.015 ;
        RECT 869.700 -520.175 870.080 -415.585 ;
        RECT 871.220 -515.605 871.600 -411.015 ;
        RECT 872.740 -520.175 873.120 -415.585 ;
        RECT 874.260 -515.605 874.640 -411.015 ;
        RECT 875.780 -520.175 876.160 -415.585 ;
        RECT 877.300 -515.605 877.680 -411.015 ;
        RECT 878.820 -520.175 879.200 -415.585 ;
        RECT 880.340 -515.605 880.720 -411.015 ;
        RECT 881.860 -520.175 882.240 -415.585 ;
        RECT 883.380 -515.605 883.760 -411.015 ;
        RECT 884.900 -520.175 885.280 -415.585 ;
        RECT 886.420 -515.605 886.800 -411.015 ;
        RECT 917.630 -490.460 943.025 -477.530 ;
        RECT -544.060 -523.010 891.540 -520.175 ;
        RECT -253.840 -538.180 -210.000 -528.150 ;
        RECT -545.580 -541.015 886.800 -538.180 ;
        RECT -572.210 -645.595 -545.890 -545.595 ;
        RECT -572.210 -856.395 -545.930 -645.595 ;
        RECT -545.580 -645.605 -545.200 -541.015 ;
        RECT -544.060 -650.175 -543.680 -545.585 ;
        RECT -542.540 -645.605 -542.160 -541.015 ;
        RECT -541.020 -650.175 -540.640 -545.585 ;
        RECT -539.500 -645.605 -539.120 -541.015 ;
        RECT -537.980 -650.175 -537.600 -545.585 ;
        RECT -536.460 -645.605 -536.080 -541.015 ;
        RECT -534.940 -650.175 -534.560 -545.585 ;
        RECT -533.420 -645.605 -533.040 -541.015 ;
        RECT -531.900 -650.175 -531.520 -545.585 ;
        RECT -530.380 -645.605 -530.000 -541.015 ;
        RECT -528.860 -650.175 -528.480 -545.585 ;
        RECT -527.340 -645.605 -526.960 -541.015 ;
        RECT -525.820 -650.175 -525.440 -545.585 ;
        RECT -524.300 -645.605 -523.920 -541.015 ;
        RECT -522.780 -650.175 -522.400 -545.585 ;
        RECT -521.260 -645.605 -520.880 -541.015 ;
        RECT -519.740 -650.175 -519.360 -545.585 ;
        RECT -518.220 -645.605 -517.840 -541.015 ;
        RECT -516.700 -650.175 -516.320 -545.585 ;
        RECT -515.180 -645.605 -514.800 -541.015 ;
        RECT -513.660 -650.175 -513.280 -545.585 ;
        RECT -512.140 -645.605 -511.760 -541.015 ;
        RECT -510.620 -650.175 -510.240 -545.585 ;
        RECT -509.100 -645.605 -508.720 -541.015 ;
        RECT -507.580 -650.175 -507.200 -545.585 ;
        RECT -506.060 -645.605 -505.680 -541.015 ;
        RECT -504.540 -650.175 -504.160 -545.585 ;
        RECT -503.020 -645.605 -502.640 -541.015 ;
        RECT -501.500 -650.175 -501.120 -545.585 ;
        RECT -499.980 -645.605 -499.600 -541.015 ;
        RECT -498.460 -650.175 -498.080 -545.585 ;
        RECT -496.940 -645.605 -496.560 -541.015 ;
        RECT -495.420 -650.175 -495.040 -545.585 ;
        RECT -493.900 -645.605 -493.520 -541.015 ;
        RECT -492.380 -650.175 -492.000 -545.585 ;
        RECT -490.860 -645.605 -490.480 -541.015 ;
        RECT -489.340 -650.175 -488.960 -545.585 ;
        RECT -487.820 -645.605 -487.440 -541.015 ;
        RECT -486.300 -650.175 -485.920 -545.585 ;
        RECT -484.780 -645.605 -484.400 -541.015 ;
        RECT -483.260 -650.175 -482.880 -545.585 ;
        RECT -481.740 -645.605 -481.360 -541.015 ;
        RECT -480.220 -650.175 -479.840 -545.585 ;
        RECT -478.700 -645.605 -478.320 -541.015 ;
        RECT -477.180 -650.175 -476.800 -545.585 ;
        RECT -475.660 -645.605 -475.280 -541.015 ;
        RECT -474.140 -650.175 -473.760 -545.585 ;
        RECT -472.620 -645.605 -472.240 -541.015 ;
        RECT -471.100 -650.175 -470.720 -545.585 ;
        RECT -469.580 -645.605 -469.200 -541.015 ;
        RECT -468.060 -650.175 -467.680 -545.585 ;
        RECT -466.540 -645.605 -466.160 -541.015 ;
        RECT -465.020 -650.175 -464.640 -545.585 ;
        RECT -463.500 -645.605 -463.120 -541.015 ;
        RECT -461.980 -650.175 -461.600 -545.585 ;
        RECT -460.460 -645.605 -460.080 -541.015 ;
        RECT -458.940 -650.175 -458.560 -545.585 ;
        RECT -457.420 -645.605 -457.040 -541.015 ;
        RECT -455.900 -650.175 -455.520 -545.585 ;
        RECT -454.380 -645.605 -454.000 -541.015 ;
        RECT -452.860 -650.175 -452.480 -545.585 ;
        RECT -451.340 -645.605 -450.960 -541.015 ;
        RECT -449.820 -650.175 -449.440 -545.585 ;
        RECT -448.300 -645.605 -447.920 -541.015 ;
        RECT -446.780 -650.175 -446.400 -545.585 ;
        RECT -445.260 -645.605 -444.880 -541.015 ;
        RECT -443.740 -650.175 -443.360 -545.585 ;
        RECT -442.220 -645.605 -441.840 -541.015 ;
        RECT -440.700 -650.175 -440.320 -545.585 ;
        RECT -439.180 -645.605 -438.800 -541.015 ;
        RECT -437.660 -650.175 -437.280 -545.585 ;
        RECT -436.140 -645.605 -435.760 -541.015 ;
        RECT -434.620 -650.175 -434.240 -545.585 ;
        RECT -433.100 -645.605 -432.720 -541.015 ;
        RECT -431.580 -650.175 -431.200 -545.585 ;
        RECT -430.060 -645.605 -429.680 -541.015 ;
        RECT -428.540 -650.175 -428.160 -545.585 ;
        RECT -427.020 -645.605 -426.640 -541.015 ;
        RECT -425.500 -650.175 -425.120 -545.585 ;
        RECT -423.980 -645.605 -423.600 -541.015 ;
        RECT -422.460 -650.175 -422.080 -545.585 ;
        RECT -420.940 -645.605 -420.560 -541.015 ;
        RECT -419.420 -650.175 -419.040 -545.585 ;
        RECT -417.900 -645.605 -417.520 -541.015 ;
        RECT -416.380 -650.175 -416.000 -545.585 ;
        RECT -414.860 -645.605 -414.480 -541.015 ;
        RECT -413.340 -650.175 -412.960 -545.585 ;
        RECT -411.820 -645.605 -411.440 -541.015 ;
        RECT -410.300 -650.175 -409.920 -545.585 ;
        RECT -408.780 -645.605 -408.400 -541.015 ;
        RECT -407.260 -650.175 -406.880 -545.585 ;
        RECT -405.740 -645.605 -405.360 -541.015 ;
        RECT -404.220 -650.175 -403.840 -545.585 ;
        RECT -402.700 -645.605 -402.320 -541.015 ;
        RECT -401.180 -650.175 -400.800 -545.585 ;
        RECT -399.660 -645.605 -399.280 -541.015 ;
        RECT -398.140 -650.175 -397.760 -545.585 ;
        RECT -396.620 -645.605 -396.240 -541.015 ;
        RECT -395.100 -650.175 -394.720 -545.585 ;
        RECT -393.580 -645.605 -393.200 -541.015 ;
        RECT -385.580 -545.595 -385.200 -541.015 ;
        RECT -386.370 -645.605 -385.200 -545.595 ;
        RECT -384.060 -650.175 -383.680 -545.585 ;
        RECT -382.540 -645.605 -382.160 -541.015 ;
        RECT -381.020 -650.175 -380.640 -545.585 ;
        RECT -379.500 -645.605 -379.120 -541.015 ;
        RECT -377.980 -650.175 -377.600 -545.585 ;
        RECT -376.460 -645.605 -376.080 -541.015 ;
        RECT -374.940 -650.175 -374.560 -545.585 ;
        RECT -373.420 -645.605 -373.040 -541.015 ;
        RECT -371.900 -650.175 -371.520 -545.585 ;
        RECT -370.380 -645.605 -370.000 -541.015 ;
        RECT -368.860 -650.175 -368.480 -545.585 ;
        RECT -367.340 -645.605 -366.960 -541.015 ;
        RECT -365.820 -650.175 -365.440 -545.585 ;
        RECT -364.300 -645.605 -363.920 -541.015 ;
        RECT -362.780 -650.175 -362.400 -545.585 ;
        RECT -361.260 -645.605 -360.880 -541.015 ;
        RECT -359.740 -650.175 -359.360 -545.585 ;
        RECT -358.220 -645.605 -357.840 -541.015 ;
        RECT -356.700 -650.175 -356.320 -545.585 ;
        RECT -355.180 -645.605 -354.800 -541.015 ;
        RECT -353.660 -650.175 -353.280 -545.585 ;
        RECT -352.140 -645.605 -351.760 -541.015 ;
        RECT -350.620 -650.175 -350.240 -545.585 ;
        RECT -349.100 -645.605 -348.720 -541.015 ;
        RECT -347.580 -650.175 -347.200 -545.585 ;
        RECT -346.060 -645.605 -345.680 -541.015 ;
        RECT -344.540 -650.175 -344.160 -545.585 ;
        RECT -343.020 -645.605 -342.640 -541.015 ;
        RECT -341.500 -650.175 -341.120 -545.585 ;
        RECT -339.980 -645.605 -339.600 -541.015 ;
        RECT -338.460 -650.175 -338.080 -545.585 ;
        RECT -336.940 -645.605 -336.560 -541.015 ;
        RECT -335.420 -650.175 -335.040 -545.585 ;
        RECT -333.900 -645.605 -333.520 -541.015 ;
        RECT -332.380 -650.175 -332.000 -545.585 ;
        RECT -330.860 -645.605 -330.480 -541.015 ;
        RECT -329.340 -650.175 -328.960 -545.585 ;
        RECT -327.820 -645.605 -327.440 -541.015 ;
        RECT -326.300 -650.175 -325.920 -545.585 ;
        RECT -324.780 -645.605 -324.400 -541.015 ;
        RECT -323.260 -650.175 -322.880 -545.585 ;
        RECT -321.740 -645.605 -321.360 -541.015 ;
        RECT -320.220 -650.175 -319.840 -545.585 ;
        RECT -318.700 -645.605 -318.320 -541.015 ;
        RECT -317.180 -650.175 -316.800 -545.585 ;
        RECT -315.660 -645.605 -315.280 -541.015 ;
        RECT -314.140 -650.175 -313.760 -545.585 ;
        RECT -312.620 -645.605 -312.240 -541.015 ;
        RECT -311.100 -650.175 -310.720 -545.585 ;
        RECT -309.580 -645.605 -309.200 -541.015 ;
        RECT -308.060 -650.175 -307.680 -545.585 ;
        RECT -306.540 -645.605 -306.160 -541.015 ;
        RECT -305.020 -650.175 -304.640 -545.585 ;
        RECT -303.500 -645.605 -303.120 -541.015 ;
        RECT -301.980 -650.175 -301.600 -545.585 ;
        RECT -300.460 -645.605 -300.080 -541.015 ;
        RECT -298.940 -650.175 -298.560 -545.585 ;
        RECT -297.420 -645.605 -297.040 -541.015 ;
        RECT -295.900 -650.175 -295.520 -545.585 ;
        RECT -294.380 -645.605 -294.000 -541.015 ;
        RECT -292.860 -650.175 -292.480 -545.585 ;
        RECT -291.340 -645.605 -290.960 -541.015 ;
        RECT -289.820 -650.175 -289.440 -545.585 ;
        RECT -288.300 -645.605 -287.920 -541.015 ;
        RECT -286.780 -650.175 -286.400 -545.585 ;
        RECT -285.260 -645.605 -284.880 -541.015 ;
        RECT -283.740 -650.175 -283.360 -545.585 ;
        RECT -282.220 -645.605 -281.840 -541.015 ;
        RECT -280.700 -650.175 -280.320 -545.585 ;
        RECT -279.180 -645.605 -278.800 -541.015 ;
        RECT -277.660 -650.175 -277.280 -545.585 ;
        RECT -276.140 -645.605 -275.760 -541.015 ;
        RECT -274.620 -650.175 -274.240 -545.585 ;
        RECT -273.100 -645.605 -272.720 -541.015 ;
        RECT -271.580 -650.175 -271.200 -545.585 ;
        RECT -270.060 -645.605 -269.680 -541.015 ;
        RECT -268.540 -650.175 -268.160 -545.585 ;
        RECT -267.020 -645.605 -266.640 -541.015 ;
        RECT -265.500 -650.175 -265.120 -545.585 ;
        RECT -263.980 -645.605 -263.600 -541.015 ;
        RECT -262.460 -650.175 -262.080 -545.585 ;
        RECT -260.940 -645.605 -260.560 -541.015 ;
        RECT -259.420 -650.175 -259.040 -545.585 ;
        RECT -257.900 -645.605 -257.520 -541.015 ;
        RECT -256.380 -650.175 -256.000 -545.585 ;
        RECT -254.860 -645.605 -254.480 -541.015 ;
        RECT -253.340 -650.175 -252.960 -545.585 ;
        RECT -251.820 -645.605 -251.440 -541.015 ;
        RECT -250.300 -650.175 -249.920 -545.585 ;
        RECT -248.780 -645.605 -248.400 -541.015 ;
        RECT -247.260 -650.175 -246.880 -545.585 ;
        RECT -245.740 -645.605 -245.360 -541.015 ;
        RECT -244.220 -650.175 -243.840 -545.585 ;
        RECT -242.700 -645.605 -242.320 -541.015 ;
        RECT -241.180 -650.175 -240.800 -545.585 ;
        RECT -239.660 -645.605 -239.280 -541.015 ;
        RECT -238.140 -650.175 -237.760 -545.585 ;
        RECT -236.620 -645.605 -236.240 -541.015 ;
        RECT -235.100 -650.175 -234.720 -545.585 ;
        RECT -233.580 -645.605 -233.200 -541.015 ;
        RECT -225.580 -545.595 -225.200 -541.015 ;
        RECT -226.370 -645.605 -225.200 -545.595 ;
        RECT -224.060 -650.175 -223.680 -545.585 ;
        RECT -222.540 -645.605 -222.160 -541.015 ;
        RECT -221.020 -650.175 -220.640 -545.585 ;
        RECT -219.500 -645.605 -219.120 -541.015 ;
        RECT -217.980 -650.175 -217.600 -545.585 ;
        RECT -216.460 -645.605 -216.080 -541.015 ;
        RECT -214.940 -650.175 -214.560 -545.585 ;
        RECT -213.420 -645.605 -213.040 -541.015 ;
        RECT -211.900 -650.175 -211.520 -545.585 ;
        RECT -210.380 -645.605 -210.000 -541.015 ;
        RECT -208.860 -650.175 -208.480 -545.585 ;
        RECT -207.340 -645.605 -206.960 -541.015 ;
        RECT -205.820 -650.175 -205.440 -545.585 ;
        RECT -204.300 -645.605 -203.920 -541.015 ;
        RECT -202.780 -650.175 -202.400 -545.585 ;
        RECT -201.260 -645.605 -200.880 -541.015 ;
        RECT -199.740 -650.175 -199.360 -545.585 ;
        RECT -198.220 -645.605 -197.840 -541.015 ;
        RECT -196.700 -650.175 -196.320 -545.585 ;
        RECT -195.180 -645.605 -194.800 -541.015 ;
        RECT -193.660 -650.175 -193.280 -545.585 ;
        RECT -192.140 -645.605 -191.760 -541.015 ;
        RECT -190.620 -650.175 -190.240 -545.585 ;
        RECT -189.100 -645.605 -188.720 -541.015 ;
        RECT -187.580 -650.175 -187.200 -545.585 ;
        RECT -186.060 -645.605 -185.680 -541.015 ;
        RECT -184.540 -650.175 -184.160 -545.585 ;
        RECT -183.020 -645.605 -182.640 -541.015 ;
        RECT -181.500 -650.175 -181.120 -545.585 ;
        RECT -179.980 -645.605 -179.600 -541.015 ;
        RECT -178.460 -650.175 -178.080 -545.585 ;
        RECT -176.940 -645.605 -176.560 -541.015 ;
        RECT -175.420 -650.175 -175.040 -545.585 ;
        RECT -173.900 -645.605 -173.520 -541.015 ;
        RECT -172.380 -650.175 -172.000 -545.585 ;
        RECT -170.860 -645.605 -170.480 -541.015 ;
        RECT -169.340 -650.175 -168.960 -545.585 ;
        RECT -167.820 -645.605 -167.440 -541.015 ;
        RECT -166.300 -650.175 -165.920 -545.585 ;
        RECT -164.780 -645.605 -164.400 -541.015 ;
        RECT -163.260 -650.175 -162.880 -545.585 ;
        RECT -161.740 -645.605 -161.360 -541.015 ;
        RECT -160.220 -650.175 -159.840 -545.585 ;
        RECT -158.700 -645.605 -158.320 -541.015 ;
        RECT -157.180 -650.175 -156.800 -545.585 ;
        RECT -155.660 -645.605 -155.280 -541.015 ;
        RECT -154.140 -650.175 -153.760 -545.585 ;
        RECT -152.620 -645.605 -152.240 -541.015 ;
        RECT -151.100 -650.175 -150.720 -545.585 ;
        RECT -149.580 -645.605 -149.200 -541.015 ;
        RECT -148.060 -650.175 -147.680 -545.585 ;
        RECT -146.540 -645.605 -146.160 -541.015 ;
        RECT -145.020 -650.175 -144.640 -545.585 ;
        RECT -143.500 -645.605 -143.120 -541.015 ;
        RECT -141.980 -650.175 -141.600 -545.585 ;
        RECT -140.460 -645.605 -140.080 -541.015 ;
        RECT -138.940 -650.175 -138.560 -545.585 ;
        RECT -137.420 -645.605 -137.040 -541.015 ;
        RECT -135.900 -650.175 -135.520 -545.585 ;
        RECT -134.380 -645.605 -134.000 -541.015 ;
        RECT -132.860 -650.175 -132.480 -545.585 ;
        RECT -131.340 -645.605 -130.960 -541.015 ;
        RECT -129.820 -650.175 -129.440 -545.585 ;
        RECT -128.300 -645.605 -127.920 -541.015 ;
        RECT -126.780 -650.175 -126.400 -545.585 ;
        RECT -125.260 -645.605 -124.880 -541.015 ;
        RECT -123.740 -650.175 -123.360 -545.585 ;
        RECT -122.220 -645.605 -121.840 -541.015 ;
        RECT -120.700 -650.175 -120.320 -545.585 ;
        RECT -119.180 -645.605 -118.800 -541.015 ;
        RECT -117.660 -650.175 -117.280 -545.585 ;
        RECT -116.140 -645.605 -115.760 -541.015 ;
        RECT -114.620 -650.175 -114.240 -545.585 ;
        RECT -113.100 -645.605 -112.720 -541.015 ;
        RECT -111.580 -650.175 -111.200 -545.585 ;
        RECT -110.060 -645.605 -109.680 -541.015 ;
        RECT -108.540 -650.175 -108.160 -545.585 ;
        RECT -107.020 -645.605 -106.640 -541.015 ;
        RECT -105.500 -650.175 -105.120 -545.585 ;
        RECT -103.980 -645.605 -103.600 -541.015 ;
        RECT -102.460 -650.175 -102.080 -545.585 ;
        RECT -100.940 -645.605 -100.560 -541.015 ;
        RECT -99.420 -650.175 -99.040 -545.585 ;
        RECT -97.900 -645.605 -97.520 -541.015 ;
        RECT -96.380 -650.175 -96.000 -545.585 ;
        RECT -94.860 -645.605 -94.480 -541.015 ;
        RECT -93.340 -650.175 -92.960 -545.585 ;
        RECT -91.820 -645.605 -91.440 -541.015 ;
        RECT -90.300 -650.175 -89.920 -545.585 ;
        RECT -88.780 -645.605 -88.400 -541.015 ;
        RECT -87.260 -650.175 -86.880 -545.585 ;
        RECT -85.740 -645.605 -85.360 -541.015 ;
        RECT -84.220 -650.175 -83.840 -545.585 ;
        RECT -82.700 -645.605 -82.320 -541.015 ;
        RECT -81.180 -650.175 -80.800 -545.585 ;
        RECT -79.660 -645.605 -79.280 -541.015 ;
        RECT -78.140 -650.175 -77.760 -545.585 ;
        RECT -76.620 -645.605 -76.240 -541.015 ;
        RECT -75.100 -650.175 -74.720 -545.585 ;
        RECT -73.580 -645.605 -73.200 -541.015 ;
        RECT -65.580 -545.595 -65.200 -541.015 ;
        RECT -66.370 -645.605 -65.200 -545.595 ;
        RECT -64.060 -650.175 -63.680 -545.585 ;
        RECT -62.540 -645.605 -62.160 -541.015 ;
        RECT -61.020 -650.175 -60.640 -545.585 ;
        RECT -59.500 -645.605 -59.120 -541.015 ;
        RECT -57.980 -650.175 -57.600 -545.585 ;
        RECT -56.460 -645.605 -56.080 -541.015 ;
        RECT -54.940 -650.175 -54.560 -545.585 ;
        RECT -53.420 -645.605 -53.040 -541.015 ;
        RECT -51.900 -650.175 -51.520 -545.585 ;
        RECT -50.380 -645.605 -50.000 -541.015 ;
        RECT -48.860 -650.175 -48.480 -545.585 ;
        RECT -47.340 -645.605 -46.960 -541.015 ;
        RECT -45.820 -650.175 -45.440 -545.585 ;
        RECT -44.300 -645.605 -43.920 -541.015 ;
        RECT -42.780 -650.175 -42.400 -545.585 ;
        RECT -41.260 -645.605 -40.880 -541.015 ;
        RECT -39.740 -650.175 -39.360 -545.585 ;
        RECT -38.220 -645.605 -37.840 -541.015 ;
        RECT -36.700 -650.175 -36.320 -545.585 ;
        RECT -35.180 -645.605 -34.800 -541.015 ;
        RECT -33.660 -650.175 -33.280 -545.585 ;
        RECT -32.140 -645.605 -31.760 -541.015 ;
        RECT -30.620 -650.175 -30.240 -545.585 ;
        RECT -29.100 -645.605 -28.720 -541.015 ;
        RECT -27.580 -650.175 -27.200 -545.585 ;
        RECT -26.060 -645.605 -25.680 -541.015 ;
        RECT -24.540 -650.175 -24.160 -545.585 ;
        RECT -23.020 -645.605 -22.640 -541.015 ;
        RECT -21.500 -650.175 -21.120 -545.585 ;
        RECT -19.980 -645.605 -19.600 -541.015 ;
        RECT -18.460 -650.175 -18.080 -545.585 ;
        RECT -16.940 -645.605 -16.560 -541.015 ;
        RECT -15.420 -650.175 -15.040 -545.585 ;
        RECT -13.900 -645.605 -13.520 -541.015 ;
        RECT -12.380 -650.175 -12.000 -545.585 ;
        RECT -10.860 -645.605 -10.480 -541.015 ;
        RECT -9.340 -650.175 -8.960 -545.585 ;
        RECT -7.820 -645.605 -7.440 -541.015 ;
        RECT -6.300 -650.175 -5.920 -545.585 ;
        RECT -4.780 -645.605 -4.400 -541.015 ;
        RECT -3.260 -650.175 -2.880 -545.585 ;
        RECT -1.740 -645.605 -1.360 -541.015 ;
        RECT -0.220 -650.175 0.160 -545.585 ;
        RECT 1.300 -645.605 1.680 -541.015 ;
        RECT 2.820 -650.175 3.200 -545.585 ;
        RECT 4.340 -645.605 4.720 -541.015 ;
        RECT 5.860 -650.175 6.240 -545.585 ;
        RECT 7.380 -645.605 7.760 -541.015 ;
        RECT 8.900 -650.175 9.280 -545.585 ;
        RECT 10.420 -645.605 10.800 -541.015 ;
        RECT 11.940 -650.175 12.320 -545.585 ;
        RECT 13.460 -645.605 13.840 -541.015 ;
        RECT 14.980 -650.175 15.360 -545.585 ;
        RECT 16.500 -645.605 16.880 -541.015 ;
        RECT 18.020 -650.175 18.400 -545.585 ;
        RECT 19.540 -645.605 19.920 -541.015 ;
        RECT 21.060 -650.175 21.440 -545.585 ;
        RECT 22.580 -645.605 22.960 -541.015 ;
        RECT 24.100 -650.175 24.480 -545.585 ;
        RECT 25.620 -645.605 26.000 -541.015 ;
        RECT 27.140 -650.175 27.520 -545.585 ;
        RECT 28.660 -645.605 29.040 -541.015 ;
        RECT 30.180 -650.175 30.560 -545.585 ;
        RECT 31.700 -645.605 32.080 -541.015 ;
        RECT 33.220 -650.175 33.600 -545.585 ;
        RECT 34.740 -645.605 35.120 -541.015 ;
        RECT 36.260 -650.175 36.640 -545.585 ;
        RECT 37.780 -645.605 38.160 -541.015 ;
        RECT 39.300 -650.175 39.680 -545.585 ;
        RECT 40.820 -645.605 41.200 -541.015 ;
        RECT 42.340 -650.175 42.720 -545.585 ;
        RECT 43.860 -645.605 44.240 -541.015 ;
        RECT 45.380 -650.175 45.760 -545.585 ;
        RECT 46.900 -645.605 47.280 -541.015 ;
        RECT 48.420 -650.175 48.800 -545.585 ;
        RECT 49.940 -645.605 50.320 -541.015 ;
        RECT 51.460 -650.175 51.840 -545.585 ;
        RECT 52.980 -645.605 53.360 -541.015 ;
        RECT 54.500 -650.175 54.880 -545.585 ;
        RECT 56.020 -645.605 56.400 -541.015 ;
        RECT 57.540 -650.175 57.920 -545.585 ;
        RECT 59.060 -645.605 59.440 -541.015 ;
        RECT 60.580 -650.175 60.960 -545.585 ;
        RECT 62.100 -645.605 62.480 -541.015 ;
        RECT 63.620 -650.175 64.000 -545.585 ;
        RECT 65.140 -645.605 65.520 -541.015 ;
        RECT 66.660 -650.175 67.040 -545.585 ;
        RECT 68.180 -645.605 68.560 -541.015 ;
        RECT 69.700 -650.175 70.080 -545.585 ;
        RECT 71.220 -645.605 71.600 -541.015 ;
        RECT 72.740 -650.175 73.120 -545.585 ;
        RECT 74.260 -645.605 74.640 -541.015 ;
        RECT 75.780 -650.175 76.160 -545.585 ;
        RECT 77.300 -645.605 77.680 -541.015 ;
        RECT 78.820 -650.175 79.200 -545.585 ;
        RECT 80.340 -645.605 80.720 -541.015 ;
        RECT 81.860 -650.175 82.240 -545.585 ;
        RECT 83.380 -645.605 83.760 -541.015 ;
        RECT 84.900 -650.175 85.280 -545.585 ;
        RECT 86.420 -645.605 86.800 -541.015 ;
        RECT 94.420 -545.595 94.800 -541.015 ;
        RECT 93.630 -645.605 94.800 -545.595 ;
        RECT 95.940 -650.175 96.320 -545.585 ;
        RECT 97.460 -645.605 97.840 -541.015 ;
        RECT 98.980 -650.175 99.360 -545.585 ;
        RECT 100.500 -645.605 100.880 -541.015 ;
        RECT 102.020 -650.175 102.400 -545.585 ;
        RECT 103.540 -645.605 103.920 -541.015 ;
        RECT 105.060 -650.175 105.440 -545.585 ;
        RECT 106.580 -645.605 106.960 -541.015 ;
        RECT 108.100 -650.175 108.480 -545.585 ;
        RECT 109.620 -645.605 110.000 -541.015 ;
        RECT 111.140 -650.175 111.520 -545.585 ;
        RECT 112.660 -645.605 113.040 -541.015 ;
        RECT 114.180 -650.175 114.560 -545.585 ;
        RECT 115.700 -645.605 116.080 -541.015 ;
        RECT 117.220 -650.175 117.600 -545.585 ;
        RECT 118.740 -645.605 119.120 -541.015 ;
        RECT 120.260 -650.175 120.640 -545.585 ;
        RECT 121.780 -645.605 122.160 -541.015 ;
        RECT 123.300 -650.175 123.680 -545.585 ;
        RECT 124.820 -645.605 125.200 -541.015 ;
        RECT 126.340 -650.175 126.720 -545.585 ;
        RECT 127.860 -645.605 128.240 -541.015 ;
        RECT 129.380 -650.175 129.760 -545.585 ;
        RECT 130.900 -645.605 131.280 -541.015 ;
        RECT 132.420 -650.175 132.800 -545.585 ;
        RECT 133.940 -645.605 134.320 -541.015 ;
        RECT 135.460 -650.175 135.840 -545.585 ;
        RECT 136.980 -645.605 137.360 -541.015 ;
        RECT 138.500 -650.175 138.880 -545.585 ;
        RECT 140.020 -645.605 140.400 -541.015 ;
        RECT 141.540 -650.175 141.920 -545.585 ;
        RECT 143.060 -645.605 143.440 -541.015 ;
        RECT 144.580 -650.175 144.960 -545.585 ;
        RECT 146.100 -645.605 146.480 -541.015 ;
        RECT 147.620 -650.175 148.000 -545.585 ;
        RECT 149.140 -645.605 149.520 -541.015 ;
        RECT 150.660 -650.175 151.040 -545.585 ;
        RECT 152.180 -645.605 152.560 -541.015 ;
        RECT 153.700 -650.175 154.080 -545.585 ;
        RECT 155.220 -645.605 155.600 -541.015 ;
        RECT 156.740 -650.175 157.120 -545.585 ;
        RECT 158.260 -645.605 158.640 -541.015 ;
        RECT 159.780 -650.175 160.160 -545.585 ;
        RECT 161.300 -645.605 161.680 -541.015 ;
        RECT 162.820 -650.175 163.200 -545.585 ;
        RECT 164.340 -645.605 164.720 -541.015 ;
        RECT 165.860 -650.175 166.240 -545.585 ;
        RECT 167.380 -645.605 167.760 -541.015 ;
        RECT 168.900 -650.175 169.280 -545.585 ;
        RECT 170.420 -645.605 170.800 -541.015 ;
        RECT 171.940 -650.175 172.320 -545.585 ;
        RECT 173.460 -645.605 173.840 -541.015 ;
        RECT 174.980 -650.175 175.360 -545.585 ;
        RECT 176.500 -645.605 176.880 -541.015 ;
        RECT 178.020 -650.175 178.400 -545.585 ;
        RECT 179.540 -645.605 179.920 -541.015 ;
        RECT 181.060 -650.175 181.440 -545.585 ;
        RECT 182.580 -645.605 182.960 -541.015 ;
        RECT 184.100 -650.175 184.480 -545.585 ;
        RECT 185.620 -645.605 186.000 -541.015 ;
        RECT 187.140 -650.175 187.520 -545.585 ;
        RECT 188.660 -645.605 189.040 -541.015 ;
        RECT 190.180 -650.175 190.560 -545.585 ;
        RECT 191.700 -645.605 192.080 -541.015 ;
        RECT 193.220 -650.175 193.600 -545.585 ;
        RECT 194.740 -645.605 195.120 -541.015 ;
        RECT 196.260 -650.175 196.640 -545.585 ;
        RECT 197.780 -645.605 198.160 -541.015 ;
        RECT 199.300 -650.175 199.680 -545.585 ;
        RECT 200.820 -645.605 201.200 -541.015 ;
        RECT 202.340 -650.175 202.720 -545.585 ;
        RECT 203.860 -645.605 204.240 -541.015 ;
        RECT 205.380 -650.175 205.760 -545.585 ;
        RECT 206.900 -645.605 207.280 -541.015 ;
        RECT 208.420 -650.175 208.800 -545.585 ;
        RECT 209.940 -645.605 210.320 -541.015 ;
        RECT 211.460 -650.175 211.840 -545.585 ;
        RECT 212.980 -645.605 213.360 -541.015 ;
        RECT 214.500 -650.175 214.880 -545.585 ;
        RECT 216.020 -645.605 216.400 -541.015 ;
        RECT 217.540 -650.175 217.920 -545.585 ;
        RECT 219.060 -645.605 219.440 -541.015 ;
        RECT 220.580 -650.175 220.960 -545.585 ;
        RECT 222.100 -645.605 222.480 -541.015 ;
        RECT 223.620 -650.175 224.000 -545.585 ;
        RECT 225.140 -645.605 225.520 -541.015 ;
        RECT 226.660 -650.175 227.040 -545.585 ;
        RECT 228.180 -645.605 228.560 -541.015 ;
        RECT 229.700 -650.175 230.080 -545.585 ;
        RECT 231.220 -645.605 231.600 -541.015 ;
        RECT 232.740 -650.175 233.120 -545.585 ;
        RECT 234.260 -645.605 234.640 -541.015 ;
        RECT 235.780 -650.175 236.160 -545.585 ;
        RECT 237.300 -645.605 237.680 -541.015 ;
        RECT 238.820 -650.175 239.200 -545.585 ;
        RECT 240.340 -645.605 240.720 -541.015 ;
        RECT 241.860 -650.175 242.240 -545.585 ;
        RECT 243.380 -645.605 243.760 -541.015 ;
        RECT 244.900 -650.175 245.280 -545.585 ;
        RECT 246.420 -645.605 246.800 -541.015 ;
        RECT 254.420 -545.595 254.800 -541.015 ;
        RECT 253.630 -645.605 254.800 -545.595 ;
        RECT 255.940 -650.175 256.320 -545.585 ;
        RECT 257.460 -645.605 257.840 -541.015 ;
        RECT 258.980 -650.175 259.360 -545.585 ;
        RECT 260.500 -645.605 260.880 -541.015 ;
        RECT 262.020 -650.175 262.400 -545.585 ;
        RECT 263.540 -645.605 263.920 -541.015 ;
        RECT 265.060 -650.175 265.440 -545.585 ;
        RECT 266.580 -645.605 266.960 -541.015 ;
        RECT 268.100 -650.175 268.480 -545.585 ;
        RECT 269.620 -645.605 270.000 -541.015 ;
        RECT 271.140 -650.175 271.520 -545.585 ;
        RECT 272.660 -645.605 273.040 -541.015 ;
        RECT 274.180 -650.175 274.560 -545.585 ;
        RECT 275.700 -645.605 276.080 -541.015 ;
        RECT 277.220 -650.175 277.600 -545.585 ;
        RECT 278.740 -645.605 279.120 -541.015 ;
        RECT 280.260 -650.175 280.640 -545.585 ;
        RECT 281.780 -645.605 282.160 -541.015 ;
        RECT 283.300 -650.175 283.680 -545.585 ;
        RECT 284.820 -645.605 285.200 -541.015 ;
        RECT 286.340 -650.175 286.720 -545.585 ;
        RECT 287.860 -645.605 288.240 -541.015 ;
        RECT 289.380 -650.175 289.760 -545.585 ;
        RECT 290.900 -645.605 291.280 -541.015 ;
        RECT 292.420 -650.175 292.800 -545.585 ;
        RECT 293.940 -645.605 294.320 -541.015 ;
        RECT 295.460 -650.175 295.840 -545.585 ;
        RECT 296.980 -645.605 297.360 -541.015 ;
        RECT 298.500 -650.175 298.880 -545.585 ;
        RECT 300.020 -645.605 300.400 -541.015 ;
        RECT 301.540 -650.175 301.920 -545.585 ;
        RECT 303.060 -645.605 303.440 -541.015 ;
        RECT 304.580 -650.175 304.960 -545.585 ;
        RECT 306.100 -645.605 306.480 -541.015 ;
        RECT 307.620 -650.175 308.000 -545.585 ;
        RECT 309.140 -645.605 309.520 -541.015 ;
        RECT 310.660 -650.175 311.040 -545.585 ;
        RECT 312.180 -645.605 312.560 -541.015 ;
        RECT 313.700 -650.175 314.080 -545.585 ;
        RECT 315.220 -645.605 315.600 -541.015 ;
        RECT 316.740 -650.175 317.120 -545.585 ;
        RECT 318.260 -645.605 318.640 -541.015 ;
        RECT 319.780 -650.175 320.160 -545.585 ;
        RECT 321.300 -645.605 321.680 -541.015 ;
        RECT 322.820 -650.175 323.200 -545.585 ;
        RECT 324.340 -645.605 324.720 -541.015 ;
        RECT 325.860 -650.175 326.240 -545.585 ;
        RECT 327.380 -645.605 327.760 -541.015 ;
        RECT 328.900 -650.175 329.280 -545.585 ;
        RECT 330.420 -645.605 330.800 -541.015 ;
        RECT 331.940 -650.175 332.320 -545.585 ;
        RECT 333.460 -645.605 333.840 -541.015 ;
        RECT 334.980 -650.175 335.360 -545.585 ;
        RECT 336.500 -645.605 336.880 -541.015 ;
        RECT 338.020 -650.175 338.400 -545.585 ;
        RECT 339.540 -645.605 339.920 -541.015 ;
        RECT 341.060 -650.175 341.440 -545.585 ;
        RECT 342.580 -645.605 342.960 -541.015 ;
        RECT 344.100 -650.175 344.480 -545.585 ;
        RECT 345.620 -645.605 346.000 -541.015 ;
        RECT 347.140 -650.175 347.520 -545.585 ;
        RECT 348.660 -645.605 349.040 -541.015 ;
        RECT 350.180 -650.175 350.560 -545.585 ;
        RECT 351.700 -645.605 352.080 -541.015 ;
        RECT 353.220 -650.175 353.600 -545.585 ;
        RECT 354.740 -645.605 355.120 -541.015 ;
        RECT 356.260 -650.175 356.640 -545.585 ;
        RECT 357.780 -645.605 358.160 -541.015 ;
        RECT 359.300 -650.175 359.680 -545.585 ;
        RECT 360.820 -645.605 361.200 -541.015 ;
        RECT 362.340 -650.175 362.720 -545.585 ;
        RECT 363.860 -645.605 364.240 -541.015 ;
        RECT 365.380 -650.175 365.760 -545.585 ;
        RECT 366.900 -645.605 367.280 -541.015 ;
        RECT 368.420 -650.175 368.800 -545.585 ;
        RECT 369.940 -645.605 370.320 -541.015 ;
        RECT 371.460 -650.175 371.840 -545.585 ;
        RECT 372.980 -645.605 373.360 -541.015 ;
        RECT 374.500 -650.175 374.880 -545.585 ;
        RECT 376.020 -645.605 376.400 -541.015 ;
        RECT 377.540 -650.175 377.920 -545.585 ;
        RECT 379.060 -645.605 379.440 -541.015 ;
        RECT 380.580 -650.175 380.960 -545.585 ;
        RECT 382.100 -645.605 382.480 -541.015 ;
        RECT 383.620 -650.175 384.000 -545.585 ;
        RECT 385.140 -645.605 385.520 -541.015 ;
        RECT 386.660 -650.175 387.040 -545.585 ;
        RECT 388.180 -645.605 388.560 -541.015 ;
        RECT 389.700 -650.175 390.080 -545.585 ;
        RECT 391.220 -645.605 391.600 -541.015 ;
        RECT 392.740 -650.175 393.120 -545.585 ;
        RECT 394.260 -645.605 394.640 -541.015 ;
        RECT 395.780 -650.175 396.160 -545.585 ;
        RECT 397.300 -645.605 397.680 -541.015 ;
        RECT 398.820 -650.175 399.200 -545.585 ;
        RECT 400.340 -645.605 400.720 -541.015 ;
        RECT 401.860 -650.175 402.240 -545.585 ;
        RECT 403.380 -645.605 403.760 -541.015 ;
        RECT 404.900 -650.175 405.280 -545.585 ;
        RECT 406.420 -645.605 406.800 -541.015 ;
        RECT 414.420 -545.595 414.800 -541.015 ;
        RECT 413.630 -645.605 414.800 -545.595 ;
        RECT 415.940 -650.175 416.320 -545.585 ;
        RECT 417.460 -645.605 417.840 -541.015 ;
        RECT 418.980 -650.175 419.360 -545.585 ;
        RECT 420.500 -645.605 420.880 -541.015 ;
        RECT 422.020 -650.175 422.400 -545.585 ;
        RECT 423.540 -645.605 423.920 -541.015 ;
        RECT 425.060 -650.175 425.440 -545.585 ;
        RECT 426.580 -645.605 426.960 -541.015 ;
        RECT 428.100 -650.175 428.480 -545.585 ;
        RECT 429.620 -645.605 430.000 -541.015 ;
        RECT 431.140 -650.175 431.520 -545.585 ;
        RECT 432.660 -645.605 433.040 -541.015 ;
        RECT 434.180 -650.175 434.560 -545.585 ;
        RECT 435.700 -645.605 436.080 -541.015 ;
        RECT 437.220 -650.175 437.600 -545.585 ;
        RECT 438.740 -645.605 439.120 -541.015 ;
        RECT 440.260 -650.175 440.640 -545.585 ;
        RECT 441.780 -645.605 442.160 -541.015 ;
        RECT 443.300 -650.175 443.680 -545.585 ;
        RECT 444.820 -645.605 445.200 -541.015 ;
        RECT 446.340 -650.175 446.720 -545.585 ;
        RECT 447.860 -645.605 448.240 -541.015 ;
        RECT 449.380 -650.175 449.760 -545.585 ;
        RECT 450.900 -645.605 451.280 -541.015 ;
        RECT 452.420 -650.175 452.800 -545.585 ;
        RECT 453.940 -645.605 454.320 -541.015 ;
        RECT 455.460 -650.175 455.840 -545.585 ;
        RECT 456.980 -645.605 457.360 -541.015 ;
        RECT 458.500 -650.175 458.880 -545.585 ;
        RECT 460.020 -645.605 460.400 -541.015 ;
        RECT 461.540 -650.175 461.920 -545.585 ;
        RECT 463.060 -645.605 463.440 -541.015 ;
        RECT 464.580 -650.175 464.960 -545.585 ;
        RECT 466.100 -645.605 466.480 -541.015 ;
        RECT 467.620 -650.175 468.000 -545.585 ;
        RECT 469.140 -645.605 469.520 -541.015 ;
        RECT 470.660 -650.175 471.040 -545.585 ;
        RECT 472.180 -645.605 472.560 -541.015 ;
        RECT 473.700 -650.175 474.080 -545.585 ;
        RECT 475.220 -645.605 475.600 -541.015 ;
        RECT 476.740 -650.175 477.120 -545.585 ;
        RECT 478.260 -645.605 478.640 -541.015 ;
        RECT 479.780 -650.175 480.160 -545.585 ;
        RECT 481.300 -645.605 481.680 -541.015 ;
        RECT 482.820 -650.175 483.200 -545.585 ;
        RECT 484.340 -645.605 484.720 -541.015 ;
        RECT 485.860 -650.175 486.240 -545.585 ;
        RECT 487.380 -645.605 487.760 -541.015 ;
        RECT 488.900 -650.175 489.280 -545.585 ;
        RECT 490.420 -645.605 490.800 -541.015 ;
        RECT 491.940 -650.175 492.320 -545.585 ;
        RECT 493.460 -645.605 493.840 -541.015 ;
        RECT 494.980 -650.175 495.360 -545.585 ;
        RECT 496.500 -645.605 496.880 -541.015 ;
        RECT 498.020 -650.175 498.400 -545.585 ;
        RECT 499.540 -645.605 499.920 -541.015 ;
        RECT 501.060 -650.175 501.440 -545.585 ;
        RECT 502.580 -645.605 502.960 -541.015 ;
        RECT 504.100 -650.175 504.480 -545.585 ;
        RECT 505.620 -645.605 506.000 -541.015 ;
        RECT 507.140 -650.175 507.520 -545.585 ;
        RECT 508.660 -645.605 509.040 -541.015 ;
        RECT 510.180 -650.175 510.560 -545.585 ;
        RECT 511.700 -645.605 512.080 -541.015 ;
        RECT 513.220 -650.175 513.600 -545.585 ;
        RECT 514.740 -645.605 515.120 -541.015 ;
        RECT 516.260 -650.175 516.640 -545.585 ;
        RECT 517.780 -645.605 518.160 -541.015 ;
        RECT 519.300 -650.175 519.680 -545.585 ;
        RECT 520.820 -645.605 521.200 -541.015 ;
        RECT 522.340 -650.175 522.720 -545.585 ;
        RECT 523.860 -645.605 524.240 -541.015 ;
        RECT 525.380 -650.175 525.760 -545.585 ;
        RECT 526.900 -645.605 527.280 -541.015 ;
        RECT 528.420 -650.175 528.800 -545.585 ;
        RECT 529.940 -645.605 530.320 -541.015 ;
        RECT 531.460 -650.175 531.840 -545.585 ;
        RECT 532.980 -645.605 533.360 -541.015 ;
        RECT 534.500 -650.175 534.880 -545.585 ;
        RECT 536.020 -645.605 536.400 -541.015 ;
        RECT 537.540 -650.175 537.920 -545.585 ;
        RECT 539.060 -645.605 539.440 -541.015 ;
        RECT 540.580 -650.175 540.960 -545.585 ;
        RECT 542.100 -645.605 542.480 -541.015 ;
        RECT 543.620 -650.175 544.000 -545.585 ;
        RECT 545.140 -645.605 545.520 -541.015 ;
        RECT 546.660 -650.175 547.040 -545.585 ;
        RECT 548.180 -645.605 548.560 -541.015 ;
        RECT 549.700 -650.175 550.080 -545.585 ;
        RECT 551.220 -645.605 551.600 -541.015 ;
        RECT 552.740 -650.175 553.120 -545.585 ;
        RECT 554.260 -645.605 554.640 -541.015 ;
        RECT 555.780 -650.175 556.160 -545.585 ;
        RECT 557.300 -645.605 557.680 -541.015 ;
        RECT 558.820 -650.175 559.200 -545.585 ;
        RECT 560.340 -645.605 560.720 -541.015 ;
        RECT 561.860 -650.175 562.240 -545.585 ;
        RECT 563.380 -645.605 563.760 -541.015 ;
        RECT 564.900 -650.175 565.280 -545.585 ;
        RECT 566.420 -645.605 566.800 -541.015 ;
        RECT 574.420 -545.595 574.800 -541.015 ;
        RECT 573.630 -645.605 574.800 -545.595 ;
        RECT 575.940 -650.175 576.320 -545.585 ;
        RECT 577.460 -645.605 577.840 -541.015 ;
        RECT 578.980 -650.175 579.360 -545.585 ;
        RECT 580.500 -645.605 580.880 -541.015 ;
        RECT 582.020 -650.175 582.400 -545.585 ;
        RECT 583.540 -645.605 583.920 -541.015 ;
        RECT 585.060 -650.175 585.440 -545.585 ;
        RECT 586.580 -645.605 586.960 -541.015 ;
        RECT 588.100 -650.175 588.480 -545.585 ;
        RECT 589.620 -645.605 590.000 -541.015 ;
        RECT 591.140 -650.175 591.520 -545.585 ;
        RECT 592.660 -645.605 593.040 -541.015 ;
        RECT 594.180 -650.175 594.560 -545.585 ;
        RECT 595.700 -645.605 596.080 -541.015 ;
        RECT 597.220 -650.175 597.600 -545.585 ;
        RECT 598.740 -645.605 599.120 -541.015 ;
        RECT 600.260 -650.175 600.640 -545.585 ;
        RECT 601.780 -645.605 602.160 -541.015 ;
        RECT 603.300 -650.175 603.680 -545.585 ;
        RECT 604.820 -645.605 605.200 -541.015 ;
        RECT 606.340 -650.175 606.720 -545.585 ;
        RECT 607.860 -645.605 608.240 -541.015 ;
        RECT 609.380 -650.175 609.760 -545.585 ;
        RECT 610.900 -645.605 611.280 -541.015 ;
        RECT 612.420 -650.175 612.800 -545.585 ;
        RECT 613.940 -645.605 614.320 -541.015 ;
        RECT 615.460 -650.175 615.840 -545.585 ;
        RECT 616.980 -645.605 617.360 -541.015 ;
        RECT 618.500 -650.175 618.880 -545.585 ;
        RECT 620.020 -645.605 620.400 -541.015 ;
        RECT 621.540 -650.175 621.920 -545.585 ;
        RECT 623.060 -645.605 623.440 -541.015 ;
        RECT 624.580 -650.175 624.960 -545.585 ;
        RECT 626.100 -645.605 626.480 -541.015 ;
        RECT 627.620 -650.175 628.000 -545.585 ;
        RECT 629.140 -645.605 629.520 -541.015 ;
        RECT 630.660 -650.175 631.040 -545.585 ;
        RECT 632.180 -645.605 632.560 -541.015 ;
        RECT 633.700 -650.175 634.080 -545.585 ;
        RECT 635.220 -645.605 635.600 -541.015 ;
        RECT 636.740 -650.175 637.120 -545.585 ;
        RECT 638.260 -645.605 638.640 -541.015 ;
        RECT 639.780 -650.175 640.160 -545.585 ;
        RECT 641.300 -645.605 641.680 -541.015 ;
        RECT 642.820 -650.175 643.200 -545.585 ;
        RECT 644.340 -645.605 644.720 -541.015 ;
        RECT 645.860 -650.175 646.240 -545.585 ;
        RECT 647.380 -645.605 647.760 -541.015 ;
        RECT 648.900 -650.175 649.280 -545.585 ;
        RECT 650.420 -645.605 650.800 -541.015 ;
        RECT 651.940 -650.175 652.320 -545.585 ;
        RECT 653.460 -645.605 653.840 -541.015 ;
        RECT 654.980 -650.175 655.360 -545.585 ;
        RECT 656.500 -645.605 656.880 -541.015 ;
        RECT 658.020 -650.175 658.400 -545.585 ;
        RECT 659.540 -645.605 659.920 -541.015 ;
        RECT 661.060 -650.175 661.440 -545.585 ;
        RECT 662.580 -645.605 662.960 -541.015 ;
        RECT 664.100 -650.175 664.480 -545.585 ;
        RECT 665.620 -645.605 666.000 -541.015 ;
        RECT 667.140 -650.175 667.520 -545.585 ;
        RECT 668.660 -645.605 669.040 -541.015 ;
        RECT 670.180 -650.175 670.560 -545.585 ;
        RECT 671.700 -645.605 672.080 -541.015 ;
        RECT 673.220 -650.175 673.600 -545.585 ;
        RECT 674.740 -645.605 675.120 -541.015 ;
        RECT 676.260 -650.175 676.640 -545.585 ;
        RECT 677.780 -645.605 678.160 -541.015 ;
        RECT 679.300 -650.175 679.680 -545.585 ;
        RECT 680.820 -645.605 681.200 -541.015 ;
        RECT 682.340 -650.175 682.720 -545.585 ;
        RECT 683.860 -645.605 684.240 -541.015 ;
        RECT 685.380 -650.175 685.760 -545.585 ;
        RECT 686.900 -645.605 687.280 -541.015 ;
        RECT 688.420 -650.175 688.800 -545.585 ;
        RECT 689.940 -645.605 690.320 -541.015 ;
        RECT 691.460 -650.175 691.840 -545.585 ;
        RECT 692.980 -645.605 693.360 -541.015 ;
        RECT 694.500 -650.175 694.880 -545.585 ;
        RECT 696.020 -645.605 696.400 -541.015 ;
        RECT 697.540 -650.175 697.920 -545.585 ;
        RECT 699.060 -645.605 699.440 -541.015 ;
        RECT 700.580 -650.175 700.960 -545.585 ;
        RECT 702.100 -645.605 702.480 -541.015 ;
        RECT 703.620 -650.175 704.000 -545.585 ;
        RECT 705.140 -645.605 705.520 -541.015 ;
        RECT 706.660 -650.175 707.040 -545.585 ;
        RECT 708.180 -645.605 708.560 -541.015 ;
        RECT 709.700 -650.175 710.080 -545.585 ;
        RECT 711.220 -645.605 711.600 -541.015 ;
        RECT 712.740 -650.175 713.120 -545.585 ;
        RECT 714.260 -645.605 714.640 -541.015 ;
        RECT 715.780 -650.175 716.160 -545.585 ;
        RECT 717.300 -645.605 717.680 -541.015 ;
        RECT 718.820 -650.175 719.200 -545.585 ;
        RECT 720.340 -645.605 720.720 -541.015 ;
        RECT 721.860 -650.175 722.240 -545.585 ;
        RECT 723.380 -645.605 723.760 -541.015 ;
        RECT 724.900 -650.175 725.280 -545.585 ;
        RECT 726.420 -645.605 726.800 -541.015 ;
        RECT 734.420 -545.595 734.800 -541.015 ;
        RECT 733.630 -645.605 734.800 -545.595 ;
        RECT 735.940 -650.175 736.320 -545.585 ;
        RECT 737.460 -645.605 737.840 -541.015 ;
        RECT 738.980 -650.175 739.360 -545.585 ;
        RECT 740.500 -645.605 740.880 -541.015 ;
        RECT 742.020 -650.175 742.400 -545.585 ;
        RECT 743.540 -645.605 743.920 -541.015 ;
        RECT 745.060 -650.175 745.440 -545.585 ;
        RECT 746.580 -645.605 746.960 -541.015 ;
        RECT 748.100 -650.175 748.480 -545.585 ;
        RECT 749.620 -645.605 750.000 -541.015 ;
        RECT 751.140 -650.175 751.520 -545.585 ;
        RECT 752.660 -645.605 753.040 -541.015 ;
        RECT 754.180 -650.175 754.560 -545.585 ;
        RECT 755.700 -645.605 756.080 -541.015 ;
        RECT 757.220 -650.175 757.600 -545.585 ;
        RECT 758.740 -645.605 759.120 -541.015 ;
        RECT 760.260 -650.175 760.640 -545.585 ;
        RECT 761.780 -645.605 762.160 -541.015 ;
        RECT 763.300 -650.175 763.680 -545.585 ;
        RECT 764.820 -645.605 765.200 -541.015 ;
        RECT 766.340 -650.175 766.720 -545.585 ;
        RECT 767.860 -645.605 768.240 -541.015 ;
        RECT 769.380 -650.175 769.760 -545.585 ;
        RECT 770.900 -645.605 771.280 -541.015 ;
        RECT 772.420 -650.175 772.800 -545.585 ;
        RECT 773.940 -645.605 774.320 -541.015 ;
        RECT 775.460 -650.175 775.840 -545.585 ;
        RECT 776.980 -645.605 777.360 -541.015 ;
        RECT 778.500 -650.175 778.880 -545.585 ;
        RECT 780.020 -645.605 780.400 -541.015 ;
        RECT 781.540 -650.175 781.920 -545.585 ;
        RECT 783.060 -645.605 783.440 -541.015 ;
        RECT 784.580 -650.175 784.960 -545.585 ;
        RECT 786.100 -645.605 786.480 -541.015 ;
        RECT 787.620 -650.175 788.000 -545.585 ;
        RECT 789.140 -645.605 789.520 -541.015 ;
        RECT 790.660 -650.175 791.040 -545.585 ;
        RECT 792.180 -645.605 792.560 -541.015 ;
        RECT 793.700 -650.175 794.080 -545.585 ;
        RECT 795.220 -645.605 795.600 -541.015 ;
        RECT 796.740 -650.175 797.120 -545.585 ;
        RECT 798.260 -645.605 798.640 -541.015 ;
        RECT 799.780 -650.175 800.160 -545.585 ;
        RECT 801.300 -645.605 801.680 -541.015 ;
        RECT 802.820 -650.175 803.200 -545.585 ;
        RECT 804.340 -645.605 804.720 -541.015 ;
        RECT 805.860 -650.175 806.240 -545.585 ;
        RECT 807.380 -645.605 807.760 -541.015 ;
        RECT 808.900 -650.175 809.280 -545.585 ;
        RECT 810.420 -645.605 810.800 -541.015 ;
        RECT 811.940 -650.175 812.320 -545.585 ;
        RECT 813.460 -645.605 813.840 -541.015 ;
        RECT 814.980 -650.175 815.360 -545.585 ;
        RECT 816.500 -645.605 816.880 -541.015 ;
        RECT 818.020 -650.175 818.400 -545.585 ;
        RECT 819.540 -645.605 819.920 -541.015 ;
        RECT 821.060 -650.175 821.440 -545.585 ;
        RECT 822.580 -645.605 822.960 -541.015 ;
        RECT 824.100 -650.175 824.480 -545.585 ;
        RECT 825.620 -645.605 826.000 -541.015 ;
        RECT 827.140 -650.175 827.520 -545.585 ;
        RECT 828.660 -645.605 829.040 -541.015 ;
        RECT 830.180 -650.175 830.560 -545.585 ;
        RECT 831.700 -645.605 832.080 -541.015 ;
        RECT 833.220 -650.175 833.600 -545.585 ;
        RECT 834.740 -645.605 835.120 -541.015 ;
        RECT 836.260 -650.175 836.640 -545.585 ;
        RECT 837.780 -645.605 838.160 -541.015 ;
        RECT 839.300 -650.175 839.680 -545.585 ;
        RECT 840.820 -645.605 841.200 -541.015 ;
        RECT 842.340 -650.175 842.720 -545.585 ;
        RECT 843.860 -645.605 844.240 -541.015 ;
        RECT 845.380 -650.175 845.760 -545.585 ;
        RECT 846.900 -645.605 847.280 -541.015 ;
        RECT 848.420 -650.175 848.800 -545.585 ;
        RECT 849.940 -645.605 850.320 -541.015 ;
        RECT 851.460 -650.175 851.840 -545.585 ;
        RECT 852.980 -645.605 853.360 -541.015 ;
        RECT 854.500 -650.175 854.880 -545.585 ;
        RECT 856.020 -645.605 856.400 -541.015 ;
        RECT 857.540 -650.175 857.920 -545.585 ;
        RECT 859.060 -645.605 859.440 -541.015 ;
        RECT 860.580 -650.175 860.960 -545.585 ;
        RECT 862.100 -645.605 862.480 -541.015 ;
        RECT 863.620 -650.175 864.000 -545.585 ;
        RECT 865.140 -645.605 865.520 -541.015 ;
        RECT 866.660 -650.175 867.040 -545.585 ;
        RECT 868.180 -645.605 868.560 -541.015 ;
        RECT 869.700 -650.175 870.080 -545.585 ;
        RECT 871.220 -645.605 871.600 -541.015 ;
        RECT 872.740 -650.175 873.120 -545.585 ;
        RECT 874.260 -645.605 874.640 -541.015 ;
        RECT 875.780 -650.175 876.160 -545.585 ;
        RECT 877.300 -645.605 877.680 -541.015 ;
        RECT 878.820 -650.175 879.200 -545.585 ;
        RECT 880.340 -645.605 880.720 -541.015 ;
        RECT 881.860 -650.175 882.240 -545.585 ;
        RECT 883.380 -645.605 883.760 -541.015 ;
        RECT 884.900 -650.175 885.280 -545.585 ;
        RECT 886.420 -645.605 886.800 -541.015 ;
        RECT 888.320 -650.175 891.540 -523.010 ;
        RECT -544.060 -653.010 891.540 -650.175 ;
        RECT -544.060 -669.335 888.320 -653.010 ;
        RECT -535.705 -856.395 -527.940 -693.905 ;
        RECT -526.800 -722.750 -479.475 -672.845 ;
        RECT -429.865 -718.750 -362.530 -691.350 ;
        RECT -516.635 -749.870 -398.300 -743.830 ;
        RECT -516.635 -813.425 -489.500 -749.870 ;
        RECT -516.635 -856.395 -490.670 -813.425 ;
        RECT -488.360 -816.960 -487.980 -753.405 ;
        RECT -486.840 -813.425 -486.460 -749.870 ;
        RECT -485.320 -816.960 -484.940 -753.405 ;
        RECT -483.800 -813.425 -483.420 -749.870 ;
        RECT -482.280 -816.960 -481.900 -753.405 ;
        RECT -480.760 -813.425 -480.380 -749.870 ;
        RECT -479.240 -816.960 -478.860 -753.405 ;
        RECT -477.720 -813.425 -477.340 -749.870 ;
        RECT -476.200 -816.960 -475.820 -753.405 ;
        RECT -474.680 -813.425 -474.300 -749.870 ;
        RECT -473.160 -816.960 -472.780 -753.405 ;
        RECT -471.640 -813.425 -471.260 -749.870 ;
        RECT -470.120 -816.960 -469.740 -753.405 ;
        RECT -468.600 -813.425 -468.220 -749.870 ;
        RECT -467.080 -816.960 -466.700 -753.405 ;
        RECT -465.560 -813.425 -465.180 -749.870 ;
        RECT -464.040 -816.960 -463.660 -753.405 ;
        RECT -462.520 -813.425 -462.140 -749.870 ;
        RECT -461.000 -816.960 -460.620 -753.405 ;
        RECT -459.480 -813.425 -459.100 -749.870 ;
        RECT -457.960 -816.960 -457.580 -753.405 ;
        RECT -456.440 -813.425 -456.060 -749.870 ;
        RECT -454.920 -816.960 -454.540 -753.405 ;
        RECT -453.400 -813.425 -453.020 -749.870 ;
        RECT -451.880 -816.960 -451.500 -753.405 ;
        RECT -450.360 -813.425 -449.980 -749.870 ;
        RECT -448.840 -816.960 -448.460 -753.405 ;
        RECT -447.320 -813.425 -446.940 -749.870 ;
        RECT -445.800 -816.960 -445.420 -753.405 ;
        RECT -444.280 -813.425 -443.900 -749.870 ;
        RECT -442.760 -816.960 -442.380 -753.405 ;
        RECT -441.240 -813.425 -440.860 -749.870 ;
        RECT -439.720 -816.960 -439.340 -753.405 ;
        RECT -438.200 -813.425 -437.820 -749.870 ;
        RECT -436.680 -816.960 -436.300 -753.405 ;
        RECT -435.160 -813.425 -434.780 -749.870 ;
        RECT -433.640 -816.960 -433.260 -753.405 ;
        RECT -432.120 -813.425 -431.740 -749.870 ;
        RECT -430.600 -816.960 -430.220 -753.405 ;
        RECT -429.080 -813.425 -428.700 -749.870 ;
        RECT -427.560 -816.960 -427.180 -753.405 ;
        RECT -426.040 -813.425 -425.660 -749.870 ;
        RECT -424.520 -816.960 -424.140 -753.405 ;
        RECT -423.000 -813.425 -422.620 -749.870 ;
        RECT -421.480 -816.960 -421.100 -753.405 ;
        RECT -419.960 -813.425 -419.580 -749.870 ;
        RECT -418.440 -816.960 -418.060 -753.405 ;
        RECT -416.920 -813.425 -416.540 -749.870 ;
        RECT -415.400 -816.960 -415.020 -753.405 ;
        RECT -413.880 -813.425 -413.500 -749.870 ;
        RECT -412.360 -816.960 -411.980 -753.405 ;
        RECT -410.840 -813.425 -410.460 -749.870 ;
        RECT -409.320 -816.960 -408.940 -753.405 ;
        RECT -407.800 -813.425 -407.420 -749.870 ;
        RECT -406.280 -816.960 -405.900 -753.405 ;
        RECT -404.760 -813.425 -404.380 -749.870 ;
        RECT -403.240 -816.960 -402.860 -753.405 ;
        RECT -401.720 -813.425 -401.340 -749.870 ;
        RECT -400.200 -816.960 -399.820 -753.405 ;
        RECT -398.680 -813.425 -398.300 -749.870 ;
        RECT -388.355 -816.960 -362.530 -718.750 ;
        RECT -301.280 -705.535 871.890 -680.075 ;
        RECT -301.280 -811.760 -300.110 -705.535 ;
        RECT -300.490 -811.770 -300.110 -811.760 ;
        RECT -488.360 -823.000 -362.530 -816.960 ;
        RECT -298.970 -817.985 -298.590 -711.750 ;
        RECT -297.450 -811.770 -297.070 -705.535 ;
        RECT -295.930 -817.985 -295.550 -711.750 ;
        RECT -294.410 -811.770 -294.030 -705.535 ;
        RECT -292.890 -817.985 -292.510 -711.750 ;
        RECT -291.370 -811.770 -290.990 -705.535 ;
        RECT -289.850 -817.985 -289.470 -711.750 ;
        RECT -288.330 -811.770 -287.950 -705.535 ;
        RECT -286.810 -817.985 -286.430 -711.750 ;
        RECT -285.290 -811.770 -284.910 -705.535 ;
        RECT -283.770 -817.985 -283.390 -711.750 ;
        RECT -282.250 -811.770 -281.870 -705.535 ;
        RECT -280.730 -817.985 -280.350 -711.750 ;
        RECT -279.210 -811.770 -278.830 -705.535 ;
        RECT -277.690 -817.985 -277.310 -711.750 ;
        RECT -276.170 -811.770 -275.790 -705.535 ;
        RECT -274.650 -817.985 -274.270 -711.750 ;
        RECT -273.130 -811.770 -272.750 -705.535 ;
        RECT -271.610 -817.985 -271.230 -711.750 ;
        RECT -270.090 -811.770 -269.710 -705.535 ;
        RECT -268.570 -817.985 -268.190 -711.750 ;
        RECT -267.050 -811.770 -266.670 -705.535 ;
        RECT -265.530 -817.985 -265.150 -711.750 ;
        RECT -264.010 -811.770 -263.630 -705.535 ;
        RECT -262.490 -817.985 -262.110 -711.750 ;
        RECT -260.970 -811.770 -260.590 -705.535 ;
        RECT -259.450 -817.985 -259.070 -711.750 ;
        RECT -257.930 -811.770 -257.550 -705.535 ;
        RECT -256.410 -817.985 -256.030 -711.750 ;
        RECT -254.890 -811.770 -254.510 -705.535 ;
        RECT -253.370 -817.985 -252.990 -711.750 ;
        RECT -251.850 -811.770 -251.470 -705.535 ;
        RECT -250.330 -817.985 -249.950 -711.750 ;
        RECT -248.810 -811.770 -248.430 -705.535 ;
        RECT -247.290 -817.985 -246.910 -711.750 ;
        RECT -245.770 -811.770 -245.390 -705.535 ;
        RECT -244.250 -817.985 -243.870 -711.750 ;
        RECT -242.730 -811.770 -242.350 -705.535 ;
        RECT -241.210 -817.985 -240.830 -711.750 ;
        RECT -239.690 -811.770 -239.310 -705.535 ;
        RECT -238.170 -817.985 -237.790 -711.750 ;
        RECT -236.650 -811.770 -236.270 -705.535 ;
        RECT -235.130 -817.985 -234.750 -711.750 ;
        RECT -233.610 -811.770 -233.230 -705.535 ;
        RECT -232.090 -817.985 -231.710 -711.750 ;
        RECT -230.570 -811.770 -230.190 -705.535 ;
        RECT -229.050 -817.985 -228.670 -711.750 ;
        RECT -227.530 -811.770 -227.150 -705.535 ;
        RECT -226.010 -817.985 -225.630 -711.750 ;
        RECT -224.490 -811.770 -224.110 -705.535 ;
        RECT -222.970 -817.985 -222.590 -711.750 ;
        RECT -221.450 -811.770 -221.070 -705.535 ;
        RECT -219.930 -817.985 -219.550 -711.750 ;
        RECT -218.410 -811.770 -218.030 -705.535 ;
        RECT -216.890 -817.985 -216.510 -711.750 ;
        RECT -215.370 -811.770 -214.990 -705.535 ;
        RECT -213.850 -817.985 -213.470 -711.750 ;
        RECT -212.330 -811.770 -211.950 -705.535 ;
        RECT -210.810 -817.985 -210.430 -711.750 ;
        RECT -209.290 -811.770 -208.910 -705.535 ;
        RECT -207.770 -817.985 -207.390 -711.750 ;
        RECT -206.250 -811.770 -205.870 -705.535 ;
        RECT -204.730 -817.985 -204.350 -711.750 ;
        RECT -203.210 -811.770 -202.830 -705.535 ;
        RECT -201.690 -817.985 -201.310 -711.750 ;
        RECT -200.170 -811.770 -199.790 -705.535 ;
        RECT -198.650 -817.985 -198.270 -711.750 ;
        RECT -197.130 -811.770 -196.750 -705.535 ;
        RECT -195.610 -817.985 -195.230 -711.750 ;
        RECT -194.090 -811.770 -193.710 -705.535 ;
        RECT -192.570 -817.985 -192.190 -711.750 ;
        RECT -191.050 -811.770 -190.670 -705.535 ;
        RECT -189.530 -817.985 -189.150 -711.750 ;
        RECT -188.010 -811.770 -187.630 -705.535 ;
        RECT -186.490 -817.985 -186.110 -711.750 ;
        RECT -184.970 -811.770 -184.590 -705.535 ;
        RECT -183.450 -817.985 -183.070 -711.750 ;
        RECT -181.930 -811.770 -181.550 -705.535 ;
        RECT -180.410 -817.985 -180.030 -711.750 ;
        RECT -178.890 -811.770 -178.510 -705.535 ;
        RECT -177.370 -817.985 -176.990 -711.750 ;
        RECT -175.850 -811.770 -175.470 -705.535 ;
        RECT -174.330 -817.985 -173.950 -711.750 ;
        RECT -172.810 -811.770 -172.430 -705.535 ;
        RECT -171.290 -817.985 -170.910 -711.750 ;
        RECT -169.770 -811.770 -169.390 -705.535 ;
        RECT -168.250 -817.985 -167.870 -711.750 ;
        RECT -166.730 -811.770 -166.350 -705.535 ;
        RECT -165.210 -817.985 -164.830 -711.750 ;
        RECT -163.690 -811.770 -163.310 -705.535 ;
        RECT -162.170 -817.985 -161.790 -711.750 ;
        RECT -160.650 -811.770 -160.270 -705.535 ;
        RECT -159.130 -817.985 -158.750 -711.750 ;
        RECT -157.610 -811.770 -157.230 -705.535 ;
        RECT -156.090 -817.985 -155.710 -711.750 ;
        RECT -154.570 -811.770 -154.190 -705.535 ;
        RECT -153.050 -817.985 -152.670 -711.750 ;
        RECT -151.530 -811.770 -151.150 -705.535 ;
        RECT -150.010 -817.985 -149.630 -711.750 ;
        RECT -148.490 -811.770 -148.110 -705.535 ;
        RECT -131.280 -811.760 -130.110 -705.535 ;
        RECT -130.490 -811.770 -130.110 -811.760 ;
        RECT -128.970 -817.985 -128.590 -711.750 ;
        RECT -127.450 -811.770 -127.070 -705.535 ;
        RECT -125.930 -817.985 -125.550 -711.750 ;
        RECT -124.410 -811.770 -124.030 -705.535 ;
        RECT -122.890 -817.985 -122.510 -711.750 ;
        RECT -121.370 -811.770 -120.990 -705.535 ;
        RECT -119.850 -817.985 -119.470 -711.750 ;
        RECT -118.330 -811.770 -117.950 -705.535 ;
        RECT -116.810 -817.985 -116.430 -711.750 ;
        RECT -115.290 -811.770 -114.910 -705.535 ;
        RECT -113.770 -817.985 -113.390 -711.750 ;
        RECT -112.250 -811.770 -111.870 -705.535 ;
        RECT -110.730 -817.985 -110.350 -711.750 ;
        RECT -109.210 -811.770 -108.830 -705.535 ;
        RECT -107.690 -817.985 -107.310 -711.750 ;
        RECT -106.170 -811.770 -105.790 -705.535 ;
        RECT -104.650 -817.985 -104.270 -711.750 ;
        RECT -103.130 -811.770 -102.750 -705.535 ;
        RECT -101.610 -817.985 -101.230 -711.750 ;
        RECT -100.090 -811.770 -99.710 -705.535 ;
        RECT -98.570 -817.985 -98.190 -711.750 ;
        RECT -97.050 -811.770 -96.670 -705.535 ;
        RECT -95.530 -817.985 -95.150 -711.750 ;
        RECT -94.010 -811.770 -93.630 -705.535 ;
        RECT -92.490 -817.985 -92.110 -711.750 ;
        RECT -90.970 -811.770 -90.590 -705.535 ;
        RECT -89.450 -817.985 -89.070 -711.750 ;
        RECT -87.930 -811.770 -87.550 -705.535 ;
        RECT -86.410 -817.985 -86.030 -711.750 ;
        RECT -84.890 -811.770 -84.510 -705.535 ;
        RECT -83.370 -817.985 -82.990 -711.750 ;
        RECT -81.850 -811.770 -81.470 -705.535 ;
        RECT -80.330 -817.985 -79.950 -711.750 ;
        RECT -78.810 -811.770 -78.430 -705.535 ;
        RECT -77.290 -817.985 -76.910 -711.750 ;
        RECT -75.770 -811.770 -75.390 -705.535 ;
        RECT -74.250 -817.985 -73.870 -711.750 ;
        RECT -72.730 -811.770 -72.350 -705.535 ;
        RECT -71.210 -817.985 -70.830 -711.750 ;
        RECT -69.690 -811.770 -69.310 -705.535 ;
        RECT -68.170 -817.985 -67.790 -711.750 ;
        RECT -66.650 -811.770 -66.270 -705.535 ;
        RECT -65.130 -817.985 -64.750 -711.750 ;
        RECT -63.610 -811.770 -63.230 -705.535 ;
        RECT -62.090 -817.985 -61.710 -711.750 ;
        RECT -60.570 -811.770 -60.190 -705.535 ;
        RECT -59.050 -817.985 -58.670 -711.750 ;
        RECT -57.530 -811.770 -57.150 -705.535 ;
        RECT -56.010 -817.985 -55.630 -711.750 ;
        RECT -54.490 -811.770 -54.110 -705.535 ;
        RECT -52.970 -817.985 -52.590 -711.750 ;
        RECT -51.450 -811.770 -51.070 -705.535 ;
        RECT -49.930 -817.985 -49.550 -711.750 ;
        RECT -48.410 -811.770 -48.030 -705.535 ;
        RECT -46.890 -817.985 -46.510 -711.750 ;
        RECT -45.370 -811.770 -44.990 -705.535 ;
        RECT -43.850 -817.985 -43.470 -711.750 ;
        RECT -42.330 -811.770 -41.950 -705.535 ;
        RECT -40.810 -817.985 -40.430 -711.750 ;
        RECT -39.290 -811.770 -38.910 -705.535 ;
        RECT -37.770 -817.985 -37.390 -711.750 ;
        RECT -36.250 -811.770 -35.870 -705.535 ;
        RECT -34.730 -817.985 -34.350 -711.750 ;
        RECT -33.210 -811.770 -32.830 -705.535 ;
        RECT -31.690 -817.985 -31.310 -711.750 ;
        RECT -30.170 -811.770 -29.790 -705.535 ;
        RECT -28.650 -817.985 -28.270 -711.750 ;
        RECT -27.130 -811.770 -26.750 -705.535 ;
        RECT -25.610 -817.985 -25.230 -711.750 ;
        RECT -24.090 -811.770 -23.710 -705.535 ;
        RECT -22.570 -817.985 -22.190 -711.750 ;
        RECT -21.050 -811.770 -20.670 -705.535 ;
        RECT -19.530 -817.985 -19.150 -711.750 ;
        RECT -18.010 -811.770 -17.630 -705.535 ;
        RECT -16.490 -817.985 -16.110 -711.750 ;
        RECT -14.970 -811.770 -14.590 -705.535 ;
        RECT -13.450 -817.985 -13.070 -711.750 ;
        RECT -11.930 -811.770 -11.550 -705.535 ;
        RECT -10.410 -817.985 -10.030 -711.750 ;
        RECT -8.890 -811.770 -8.510 -705.535 ;
        RECT -7.370 -817.985 -6.990 -711.750 ;
        RECT -5.850 -811.770 -5.470 -705.535 ;
        RECT -4.330 -817.985 -3.950 -711.750 ;
        RECT -2.810 -811.770 -2.430 -705.535 ;
        RECT -1.290 -817.985 -0.910 -711.750 ;
        RECT 0.230 -811.770 0.610 -705.535 ;
        RECT 1.750 -817.985 2.130 -711.750 ;
        RECT 3.270 -811.770 3.650 -705.535 ;
        RECT 4.790 -817.985 5.170 -711.750 ;
        RECT 6.310 -811.770 6.690 -705.535 ;
        RECT 7.830 -817.985 8.210 -711.750 ;
        RECT 9.350 -811.770 9.730 -705.535 ;
        RECT 10.870 -817.985 11.250 -711.750 ;
        RECT 12.390 -811.770 12.770 -705.535 ;
        RECT 13.910 -817.985 14.290 -711.750 ;
        RECT 15.430 -811.770 15.810 -705.535 ;
        RECT 16.950 -817.985 17.330 -711.750 ;
        RECT 18.470 -811.770 18.850 -705.535 ;
        RECT 19.990 -817.985 20.370 -711.750 ;
        RECT 21.510 -811.770 21.890 -705.535 ;
        RECT 38.720 -811.760 39.890 -705.535 ;
        RECT 39.510 -811.770 39.890 -811.760 ;
        RECT 41.030 -817.985 41.410 -711.750 ;
        RECT 42.550 -811.770 42.930 -705.535 ;
        RECT 44.070 -817.985 44.450 -711.750 ;
        RECT 45.590 -811.770 45.970 -705.535 ;
        RECT 47.110 -817.985 47.490 -711.750 ;
        RECT 48.630 -811.770 49.010 -705.535 ;
        RECT 50.150 -817.985 50.530 -711.750 ;
        RECT 51.670 -811.770 52.050 -705.535 ;
        RECT 53.190 -817.985 53.570 -711.750 ;
        RECT 54.710 -811.770 55.090 -705.535 ;
        RECT 56.230 -817.985 56.610 -711.750 ;
        RECT 57.750 -811.770 58.130 -705.535 ;
        RECT 59.270 -817.985 59.650 -711.750 ;
        RECT 60.790 -811.770 61.170 -705.535 ;
        RECT 62.310 -817.985 62.690 -711.750 ;
        RECT 63.830 -811.770 64.210 -705.535 ;
        RECT 65.350 -817.985 65.730 -711.750 ;
        RECT 66.870 -811.770 67.250 -705.535 ;
        RECT 68.390 -817.985 68.770 -711.750 ;
        RECT 69.910 -811.770 70.290 -705.535 ;
        RECT 71.430 -817.985 71.810 -711.750 ;
        RECT 72.950 -811.770 73.330 -705.535 ;
        RECT 74.470 -817.985 74.850 -711.750 ;
        RECT 75.990 -811.770 76.370 -705.535 ;
        RECT 77.510 -817.985 77.890 -711.750 ;
        RECT 79.030 -811.770 79.410 -705.535 ;
        RECT 80.550 -817.985 80.930 -711.750 ;
        RECT 82.070 -811.770 82.450 -705.535 ;
        RECT 83.590 -817.985 83.970 -711.750 ;
        RECT 85.110 -811.770 85.490 -705.535 ;
        RECT 86.630 -817.985 87.010 -711.750 ;
        RECT 88.150 -811.770 88.530 -705.535 ;
        RECT 89.670 -817.985 90.050 -711.750 ;
        RECT 91.190 -811.770 91.570 -705.535 ;
        RECT 92.710 -817.985 93.090 -711.750 ;
        RECT 94.230 -811.770 94.610 -705.535 ;
        RECT 95.750 -817.985 96.130 -711.750 ;
        RECT 97.270 -811.770 97.650 -705.535 ;
        RECT 98.790 -817.985 99.170 -711.750 ;
        RECT 100.310 -811.770 100.690 -705.535 ;
        RECT 101.830 -817.985 102.210 -711.750 ;
        RECT 103.350 -811.770 103.730 -705.535 ;
        RECT 104.870 -817.985 105.250 -711.750 ;
        RECT 106.390 -811.770 106.770 -705.535 ;
        RECT 107.910 -817.985 108.290 -711.750 ;
        RECT 109.430 -811.770 109.810 -705.535 ;
        RECT 110.950 -817.985 111.330 -711.750 ;
        RECT 112.470 -811.770 112.850 -705.535 ;
        RECT 113.990 -817.985 114.370 -711.750 ;
        RECT 115.510 -811.770 115.890 -705.535 ;
        RECT 117.030 -817.985 117.410 -711.750 ;
        RECT 118.550 -811.770 118.930 -705.535 ;
        RECT 120.070 -817.985 120.450 -711.750 ;
        RECT 121.590 -811.770 121.970 -705.535 ;
        RECT 123.110 -817.985 123.490 -711.750 ;
        RECT 124.630 -811.770 125.010 -705.535 ;
        RECT 126.150 -817.985 126.530 -711.750 ;
        RECT 127.670 -811.770 128.050 -705.535 ;
        RECT 129.190 -817.985 129.570 -711.750 ;
        RECT 130.710 -811.770 131.090 -705.535 ;
        RECT 132.230 -817.985 132.610 -711.750 ;
        RECT 133.750 -811.770 134.130 -705.535 ;
        RECT 135.270 -817.985 135.650 -711.750 ;
        RECT 136.790 -811.770 137.170 -705.535 ;
        RECT 138.310 -817.985 138.690 -711.750 ;
        RECT 139.830 -811.770 140.210 -705.535 ;
        RECT 141.350 -817.985 141.730 -711.750 ;
        RECT 142.870 -811.770 143.250 -705.535 ;
        RECT 144.390 -817.985 144.770 -711.750 ;
        RECT 145.910 -811.770 146.290 -705.535 ;
        RECT 147.430 -817.985 147.810 -711.750 ;
        RECT 148.950 -811.770 149.330 -705.535 ;
        RECT 150.470 -817.985 150.850 -711.750 ;
        RECT 151.990 -811.770 152.370 -705.535 ;
        RECT 153.510 -817.985 153.890 -711.750 ;
        RECT 155.030 -811.770 155.410 -705.535 ;
        RECT 156.550 -817.985 156.930 -711.750 ;
        RECT 158.070 -811.770 158.450 -705.535 ;
        RECT 159.590 -817.985 159.970 -711.750 ;
        RECT 161.110 -811.770 161.490 -705.535 ;
        RECT 162.630 -817.985 163.010 -711.750 ;
        RECT 164.150 -811.770 164.530 -705.535 ;
        RECT 165.670 -817.985 166.050 -711.750 ;
        RECT 167.190 -811.770 167.570 -705.535 ;
        RECT 168.710 -817.985 169.090 -711.750 ;
        RECT 170.230 -811.770 170.610 -705.535 ;
        RECT 171.750 -817.985 172.130 -711.750 ;
        RECT 173.270 -811.770 173.650 -705.535 ;
        RECT 174.790 -817.985 175.170 -711.750 ;
        RECT 176.310 -811.770 176.690 -705.535 ;
        RECT 177.830 -817.985 178.210 -711.750 ;
        RECT 179.350 -811.770 179.730 -705.535 ;
        RECT 180.870 -817.985 181.250 -711.750 ;
        RECT 182.390 -811.770 182.770 -705.535 ;
        RECT 183.910 -817.985 184.290 -711.750 ;
        RECT 185.430 -811.770 185.810 -705.535 ;
        RECT 186.950 -817.985 187.330 -711.750 ;
        RECT 188.470 -811.770 188.850 -705.535 ;
        RECT 189.990 -817.985 190.370 -711.750 ;
        RECT 191.510 -811.770 191.890 -705.535 ;
        RECT 208.720 -811.760 209.890 -705.535 ;
        RECT 209.510 -811.770 209.890 -811.760 ;
        RECT 211.030 -817.985 211.410 -711.750 ;
        RECT 212.550 -811.770 212.930 -705.535 ;
        RECT 214.070 -817.985 214.450 -711.750 ;
        RECT 215.590 -811.770 215.970 -705.535 ;
        RECT 217.110 -817.985 217.490 -711.750 ;
        RECT 218.630 -811.770 219.010 -705.535 ;
        RECT 220.150 -817.985 220.530 -711.750 ;
        RECT 221.670 -811.770 222.050 -705.535 ;
        RECT 223.190 -817.985 223.570 -711.750 ;
        RECT 224.710 -811.770 225.090 -705.535 ;
        RECT 226.230 -817.985 226.610 -711.750 ;
        RECT 227.750 -811.770 228.130 -705.535 ;
        RECT 229.270 -817.985 229.650 -711.750 ;
        RECT 230.790 -811.770 231.170 -705.535 ;
        RECT 232.310 -817.985 232.690 -711.750 ;
        RECT 233.830 -811.770 234.210 -705.535 ;
        RECT 235.350 -817.985 235.730 -711.750 ;
        RECT 236.870 -811.770 237.250 -705.535 ;
        RECT 238.390 -817.985 238.770 -711.750 ;
        RECT 239.910 -811.770 240.290 -705.535 ;
        RECT 241.430 -817.985 241.810 -711.750 ;
        RECT 242.950 -811.770 243.330 -705.535 ;
        RECT 244.470 -817.985 244.850 -711.750 ;
        RECT 245.990 -811.770 246.370 -705.535 ;
        RECT 247.510 -817.985 247.890 -711.750 ;
        RECT 249.030 -811.770 249.410 -705.535 ;
        RECT 250.550 -817.985 250.930 -711.750 ;
        RECT 252.070 -811.770 252.450 -705.535 ;
        RECT 253.590 -817.985 253.970 -711.750 ;
        RECT 255.110 -811.770 255.490 -705.535 ;
        RECT 256.630 -817.985 257.010 -711.750 ;
        RECT 258.150 -811.770 258.530 -705.535 ;
        RECT 259.670 -817.985 260.050 -711.750 ;
        RECT 261.190 -811.770 261.570 -705.535 ;
        RECT 262.710 -817.985 263.090 -711.750 ;
        RECT 264.230 -811.770 264.610 -705.535 ;
        RECT 265.750 -817.985 266.130 -711.750 ;
        RECT 267.270 -811.770 267.650 -705.535 ;
        RECT 268.790 -817.985 269.170 -711.750 ;
        RECT 270.310 -811.770 270.690 -705.535 ;
        RECT 271.830 -817.985 272.210 -711.750 ;
        RECT 273.350 -811.770 273.730 -705.535 ;
        RECT 274.870 -817.985 275.250 -711.750 ;
        RECT 276.390 -811.770 276.770 -705.535 ;
        RECT 277.910 -817.985 278.290 -711.750 ;
        RECT 279.430 -811.770 279.810 -705.535 ;
        RECT 280.950 -817.985 281.330 -711.750 ;
        RECT 282.470 -811.770 282.850 -705.535 ;
        RECT 283.990 -817.985 284.370 -711.750 ;
        RECT 285.510 -811.770 285.890 -705.535 ;
        RECT 287.030 -817.985 287.410 -711.750 ;
        RECT 288.550 -811.770 288.930 -705.535 ;
        RECT 290.070 -817.985 290.450 -711.750 ;
        RECT 291.590 -811.770 291.970 -705.535 ;
        RECT 293.110 -817.985 293.490 -711.750 ;
        RECT 294.630 -811.770 295.010 -705.535 ;
        RECT 296.150 -817.985 296.530 -711.750 ;
        RECT 297.670 -811.770 298.050 -705.535 ;
        RECT 299.190 -817.985 299.570 -711.750 ;
        RECT 300.710 -811.770 301.090 -705.535 ;
        RECT 302.230 -817.985 302.610 -711.750 ;
        RECT 303.750 -811.770 304.130 -705.535 ;
        RECT 305.270 -817.985 305.650 -711.750 ;
        RECT 306.790 -811.770 307.170 -705.535 ;
        RECT 308.310 -817.985 308.690 -711.750 ;
        RECT 309.830 -811.770 310.210 -705.535 ;
        RECT 311.350 -817.985 311.730 -711.750 ;
        RECT 312.870 -811.770 313.250 -705.535 ;
        RECT 314.390 -817.985 314.770 -711.750 ;
        RECT 315.910 -811.770 316.290 -705.535 ;
        RECT 317.430 -817.985 317.810 -711.750 ;
        RECT 318.950 -811.770 319.330 -705.535 ;
        RECT 320.470 -817.985 320.850 -711.750 ;
        RECT 321.990 -811.770 322.370 -705.535 ;
        RECT 323.510 -817.985 323.890 -711.750 ;
        RECT 325.030 -811.770 325.410 -705.535 ;
        RECT 326.550 -817.985 326.930 -711.750 ;
        RECT 328.070 -811.770 328.450 -705.535 ;
        RECT 329.590 -817.985 329.970 -711.750 ;
        RECT 331.110 -811.770 331.490 -705.535 ;
        RECT 332.630 -817.985 333.010 -711.750 ;
        RECT 334.150 -811.770 334.530 -705.535 ;
        RECT 335.670 -817.985 336.050 -711.750 ;
        RECT 337.190 -811.770 337.570 -705.535 ;
        RECT 338.710 -817.985 339.090 -711.750 ;
        RECT 340.230 -811.770 340.610 -705.535 ;
        RECT 341.750 -817.985 342.130 -711.750 ;
        RECT 343.270 -811.770 343.650 -705.535 ;
        RECT 344.790 -817.985 345.170 -711.750 ;
        RECT 346.310 -811.770 346.690 -705.535 ;
        RECT 347.830 -817.985 348.210 -711.750 ;
        RECT 349.350 -811.770 349.730 -705.535 ;
        RECT 350.870 -817.985 351.250 -711.750 ;
        RECT 352.390 -811.770 352.770 -705.535 ;
        RECT 353.910 -817.985 354.290 -711.750 ;
        RECT 355.430 -811.770 355.810 -705.535 ;
        RECT 356.950 -817.985 357.330 -711.750 ;
        RECT 358.470 -811.770 358.850 -705.535 ;
        RECT 359.990 -817.985 360.370 -711.750 ;
        RECT 361.510 -811.770 361.890 -705.535 ;
        RECT 378.720 -811.760 379.890 -705.535 ;
        RECT 379.510 -811.770 379.890 -811.760 ;
        RECT 381.030 -817.985 381.410 -711.750 ;
        RECT 382.550 -811.770 382.930 -705.535 ;
        RECT 384.070 -817.985 384.450 -711.750 ;
        RECT 385.590 -811.770 385.970 -705.535 ;
        RECT 387.110 -817.985 387.490 -711.750 ;
        RECT 388.630 -811.770 389.010 -705.535 ;
        RECT 390.150 -817.985 390.530 -711.750 ;
        RECT 391.670 -811.770 392.050 -705.535 ;
        RECT 393.190 -817.985 393.570 -711.750 ;
        RECT 394.710 -811.770 395.090 -705.535 ;
        RECT 396.230 -817.985 396.610 -711.750 ;
        RECT 397.750 -811.770 398.130 -705.535 ;
        RECT 399.270 -817.985 399.650 -711.750 ;
        RECT 400.790 -811.770 401.170 -705.535 ;
        RECT 402.310 -817.985 402.690 -711.750 ;
        RECT 403.830 -811.770 404.210 -705.535 ;
        RECT 405.350 -817.985 405.730 -711.750 ;
        RECT 406.870 -811.770 407.250 -705.535 ;
        RECT 408.390 -817.985 408.770 -711.750 ;
        RECT 409.910 -811.770 410.290 -705.535 ;
        RECT 411.430 -817.985 411.810 -711.750 ;
        RECT 412.950 -811.770 413.330 -705.535 ;
        RECT 414.470 -817.985 414.850 -711.750 ;
        RECT 415.990 -811.770 416.370 -705.535 ;
        RECT 417.510 -817.985 417.890 -711.750 ;
        RECT 419.030 -811.770 419.410 -705.535 ;
        RECT 420.550 -817.985 420.930 -711.750 ;
        RECT 422.070 -811.770 422.450 -705.535 ;
        RECT 423.590 -817.985 423.970 -711.750 ;
        RECT 425.110 -811.770 425.490 -705.535 ;
        RECT 426.630 -817.985 427.010 -711.750 ;
        RECT 428.150 -811.770 428.530 -705.535 ;
        RECT 429.670 -817.985 430.050 -711.750 ;
        RECT 431.190 -811.770 431.570 -705.535 ;
        RECT 432.710 -817.985 433.090 -711.750 ;
        RECT 434.230 -811.770 434.610 -705.535 ;
        RECT 435.750 -817.985 436.130 -711.750 ;
        RECT 437.270 -811.770 437.650 -705.535 ;
        RECT 438.790 -817.985 439.170 -711.750 ;
        RECT 440.310 -811.770 440.690 -705.535 ;
        RECT 441.830 -817.985 442.210 -711.750 ;
        RECT 443.350 -811.770 443.730 -705.535 ;
        RECT 444.870 -817.985 445.250 -711.750 ;
        RECT 446.390 -811.770 446.770 -705.535 ;
        RECT 447.910 -817.985 448.290 -711.750 ;
        RECT 449.430 -811.770 449.810 -705.535 ;
        RECT 450.950 -817.985 451.330 -711.750 ;
        RECT 452.470 -811.770 452.850 -705.535 ;
        RECT 453.990 -817.985 454.370 -711.750 ;
        RECT 455.510 -811.770 455.890 -705.535 ;
        RECT 457.030 -817.985 457.410 -711.750 ;
        RECT 458.550 -811.770 458.930 -705.535 ;
        RECT 460.070 -817.985 460.450 -711.750 ;
        RECT 461.590 -811.770 461.970 -705.535 ;
        RECT 463.110 -817.985 463.490 -711.750 ;
        RECT 464.630 -811.770 465.010 -705.535 ;
        RECT 466.150 -817.985 466.530 -711.750 ;
        RECT 467.670 -811.770 468.050 -705.535 ;
        RECT 469.190 -817.985 469.570 -711.750 ;
        RECT 470.710 -811.770 471.090 -705.535 ;
        RECT 472.230 -817.985 472.610 -711.750 ;
        RECT 473.750 -811.770 474.130 -705.535 ;
        RECT 475.270 -817.985 475.650 -711.750 ;
        RECT 476.790 -811.770 477.170 -705.535 ;
        RECT 478.310 -817.985 478.690 -711.750 ;
        RECT 479.830 -811.770 480.210 -705.535 ;
        RECT 481.350 -817.985 481.730 -711.750 ;
        RECT 482.870 -811.770 483.250 -705.535 ;
        RECT 484.390 -817.985 484.770 -711.750 ;
        RECT 485.910 -811.770 486.290 -705.535 ;
        RECT 487.430 -817.985 487.810 -711.750 ;
        RECT 488.950 -811.770 489.330 -705.535 ;
        RECT 490.470 -817.985 490.850 -711.750 ;
        RECT 491.990 -811.770 492.370 -705.535 ;
        RECT 493.510 -817.985 493.890 -711.750 ;
        RECT 495.030 -811.770 495.410 -705.535 ;
        RECT 496.550 -817.985 496.930 -711.750 ;
        RECT 498.070 -811.770 498.450 -705.535 ;
        RECT 499.590 -817.985 499.970 -711.750 ;
        RECT 501.110 -811.770 501.490 -705.535 ;
        RECT 502.630 -817.985 503.010 -711.750 ;
        RECT 504.150 -811.770 504.530 -705.535 ;
        RECT 505.670 -817.985 506.050 -711.750 ;
        RECT 507.190 -811.770 507.570 -705.535 ;
        RECT 508.710 -817.985 509.090 -711.750 ;
        RECT 510.230 -811.770 510.610 -705.535 ;
        RECT 511.750 -817.985 512.130 -711.750 ;
        RECT 513.270 -811.770 513.650 -705.535 ;
        RECT 514.790 -817.985 515.170 -711.750 ;
        RECT 516.310 -811.770 516.690 -705.535 ;
        RECT 517.830 -817.985 518.210 -711.750 ;
        RECT 519.350 -811.770 519.730 -705.535 ;
        RECT 520.870 -817.985 521.250 -711.750 ;
        RECT 522.390 -811.770 522.770 -705.535 ;
        RECT 523.910 -817.985 524.290 -711.750 ;
        RECT 525.430 -811.770 525.810 -705.535 ;
        RECT 526.950 -817.985 527.330 -711.750 ;
        RECT 528.470 -811.770 528.850 -705.535 ;
        RECT 529.990 -817.985 530.370 -711.750 ;
        RECT 531.510 -811.770 531.890 -705.535 ;
        RECT 548.720 -811.760 549.890 -705.535 ;
        RECT 549.510 -811.770 549.890 -811.760 ;
        RECT 551.030 -817.985 551.410 -711.750 ;
        RECT 552.550 -811.770 552.930 -705.535 ;
        RECT 554.070 -817.985 554.450 -711.750 ;
        RECT 555.590 -811.770 555.970 -705.535 ;
        RECT 557.110 -817.985 557.490 -711.750 ;
        RECT 558.630 -811.770 559.010 -705.535 ;
        RECT 560.150 -817.985 560.530 -711.750 ;
        RECT 561.670 -811.770 562.050 -705.535 ;
        RECT 563.190 -817.985 563.570 -711.750 ;
        RECT 564.710 -811.770 565.090 -705.535 ;
        RECT 566.230 -817.985 566.610 -711.750 ;
        RECT 567.750 -811.770 568.130 -705.535 ;
        RECT 569.270 -817.985 569.650 -711.750 ;
        RECT 570.790 -811.770 571.170 -705.535 ;
        RECT 572.310 -817.985 572.690 -711.750 ;
        RECT 573.830 -811.770 574.210 -705.535 ;
        RECT 575.350 -817.985 575.730 -711.750 ;
        RECT 576.870 -811.770 577.250 -705.535 ;
        RECT 578.390 -817.985 578.770 -711.750 ;
        RECT 579.910 -811.770 580.290 -705.535 ;
        RECT 581.430 -817.985 581.810 -711.750 ;
        RECT 582.950 -811.770 583.330 -705.535 ;
        RECT 584.470 -817.985 584.850 -711.750 ;
        RECT 585.990 -811.770 586.370 -705.535 ;
        RECT 587.510 -817.985 587.890 -711.750 ;
        RECT 589.030 -811.770 589.410 -705.535 ;
        RECT 590.550 -817.985 590.930 -711.750 ;
        RECT 592.070 -811.770 592.450 -705.535 ;
        RECT 593.590 -817.985 593.970 -711.750 ;
        RECT 595.110 -811.770 595.490 -705.535 ;
        RECT 596.630 -817.985 597.010 -711.750 ;
        RECT 598.150 -811.770 598.530 -705.535 ;
        RECT 599.670 -817.985 600.050 -711.750 ;
        RECT 601.190 -811.770 601.570 -705.535 ;
        RECT 602.710 -817.985 603.090 -711.750 ;
        RECT 604.230 -811.770 604.610 -705.535 ;
        RECT 605.750 -817.985 606.130 -711.750 ;
        RECT 607.270 -811.770 607.650 -705.535 ;
        RECT 608.790 -817.985 609.170 -711.750 ;
        RECT 610.310 -811.770 610.690 -705.535 ;
        RECT 611.830 -817.985 612.210 -711.750 ;
        RECT 613.350 -811.770 613.730 -705.535 ;
        RECT 614.870 -817.985 615.250 -711.750 ;
        RECT 616.390 -811.770 616.770 -705.535 ;
        RECT 617.910 -817.985 618.290 -711.750 ;
        RECT 619.430 -811.770 619.810 -705.535 ;
        RECT 620.950 -817.985 621.330 -711.750 ;
        RECT 622.470 -811.770 622.850 -705.535 ;
        RECT 623.990 -817.985 624.370 -711.750 ;
        RECT 625.510 -811.770 625.890 -705.535 ;
        RECT 627.030 -817.985 627.410 -711.750 ;
        RECT 628.550 -811.770 628.930 -705.535 ;
        RECT 630.070 -817.985 630.450 -711.750 ;
        RECT 631.590 -811.770 631.970 -705.535 ;
        RECT 633.110 -817.985 633.490 -711.750 ;
        RECT 634.630 -811.770 635.010 -705.535 ;
        RECT 636.150 -817.985 636.530 -711.750 ;
        RECT 637.670 -811.770 638.050 -705.535 ;
        RECT 639.190 -817.985 639.570 -711.750 ;
        RECT 640.710 -811.770 641.090 -705.535 ;
        RECT 642.230 -817.985 642.610 -711.750 ;
        RECT 643.750 -811.770 644.130 -705.535 ;
        RECT 645.270 -817.985 645.650 -711.750 ;
        RECT 646.790 -811.770 647.170 -705.535 ;
        RECT 648.310 -817.985 648.690 -711.750 ;
        RECT 649.830 -811.770 650.210 -705.535 ;
        RECT 651.350 -817.985 651.730 -711.750 ;
        RECT 652.870 -811.770 653.250 -705.535 ;
        RECT 654.390 -817.985 654.770 -711.750 ;
        RECT 655.910 -811.770 656.290 -705.535 ;
        RECT 657.430 -817.985 657.810 -711.750 ;
        RECT 658.950 -811.770 659.330 -705.535 ;
        RECT 660.470 -817.985 660.850 -711.750 ;
        RECT 661.990 -811.770 662.370 -705.535 ;
        RECT 663.510 -817.985 663.890 -711.750 ;
        RECT 665.030 -811.770 665.410 -705.535 ;
        RECT 666.550 -817.985 666.930 -711.750 ;
        RECT 668.070 -811.770 668.450 -705.535 ;
        RECT 669.590 -817.985 669.970 -711.750 ;
        RECT 671.110 -811.770 671.490 -705.535 ;
        RECT 672.630 -817.985 673.010 -711.750 ;
        RECT 674.150 -811.770 674.530 -705.535 ;
        RECT 675.670 -817.985 676.050 -711.750 ;
        RECT 677.190 -811.770 677.570 -705.535 ;
        RECT 678.710 -817.985 679.090 -711.750 ;
        RECT 680.230 -811.770 680.610 -705.535 ;
        RECT 681.750 -817.985 682.130 -711.750 ;
        RECT 683.270 -811.770 683.650 -705.535 ;
        RECT 684.790 -817.985 685.170 -711.750 ;
        RECT 686.310 -811.770 686.690 -705.535 ;
        RECT 687.830 -817.985 688.210 -711.750 ;
        RECT 689.350 -811.770 689.730 -705.535 ;
        RECT 690.870 -817.985 691.250 -711.750 ;
        RECT 692.390 -811.770 692.770 -705.535 ;
        RECT 693.910 -817.985 694.290 -711.750 ;
        RECT 695.430 -811.770 695.810 -705.535 ;
        RECT 696.950 -817.985 697.330 -711.750 ;
        RECT 698.470 -811.770 698.850 -705.535 ;
        RECT 699.990 -817.985 700.370 -711.750 ;
        RECT 701.510 -811.770 701.890 -705.535 ;
        RECT 718.720 -811.760 719.890 -705.535 ;
        RECT 719.510 -811.770 719.890 -811.760 ;
        RECT 721.030 -817.985 721.410 -711.750 ;
        RECT 722.550 -811.770 722.930 -705.535 ;
        RECT 724.070 -817.985 724.450 -711.750 ;
        RECT 725.590 -811.770 725.970 -705.535 ;
        RECT 727.110 -817.985 727.490 -711.750 ;
        RECT 728.630 -811.770 729.010 -705.535 ;
        RECT 730.150 -817.985 730.530 -711.750 ;
        RECT 731.670 -811.770 732.050 -705.535 ;
        RECT 733.190 -817.985 733.570 -711.750 ;
        RECT 734.710 -811.770 735.090 -705.535 ;
        RECT 736.230 -817.985 736.610 -711.750 ;
        RECT 737.750 -811.770 738.130 -705.535 ;
        RECT 739.270 -817.985 739.650 -711.750 ;
        RECT 740.790 -811.770 741.170 -705.535 ;
        RECT 742.310 -817.985 742.690 -711.750 ;
        RECT 743.830 -811.770 744.210 -705.535 ;
        RECT 745.350 -817.985 745.730 -711.750 ;
        RECT 746.870 -811.770 747.250 -705.535 ;
        RECT 748.390 -817.985 748.770 -711.750 ;
        RECT 749.910 -811.770 750.290 -705.535 ;
        RECT 751.430 -817.985 751.810 -711.750 ;
        RECT 752.950 -811.770 753.330 -705.535 ;
        RECT 754.470 -817.985 754.850 -711.750 ;
        RECT 755.990 -811.770 756.370 -705.535 ;
        RECT 757.510 -817.985 757.890 -711.750 ;
        RECT 759.030 -811.770 759.410 -705.535 ;
        RECT 760.550 -817.985 760.930 -711.750 ;
        RECT 762.070 -811.770 762.450 -705.535 ;
        RECT 763.590 -817.985 763.970 -711.750 ;
        RECT 765.110 -811.770 765.490 -705.535 ;
        RECT 766.630 -817.985 767.010 -711.750 ;
        RECT 768.150 -811.770 768.530 -705.535 ;
        RECT 769.670 -817.985 770.050 -711.750 ;
        RECT 771.190 -811.770 771.570 -705.535 ;
        RECT 772.710 -817.985 773.090 -711.750 ;
        RECT 774.230 -811.770 774.610 -705.535 ;
        RECT 775.750 -817.985 776.130 -711.750 ;
        RECT 777.270 -811.770 777.650 -705.535 ;
        RECT 778.790 -817.985 779.170 -711.750 ;
        RECT 780.310 -811.770 780.690 -705.535 ;
        RECT 781.830 -817.985 782.210 -711.750 ;
        RECT 783.350 -811.770 783.730 -705.535 ;
        RECT 784.870 -817.985 785.250 -711.750 ;
        RECT 786.390 -811.770 786.770 -705.535 ;
        RECT 787.910 -817.985 788.290 -711.750 ;
        RECT 789.430 -811.770 789.810 -705.535 ;
        RECT 790.950 -817.985 791.330 -711.750 ;
        RECT 792.470 -811.770 792.850 -705.535 ;
        RECT 793.990 -817.985 794.370 -711.750 ;
        RECT 795.510 -811.770 795.890 -705.535 ;
        RECT 797.030 -817.985 797.410 -711.750 ;
        RECT 798.550 -811.770 798.930 -705.535 ;
        RECT 800.070 -817.985 800.450 -711.750 ;
        RECT 801.590 -811.770 801.970 -705.535 ;
        RECT 803.110 -817.985 803.490 -711.750 ;
        RECT 804.630 -811.770 805.010 -705.535 ;
        RECT 806.150 -817.985 806.530 -711.750 ;
        RECT 807.670 -811.770 808.050 -705.535 ;
        RECT 809.190 -817.985 809.570 -711.750 ;
        RECT 810.710 -811.770 811.090 -705.535 ;
        RECT 812.230 -817.985 812.610 -711.750 ;
        RECT 813.750 -811.770 814.130 -705.535 ;
        RECT 815.270 -817.985 815.650 -711.750 ;
        RECT 816.790 -811.770 817.170 -705.535 ;
        RECT 818.310 -817.985 818.690 -711.750 ;
        RECT 819.830 -811.770 820.210 -705.535 ;
        RECT 821.350 -817.985 821.730 -711.750 ;
        RECT 822.870 -811.770 823.250 -705.535 ;
        RECT 824.390 -817.985 824.770 -711.750 ;
        RECT 825.910 -811.770 826.290 -705.535 ;
        RECT 827.430 -817.985 827.810 -711.750 ;
        RECT 828.950 -811.770 829.330 -705.535 ;
        RECT 830.470 -817.985 830.850 -711.750 ;
        RECT 831.990 -811.770 832.370 -705.535 ;
        RECT 833.510 -817.985 833.890 -711.750 ;
        RECT 835.030 -811.770 835.410 -705.535 ;
        RECT 836.550 -817.985 836.930 -711.750 ;
        RECT 838.070 -811.770 838.450 -705.535 ;
        RECT 839.590 -817.985 839.970 -711.750 ;
        RECT 841.110 -811.770 841.490 -705.535 ;
        RECT 842.630 -817.985 843.010 -711.750 ;
        RECT 844.150 -811.770 844.530 -705.535 ;
        RECT 845.670 -817.985 846.050 -711.750 ;
        RECT 847.190 -811.770 847.570 -705.535 ;
        RECT 848.710 -817.985 849.090 -711.750 ;
        RECT 850.230 -811.770 850.610 -705.535 ;
        RECT 851.750 -817.985 852.130 -711.750 ;
        RECT 853.270 -811.770 853.650 -705.535 ;
        RECT 854.790 -817.985 855.170 -711.750 ;
        RECT 856.310 -811.770 856.690 -705.535 ;
        RECT 857.830 -817.985 858.210 -711.750 ;
        RECT 859.350 -811.770 859.730 -705.535 ;
        RECT 860.870 -817.985 861.250 -711.750 ;
        RECT 862.390 -811.770 862.770 -705.535 ;
        RECT 863.910 -817.985 864.290 -711.750 ;
        RECT 865.430 -811.770 865.810 -705.535 ;
        RECT 866.950 -817.985 867.330 -711.750 ;
        RECT 868.470 -811.770 868.850 -705.535 ;
        RECT 869.990 -817.985 870.370 -711.750 ;
        RECT 871.510 -811.770 871.890 -705.535 ;
        RECT -298.970 -843.445 873.410 -817.985 ;
        RECT 408.135 -882.355 892.360 -856.395 ;
      LAYER Metal2 ;
        RECT -527.150 1.895 -91.505 25.205 ;
        RECT -527.150 -686.875 -481.345 1.895 ;
        RECT -83.605 -14.790 591.125 -10.530 ;
        RECT 604.575 -14.790 623.570 15.700 ;
        RECT -83.605 -22.360 627.005 -14.790 ;
        RECT -83.605 -24.020 591.125 -22.360 ;
        RECT 604.575 -23.340 623.570 -22.360 ;
        RECT -83.605 -40.875 -17.185 -24.020 ;
        RECT -71.065 -55.045 -25.115 -40.875 ;
        RECT -435.970 -724.945 -358.995 -115.075 ;
        RECT -253.840 -542.990 -210.000 -401.350 ;
        RECT -82.045 -669.335 -14.465 -55.045 ;
        RECT 35.970 -387.375 91.820 -35.970 ;
        RECT 171.035 -669.335 239.765 -37.425 ;
        RECT 892.305 -59.890 906.660 53.180 ;
        RECT 865.660 -67.230 906.660 -59.890 ;
        RECT 398.980 -416.210 446.270 -115.075 ;
        RECT 542.480 -270.595 585.980 -115.075 ;
        RECT 405.305 -878.275 448.700 -680.075 ;
        RECT 713.300 -843.335 774.745 -79.430 ;
        RECT 865.660 -93.085 873.700 -67.230 ;
        RECT 943.025 -860.320 962.020 34.935 ;
        RECT 812.035 -877.875 962.020 -860.320 ;
        RECT 943.025 -880.770 962.020 -877.875 ;
      LAYER Metal3 ;
        RECT 893.970 44.330 903.255 85.505 ;
        RECT 944.990 28.415 960.480 43.190 ;
        RECT 606.540 9.180 622.030 23.955 ;
      LAYER Metal4 ;
        RECT 565.125 158.715 671.125 161.715 ;
        RECT 565.125 33.715 568.125 158.715 ;
        RECT 668.125 33.715 671.125 158.715 ;
        RECT 565.125 24.715 671.125 33.715 ;
        RECT 674.125 158.715 780.125 161.715 ;
        RECT 674.125 33.715 677.125 158.715 ;
        RECT 777.125 33.715 780.125 158.715 ;
        RECT 674.125 24.715 780.125 33.715 ;
        RECT 783.125 158.715 889.125 161.715 ;
        RECT 783.125 33.715 786.125 158.715 ;
        RECT 886.125 33.715 889.125 158.715 ;
        RECT 929.525 148.580 1066.525 151.580 ;
        RECT 893.970 78.935 902.465 101.275 ;
        RECT 929.525 48.580 932.525 148.580 ;
        RECT 1057.525 48.580 1066.525 148.580 ;
        RECT 929.525 45.580 1066.525 48.580 ;
        RECT 946.180 36.895 959.215 45.580 ;
        RECT 783.125 24.715 889.125 33.715 ;
        RECT 607.730 17.660 620.765 24.715 ;
      LAYER Metal5 ;
        RECT 570.125 98.865 666.125 156.715 ;
        RECT 679.125 98.865 775.125 156.715 ;
        RECT 788.125 98.865 884.125 156.715 ;
        RECT 934.525 100.140 1055.525 146.580 ;
        RECT 890.290 98.865 1055.525 100.140 ;
        RECT 563.625 93.565 1055.525 98.865 ;
        RECT 570.125 35.715 666.125 93.565 ;
        RECT 679.125 35.715 775.125 93.565 ;
        RECT 788.125 35.715 884.125 93.565 ;
        RECT 934.525 50.580 1055.525 93.565 ;
        RECT 1062.775 47.005 1064.975 150.155 ;
        RECT 563.625 24.715 890.625 30.015 ;
  END
END OTA_2stage
END LIBRARY

