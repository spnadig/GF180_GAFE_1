VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OTA_2stage_macro
  CLASS BLOCK ;
  FOREIGN OTA_2stage_macro ;
  ORIGIN 0.000 0.000 ;
  SIZE 1804.180 BY 1218.995 ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 106.565 349.955 187.040 409.555 ;
    END
  END vss
  PIN vin2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 106.565 275.300 152.710 334.780 ;
    END
  END vin2
  PIN vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 106.565 198.065 125.530 257.060 ;
    END
  END vout
  PIN vin1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 106.565 426.605 153.105 483.565 ;
    END
  END vin1
  PIN vp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 106.565 503.490 128.500 557.990 ;
    END
  END vp
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 45.090 628.080 109.565 720.005 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 10.530 720.305 1782.660 1153.455 ;
        RECT 10.530 627.780 44.790 720.305 ;
        RECT 109.865 627.780 1782.660 720.305 ;
        RECT 10.530 558.290 1782.660 627.780 ;
        RECT 10.530 503.190 106.265 558.290 ;
        RECT 128.800 503.190 1782.660 558.290 ;
        RECT 10.530 483.865 1782.660 503.190 ;
        RECT 10.530 426.305 106.265 483.865 ;
        RECT 153.405 426.305 1782.660 483.865 ;
        RECT 10.530 409.855 1782.660 426.305 ;
        RECT 10.530 349.655 106.265 409.855 ;
        RECT 187.340 349.655 1782.660 409.855 ;
        RECT 10.530 335.080 1782.660 349.655 ;
        RECT 10.530 275.000 106.265 335.080 ;
        RECT 153.010 275.000 1782.660 335.080 ;
        RECT 10.530 257.360 1782.660 275.000 ;
        RECT 10.530 197.765 106.265 257.360 ;
        RECT 125.830 197.765 1782.660 257.360 ;
        RECT 10.530 3.905 1782.660 197.765 ;
      LAYER Metal2 ;
        RECT 10.690 32.950 1695.285 1218.995 ;
      LAYER Metal3 ;
        RECT 10.690 112.505 1732.275 1218.995 ;
      LAYER Metal4 ;
        RECT 10.690 112.505 1799.790 1218.995 ;
      LAYER Metal5 ;
        RECT 10.690 112.505 1798.240 1218.995 ;
  END
END OTA_2stage_macro
END LIBRARY

