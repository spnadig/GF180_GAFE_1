VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OTA_2stage
  CLASS BLOCK ;
  FOREIGN OTA_2stage ;
  ORIGIN 0.000 0.000 ;
  SIZE 1950.000 BY 1250.000 ;
  PIN vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1679.325 851.115 1896.265 880.615 ;
    END
  END vout
  PIN vin1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.485 765.035 145.415 778.985 ;
    END
  END vin1
  PIN vp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 619.445 1059.895 659.415 1165.190 ;
    END
  END vp
  PIN vin2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1706.630 465.030 1889.190 495.195 ;
    END
  END vin2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 205.205 73.135 1185.550 99.095 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 776.875 1008.880 903.255 1116.735 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 8.485 1165.490 1744.395 1168.515 ;
        RECT 8.485 1059.595 619.145 1165.490 ;
        RECT 659.715 1117.035 1744.395 1165.490 ;
        RECT 659.715 1059.595 776.575 1117.035 ;
        RECT 8.485 1008.580 776.575 1059.595 ;
        RECT 903.555 1008.580 1744.395 1117.035 ;
        RECT 8.485 880.915 1744.395 1008.580 ;
        RECT 8.485 850.815 1679.025 880.915 ;
        RECT 8.485 779.285 1744.395 850.815 ;
        RECT 8.485 778.985 127.030 779.285 ;
        RECT 145.715 764.735 1744.395 779.285 ;
        RECT 8.485 495.495 1744.395 764.735 ;
        RECT 8.485 464.730 1706.330 495.495 ;
        RECT 8.485 99.395 1744.395 464.730 ;
        RECT 8.485 72.835 204.905 99.395 ;
        RECT 1185.850 72.835 1744.395 99.395 ;
        RECT 8.485 10.950 1744.395 72.835 ;
      LAYER Metal2 ;
        RECT 250.265 63.955 1739.435 1011.080 ;
      LAYER Metal3 ;
        RECT 89.615 143.510 1776.425 1107.145 ;
      LAYER Metal4 ;
        RECT 89.615 143.510 1843.940 1117.205 ;
      LAYER Metal5 ;
        RECT 105.315 143.510 1842.390 1112.205 ;
  END
END OTA_2stage
END LIBRARY

