* SPICE3 file created from top.ext - technology: gf180mcuC


.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VNW VPW
X0 Z a_36_113# VDD VNW pfet_06v0 ad=0.5368p pd=3.32u as=0.803p ps=3.84u w=1.22u l=0.5u
X1 Z a_36_113# VSS VPW nfet_06v0 ad=0.2178p pd=1.87u as=0.306p ps=2.39u w=0.495u l=0.6u
X2 VSS I a_36_113# VPW nfet_06v0 ad=0p pd=0u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3 VDD I a_36_113# VNW pfet_06v0 ad=0p pd=0u as=0.462p ps=2.98u w=1.05u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VNW VPW
X0 a_244_159# A1 a_36_159# VPW nfet_06v0 ad=0.1168p pd=1.37u as=0.1606p ps=1.61u w=0.365u l=0.6u
X1 a_36_159# A1 VDD VNW pfet_06v0 ad=0.312p pd=2.24u as=1.0755p ps=6.19u w=0.6u l=0.5u
X2 VDD A2 a_36_159# VNW pfet_06v0 ad=0p pd=0u as=0p ps=0u w=0.6u l=0.5u
X3 Z a_36_159# VDD VNW pfet_06v0 ad=0.5346p pd=3.31u as=0p ps=0u w=1.215u l=0.5u
X4 Z a_36_159# VSS VPW nfet_06v0 ad=0.3586p pd=2.51u as=0.4681p ps=3.11u w=0.815u l=0.6u
X5 VSS A2 a_244_159# VPW nfet_06v0 ad=0p pd=0u as=0p ps=0u w=0.365u l=0.6u
.ends

.subckt TopLevel_oscillator Y VP GND
X0 a_1067_4019# a_n3996_4046# VP VP pfet_03v3 ad=0.22p pd=1.88u as=0.66p ps=5.64u w=0.5u l=5u
X1 a_1067_4019# a_n3996_4046# GND GND nfet_03v3 ad=0.22p pd=1.88u as=0.66p ps=5.64u w=0.5u l=5u
X2 a_n3996_4046# Y GND GND nfet_03v3 ad=0.22p pd=1.88u as=0p ps=0u w=0.5u l=5u
X3 Y a_1067_4019# VP VP pfet_03v3 ad=0.22p pd=1.88u as=0p ps=0u w=0.5u l=5u
X4 Y a_1067_4019# GND GND nfet_03v3 ad=0.22p pd=1.88u as=0p ps=0u w=0.5u l=5u
X5 a_n3996_4046# Y VP VP pfet_03v3 ad=0.22p pd=1.88u as=0p ps=0u w=0.5u l=5u
C0 Y GND 30.75fF
C1 VP GND 5.07fF
C2 a_1067_4019# GND 11.97fF
C3 a_n3996_4046# GND 12.06fF
.ends

.subckt top VDD osc_out VSS osc_en
Xinput1 VSS net1 osc_en VDD input1/VNW VSUBS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0_ VDD VSS osc_out net1 osc_sig _0_/VNW VSUBS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xosc0 osc_sig osc0/VP VSUBS TopLevel_oscillator
C0 VDD VSS 61.32fF
C1 osc_out VSS 3.54fF
C2 net1 VSS 4.22fF
C3 VSS VSUBS 188.76fF
C4 VDD VSUBS 177.25fF
C5 osc_sig VSUBS 31.49fF
C6 osc0/VP VSUBS 5.07fF
C11 _0_/VNW VSUBS 3.40fF
.ends

