VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO TopLevel_oscillator_macro
  CLASS BLOCK ;
  FOREIGN TopLevel_oscillator_macro ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 570.000 ;
  PIN VP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 309.060 478.920 309.070 478.930 ;
    END
  END VP
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 388.440 493.585 388.450 493.595 ;
    END
  END GND
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 223.185 500.770 223.195 500.780 ;
    END
  END Y
  PIN ASIG5V
    PORT
      LAYER Metal5 ;
        RECT -112.600 123.490 -112.590 123.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -27.600 123.490 -27.590 123.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 14.480 123.085 89.480 123.515 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 99.480 123.085 174.480 123.515 ;
    END
  END ASIG5V
  PIN CLK_EN
    PORT
      LAYER Metal2 ;
        RECT 46.780 501.020 46.790 501.030 ;
    END
  END CLK_EN
  PIN AND_OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 121.940 491.525 123.640 491.955 ;
    END
  END AND_OUT
  OBS
      LAYER Metal1 ;
        RECT 14.320 78.310 429.640 429.980 ;
      LAYER Metal2 ;
        RECT 14.480 501.330 429.480 529.365 ;
        RECT 14.480 500.720 46.480 501.330 ;
        RECT 47.090 500.720 429.480 501.330 ;
        RECT 14.480 492.255 429.480 500.720 ;
        RECT 14.480 491.225 121.640 492.255 ;
        RECT 123.940 491.225 429.480 492.255 ;
        RECT 14.480 12.770 429.480 491.225 ;
      LAYER Metal3 ;
        RECT 14.480 12.770 429.480 529.365 ;
      LAYER Metal4 ;
        RECT 14.480 12.770 429.480 529.365 ;
      LAYER Metal5 ;
        RECT 14.480 124.015 429.480 529.365 ;
        RECT 89.980 122.585 98.980 124.015 ;
        RECT 174.980 122.585 429.480 124.015 ;
        RECT 14.480 12.770 429.480 122.585 ;
  END
END TopLevel_oscillator_macro
END LIBRARY

