* Extracted by KLayout with GF180 LVS runset on : 07/02/2023 03:42

.SUBCKT TopLevel_oscillator GND
X$1 \$4 \$2 \$5 \$1 GND inverter
X$2 \$5 \$2 \$3 \$1 GND inverter
X$3 \$3 \$2 \$4 \$1 GND inverter
.ENDS TopLevel_oscillator

.SUBCKT inverter A GND Y VP GND$1
M$1 GND A Y GND$1 nfet_03v3 L=5U W=0.5U AS=0.22P AD=0.22P PS=1.88U PD=1.88U
M$2 VP A Y VP pfet_03v3 L=5U W=0.5U AS=0.22P AD=0.22P PS=1.88U PD=1.88U
.ENDS inverter
