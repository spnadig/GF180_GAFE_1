VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OTA_2stage
  CLASS BLOCK ;
  FOREIGN OTA_2stage ;
  ORIGIN 0.000 0.000 ;
  SIZE 2046.900 BY 1307.330 ;
  PIN vin1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 162.150 808.940 187.920 822.890 ;
    END
  END vin1
  PIN vp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 661.950 1103.800 701.920 1135.355 ;
    END
  END vp
  PIN vin2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1737.550 521.860 1762.945 539.095 ;
    END
  END vin2
  PIN vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1690.540 895.020 1710.630 924.520 ;
    END
  END vout
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 247.710 117.035 1228.055 142.995 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 819.380 1052.785 945.760 1160.640 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 162.150 1135.655 819.080 1160.640 ;
        RECT 162.150 1103.500 661.650 1135.655 ;
        RECT 702.220 1103.500 819.080 1135.655 ;
        RECT 162.150 1052.485 819.080 1103.500 ;
        RECT 946.060 1052.485 1762.945 1160.640 ;
        RECT 162.150 924.820 1762.945 1052.485 ;
        RECT 162.150 894.720 1690.240 924.820 ;
        RECT 1710.930 894.720 1762.945 924.820 ;
        RECT 162.150 823.190 1762.945 894.720 ;
        RECT 188.220 808.640 1762.945 823.190 ;
        RECT 162.150 539.395 1762.945 808.640 ;
        RECT 162.150 521.560 1737.250 539.395 ;
        RECT 162.150 143.295 1762.945 521.560 ;
        RECT 162.150 117.035 247.410 143.295 ;
        RECT 1228.355 117.035 1762.945 143.295 ;
      LAYER Metal2 ;
        RECT 292.770 118.620 1781.940 1052.575 ;
      LAYER Metal3 ;
        RECT 1426.460 1008.575 1780.400 1084.900 ;
      LAYER Metal4 ;
        RECT 1385.045 1017.055 1886.445 1161.110 ;
      LAYER Metal5 ;
        RECT 1383.545 1024.110 1884.895 1156.110 ;
  END
END OTA_2stage
END LIBRARY

