magic
tech gf180mcuC
magscale 1 10
timestamp 1676577649
<< error_p >>
rect -66 0 -64 20000
rect 0 0 2 20000
<< nmos >>
rect 88 0 288 20000
rect 392 0 592 20000
rect 696 0 896 20000
rect 1000 0 1200 20000
rect 1304 0 1504 20000
rect 1608 0 1808 20000
rect 1912 0 2112 20000
rect 2216 0 2416 20000
rect 2520 0 2720 20000
rect 2824 0 3024 20000
rect 3128 0 3328 20000
rect 3432 0 3632 20000
rect 3736 0 3936 20000
rect 4040 0 4240 20000
rect 4344 0 4544 20000
rect 4648 0 4848 20000
rect 4952 0 5152 20000
rect 5256 0 5456 20000
rect 5560 0 5760 20000
rect 5864 0 6064 20000
rect 6168 0 6368 20000
rect 6472 0 6672 20000
rect 6776 0 6976 20000
rect 7080 0 7280 20000
rect 7384 0 7584 20000
rect 7688 0 7888 20000
rect 7992 0 8192 20000
rect 8296 0 8496 20000
rect 8600 0 8800 20000
rect 8904 0 9104 20000
rect 9208 0 9408 20000
rect 9512 0 9712 20000
rect 9816 0 10016 20000
rect 10120 0 10320 20000
rect 10424 0 10624 20000
rect 10728 0 10928 20000
rect 11032 0 11232 20000
rect 11336 0 11536 20000
rect 11640 0 11840 20000
rect 11944 0 12144 20000
rect 12248 0 12448 20000
rect 12552 0 12752 20000
rect 12856 0 13056 20000
rect 13160 0 13360 20000
rect 13464 0 13664 20000
rect 13768 0 13968 20000
rect 14072 0 14272 20000
rect 14376 0 14576 20000
rect 14680 0 14880 20000
rect 14984 0 15184 20000
rect 15288 0 15488 20000
rect 15592 0 15792 20000
rect 15896 0 16096 20000
rect 16200 0 16400 20000
rect 16504 0 16704 20000
rect 16808 0 17008 20000
rect 17112 0 17312 20000
rect 17416 0 17616 20000
rect 17720 0 17920 20000
rect 18024 0 18224 20000
rect 18328 0 18528 20000
rect 18632 0 18832 20000
rect 18936 0 19136 20000
rect 19240 0 19440 20000
rect 19544 0 19744 20000
rect 19848 0 20048 20000
rect 20152 0 20352 20000
rect 20456 0 20656 20000
rect 20760 0 20960 20000
rect 21064 0 21264 20000
rect 21368 0 21568 20000
rect 21672 0 21872 20000
rect 21976 0 22176 20000
rect 22280 0 22480 20000
rect 22584 0 22784 20000
rect 22888 0 23088 20000
rect 23192 0 23392 20000
rect 23496 0 23696 20000
rect 23800 0 24000 20000
rect 24104 0 24304 20000
rect 24408 0 24608 20000
rect 24712 0 24912 20000
rect 25016 0 25216 20000
rect 25320 0 25520 20000
rect 25624 0 25824 20000
rect 25928 0 26128 20000
rect 26232 0 26432 20000
rect 26536 0 26736 20000
rect 26840 0 27040 20000
rect 27144 0 27344 20000
rect 27448 0 27648 20000
rect 27752 0 27952 20000
rect 28056 0 28256 20000
rect 28360 0 28560 20000
rect 28664 0 28864 20000
rect 28968 0 29168 20000
rect 29272 0 29472 20000
rect 29576 0 29776 20000
rect 29880 0 30080 20000
rect 30184 0 30384 20000
<< ndiff >>
rect 0 19973 88 20000
rect 0 27 13 19973
rect 59 27 88 19973
rect 0 0 88 27
rect 288 19973 392 20000
rect 288 27 317 19973
rect 363 27 392 19973
rect 288 0 392 27
rect 592 19973 696 20000
rect 592 27 621 19973
rect 667 27 696 19973
rect 592 0 696 27
rect 896 19973 1000 20000
rect 896 27 925 19973
rect 971 27 1000 19973
rect 896 0 1000 27
rect 1200 19973 1304 20000
rect 1200 27 1229 19973
rect 1275 27 1304 19973
rect 1200 0 1304 27
rect 1504 19973 1608 20000
rect 1504 27 1533 19973
rect 1579 27 1608 19973
rect 1504 0 1608 27
rect 1808 19973 1912 20000
rect 1808 27 1837 19973
rect 1883 27 1912 19973
rect 1808 0 1912 27
rect 2112 19973 2216 20000
rect 2112 27 2141 19973
rect 2187 27 2216 19973
rect 2112 0 2216 27
rect 2416 19973 2520 20000
rect 2416 27 2445 19973
rect 2491 27 2520 19973
rect 2416 0 2520 27
rect 2720 19973 2824 20000
rect 2720 27 2749 19973
rect 2795 27 2824 19973
rect 2720 0 2824 27
rect 3024 19973 3128 20000
rect 3024 27 3053 19973
rect 3099 27 3128 19973
rect 3024 0 3128 27
rect 3328 19973 3432 20000
rect 3328 27 3357 19973
rect 3403 27 3432 19973
rect 3328 0 3432 27
rect 3632 19973 3736 20000
rect 3632 27 3661 19973
rect 3707 27 3736 19973
rect 3632 0 3736 27
rect 3936 19973 4040 20000
rect 3936 27 3965 19973
rect 4011 27 4040 19973
rect 3936 0 4040 27
rect 4240 19973 4344 20000
rect 4240 27 4269 19973
rect 4315 27 4344 19973
rect 4240 0 4344 27
rect 4544 19973 4648 20000
rect 4544 27 4573 19973
rect 4619 27 4648 19973
rect 4544 0 4648 27
rect 4848 19973 4952 20000
rect 4848 27 4877 19973
rect 4923 27 4952 19973
rect 4848 0 4952 27
rect 5152 19973 5256 20000
rect 5152 27 5181 19973
rect 5227 27 5256 19973
rect 5152 0 5256 27
rect 5456 19973 5560 20000
rect 5456 27 5485 19973
rect 5531 27 5560 19973
rect 5456 0 5560 27
rect 5760 19973 5864 20000
rect 5760 27 5789 19973
rect 5835 27 5864 19973
rect 5760 0 5864 27
rect 6064 19973 6168 20000
rect 6064 27 6093 19973
rect 6139 27 6168 19973
rect 6064 0 6168 27
rect 6368 19973 6472 20000
rect 6368 27 6397 19973
rect 6443 27 6472 19973
rect 6368 0 6472 27
rect 6672 19973 6776 20000
rect 6672 27 6701 19973
rect 6747 27 6776 19973
rect 6672 0 6776 27
rect 6976 19973 7080 20000
rect 6976 27 7005 19973
rect 7051 27 7080 19973
rect 6976 0 7080 27
rect 7280 19973 7384 20000
rect 7280 27 7309 19973
rect 7355 27 7384 19973
rect 7280 0 7384 27
rect 7584 19973 7688 20000
rect 7584 27 7613 19973
rect 7659 27 7688 19973
rect 7584 0 7688 27
rect 7888 19973 7992 20000
rect 7888 27 7917 19973
rect 7963 27 7992 19973
rect 7888 0 7992 27
rect 8192 19973 8296 20000
rect 8192 27 8221 19973
rect 8267 27 8296 19973
rect 8192 0 8296 27
rect 8496 19973 8600 20000
rect 8496 27 8525 19973
rect 8571 27 8600 19973
rect 8496 0 8600 27
rect 8800 19973 8904 20000
rect 8800 27 8829 19973
rect 8875 27 8904 19973
rect 8800 0 8904 27
rect 9104 19973 9208 20000
rect 9104 27 9133 19973
rect 9179 27 9208 19973
rect 9104 0 9208 27
rect 9408 19973 9512 20000
rect 9408 27 9437 19973
rect 9483 27 9512 19973
rect 9408 0 9512 27
rect 9712 19973 9816 20000
rect 9712 27 9741 19973
rect 9787 27 9816 19973
rect 9712 0 9816 27
rect 10016 19973 10120 20000
rect 10016 27 10045 19973
rect 10091 27 10120 19973
rect 10016 0 10120 27
rect 10320 19973 10424 20000
rect 10320 27 10349 19973
rect 10395 27 10424 19973
rect 10320 0 10424 27
rect 10624 19973 10728 20000
rect 10624 27 10653 19973
rect 10699 27 10728 19973
rect 10624 0 10728 27
rect 10928 19973 11032 20000
rect 10928 27 10957 19973
rect 11003 27 11032 19973
rect 10928 0 11032 27
rect 11232 19973 11336 20000
rect 11232 27 11261 19973
rect 11307 27 11336 19973
rect 11232 0 11336 27
rect 11536 19973 11640 20000
rect 11536 27 11565 19973
rect 11611 27 11640 19973
rect 11536 0 11640 27
rect 11840 19973 11944 20000
rect 11840 27 11869 19973
rect 11915 27 11944 19973
rect 11840 0 11944 27
rect 12144 19973 12248 20000
rect 12144 27 12173 19973
rect 12219 27 12248 19973
rect 12144 0 12248 27
rect 12448 19973 12552 20000
rect 12448 27 12477 19973
rect 12523 27 12552 19973
rect 12448 0 12552 27
rect 12752 19973 12856 20000
rect 12752 27 12781 19973
rect 12827 27 12856 19973
rect 12752 0 12856 27
rect 13056 19973 13160 20000
rect 13056 27 13085 19973
rect 13131 27 13160 19973
rect 13056 0 13160 27
rect 13360 19973 13464 20000
rect 13360 27 13389 19973
rect 13435 27 13464 19973
rect 13360 0 13464 27
rect 13664 19973 13768 20000
rect 13664 27 13693 19973
rect 13739 27 13768 19973
rect 13664 0 13768 27
rect 13968 19973 14072 20000
rect 13968 27 13997 19973
rect 14043 27 14072 19973
rect 13968 0 14072 27
rect 14272 19973 14376 20000
rect 14272 27 14301 19973
rect 14347 27 14376 19973
rect 14272 0 14376 27
rect 14576 19973 14680 20000
rect 14576 27 14605 19973
rect 14651 27 14680 19973
rect 14576 0 14680 27
rect 14880 19973 14984 20000
rect 14880 27 14909 19973
rect 14955 27 14984 19973
rect 14880 0 14984 27
rect 15184 19973 15288 20000
rect 15184 27 15213 19973
rect 15259 27 15288 19973
rect 15184 0 15288 27
rect 15488 19973 15592 20000
rect 15488 27 15517 19973
rect 15563 27 15592 19973
rect 15488 0 15592 27
rect 15792 19973 15896 20000
rect 15792 27 15821 19973
rect 15867 27 15896 19973
rect 15792 0 15896 27
rect 16096 19973 16200 20000
rect 16096 27 16125 19973
rect 16171 27 16200 19973
rect 16096 0 16200 27
rect 16400 19973 16504 20000
rect 16400 27 16429 19973
rect 16475 27 16504 19973
rect 16400 0 16504 27
rect 16704 19973 16808 20000
rect 16704 27 16733 19973
rect 16779 27 16808 19973
rect 16704 0 16808 27
rect 17008 19973 17112 20000
rect 17008 27 17037 19973
rect 17083 27 17112 19973
rect 17008 0 17112 27
rect 17312 19973 17416 20000
rect 17312 27 17341 19973
rect 17387 27 17416 19973
rect 17312 0 17416 27
rect 17616 19973 17720 20000
rect 17616 27 17645 19973
rect 17691 27 17720 19973
rect 17616 0 17720 27
rect 17920 19973 18024 20000
rect 17920 27 17949 19973
rect 17995 27 18024 19973
rect 17920 0 18024 27
rect 18224 19973 18328 20000
rect 18224 27 18253 19973
rect 18299 27 18328 19973
rect 18224 0 18328 27
rect 18528 19973 18632 20000
rect 18528 27 18557 19973
rect 18603 27 18632 19973
rect 18528 0 18632 27
rect 18832 19973 18936 20000
rect 18832 27 18861 19973
rect 18907 27 18936 19973
rect 18832 0 18936 27
rect 19136 19973 19240 20000
rect 19136 27 19165 19973
rect 19211 27 19240 19973
rect 19136 0 19240 27
rect 19440 19973 19544 20000
rect 19440 27 19469 19973
rect 19515 27 19544 19973
rect 19440 0 19544 27
rect 19744 19973 19848 20000
rect 19744 27 19773 19973
rect 19819 27 19848 19973
rect 19744 0 19848 27
rect 20048 19973 20152 20000
rect 20048 27 20077 19973
rect 20123 27 20152 19973
rect 20048 0 20152 27
rect 20352 19973 20456 20000
rect 20352 27 20381 19973
rect 20427 27 20456 19973
rect 20352 0 20456 27
rect 20656 19973 20760 20000
rect 20656 27 20685 19973
rect 20731 27 20760 19973
rect 20656 0 20760 27
rect 20960 19973 21064 20000
rect 20960 27 20989 19973
rect 21035 27 21064 19973
rect 20960 0 21064 27
rect 21264 19973 21368 20000
rect 21264 27 21293 19973
rect 21339 27 21368 19973
rect 21264 0 21368 27
rect 21568 19973 21672 20000
rect 21568 27 21597 19973
rect 21643 27 21672 19973
rect 21568 0 21672 27
rect 21872 19973 21976 20000
rect 21872 27 21901 19973
rect 21947 27 21976 19973
rect 21872 0 21976 27
rect 22176 19973 22280 20000
rect 22176 27 22205 19973
rect 22251 27 22280 19973
rect 22176 0 22280 27
rect 22480 19973 22584 20000
rect 22480 27 22509 19973
rect 22555 27 22584 19973
rect 22480 0 22584 27
rect 22784 19973 22888 20000
rect 22784 27 22813 19973
rect 22859 27 22888 19973
rect 22784 0 22888 27
rect 23088 19973 23192 20000
rect 23088 27 23117 19973
rect 23163 27 23192 19973
rect 23088 0 23192 27
rect 23392 19973 23496 20000
rect 23392 27 23421 19973
rect 23467 27 23496 19973
rect 23392 0 23496 27
rect 23696 19973 23800 20000
rect 23696 27 23725 19973
rect 23771 27 23800 19973
rect 23696 0 23800 27
rect 24000 19973 24104 20000
rect 24000 27 24029 19973
rect 24075 27 24104 19973
rect 24000 0 24104 27
rect 24304 19973 24408 20000
rect 24304 27 24333 19973
rect 24379 27 24408 19973
rect 24304 0 24408 27
rect 24608 19973 24712 20000
rect 24608 27 24637 19973
rect 24683 27 24712 19973
rect 24608 0 24712 27
rect 24912 19973 25016 20000
rect 24912 27 24941 19973
rect 24987 27 25016 19973
rect 24912 0 25016 27
rect 25216 19973 25320 20000
rect 25216 27 25245 19973
rect 25291 27 25320 19973
rect 25216 0 25320 27
rect 25520 19973 25624 20000
rect 25520 27 25549 19973
rect 25595 27 25624 19973
rect 25520 0 25624 27
rect 25824 19973 25928 20000
rect 25824 27 25853 19973
rect 25899 27 25928 19973
rect 25824 0 25928 27
rect 26128 19973 26232 20000
rect 26128 27 26157 19973
rect 26203 27 26232 19973
rect 26128 0 26232 27
rect 26432 19973 26536 20000
rect 26432 27 26461 19973
rect 26507 27 26536 19973
rect 26432 0 26536 27
rect 26736 19973 26840 20000
rect 26736 27 26765 19973
rect 26811 27 26840 19973
rect 26736 0 26840 27
rect 27040 19973 27144 20000
rect 27040 27 27069 19973
rect 27115 27 27144 19973
rect 27040 0 27144 27
rect 27344 19973 27448 20000
rect 27344 27 27373 19973
rect 27419 27 27448 19973
rect 27344 0 27448 27
rect 27648 19973 27752 20000
rect 27648 27 27677 19973
rect 27723 27 27752 19973
rect 27648 0 27752 27
rect 27952 19973 28056 20000
rect 27952 27 27981 19973
rect 28027 27 28056 19973
rect 27952 0 28056 27
rect 28256 19973 28360 20000
rect 28256 27 28285 19973
rect 28331 27 28360 19973
rect 28256 0 28360 27
rect 28560 19973 28664 20000
rect 28560 27 28589 19973
rect 28635 27 28664 19973
rect 28560 0 28664 27
rect 28864 19973 28968 20000
rect 28864 27 28893 19973
rect 28939 27 28968 19973
rect 28864 0 28968 27
rect 29168 19973 29272 20000
rect 29168 27 29197 19973
rect 29243 27 29272 19973
rect 29168 0 29272 27
rect 29472 19973 29576 20000
rect 29472 27 29501 19973
rect 29547 27 29576 19973
rect 29472 0 29576 27
rect 29776 19973 29880 20000
rect 29776 27 29805 19973
rect 29851 27 29880 19973
rect 29776 0 29880 27
rect 30080 19973 30184 20000
rect 30080 27 30109 19973
rect 30155 27 30184 19973
rect 30080 0 30184 27
rect 30384 19973 30472 20000
rect 30384 27 30413 19973
rect 30459 27 30472 19973
rect 30384 0 30472 27
<< ndiffc >>
rect 13 27 59 19973
rect 317 27 363 19973
rect 621 27 667 19973
rect 925 27 971 19973
rect 1229 27 1275 19973
rect 1533 27 1579 19973
rect 1837 27 1883 19973
rect 2141 27 2187 19973
rect 2445 27 2491 19973
rect 2749 27 2795 19973
rect 3053 27 3099 19973
rect 3357 27 3403 19973
rect 3661 27 3707 19973
rect 3965 27 4011 19973
rect 4269 27 4315 19973
rect 4573 27 4619 19973
rect 4877 27 4923 19973
rect 5181 27 5227 19973
rect 5485 27 5531 19973
rect 5789 27 5835 19973
rect 6093 27 6139 19973
rect 6397 27 6443 19973
rect 6701 27 6747 19973
rect 7005 27 7051 19973
rect 7309 27 7355 19973
rect 7613 27 7659 19973
rect 7917 27 7963 19973
rect 8221 27 8267 19973
rect 8525 27 8571 19973
rect 8829 27 8875 19973
rect 9133 27 9179 19973
rect 9437 27 9483 19973
rect 9741 27 9787 19973
rect 10045 27 10091 19973
rect 10349 27 10395 19973
rect 10653 27 10699 19973
rect 10957 27 11003 19973
rect 11261 27 11307 19973
rect 11565 27 11611 19973
rect 11869 27 11915 19973
rect 12173 27 12219 19973
rect 12477 27 12523 19973
rect 12781 27 12827 19973
rect 13085 27 13131 19973
rect 13389 27 13435 19973
rect 13693 27 13739 19973
rect 13997 27 14043 19973
rect 14301 27 14347 19973
rect 14605 27 14651 19973
rect 14909 27 14955 19973
rect 15213 27 15259 19973
rect 15517 27 15563 19973
rect 15821 27 15867 19973
rect 16125 27 16171 19973
rect 16429 27 16475 19973
rect 16733 27 16779 19973
rect 17037 27 17083 19973
rect 17341 27 17387 19973
rect 17645 27 17691 19973
rect 17949 27 17995 19973
rect 18253 27 18299 19973
rect 18557 27 18603 19973
rect 18861 27 18907 19973
rect 19165 27 19211 19973
rect 19469 27 19515 19973
rect 19773 27 19819 19973
rect 20077 27 20123 19973
rect 20381 27 20427 19973
rect 20685 27 20731 19973
rect 20989 27 21035 19973
rect 21293 27 21339 19973
rect 21597 27 21643 19973
rect 21901 27 21947 19973
rect 22205 27 22251 19973
rect 22509 27 22555 19973
rect 22813 27 22859 19973
rect 23117 27 23163 19973
rect 23421 27 23467 19973
rect 23725 27 23771 19973
rect 24029 27 24075 19973
rect 24333 27 24379 19973
rect 24637 27 24683 19973
rect 24941 27 24987 19973
rect 25245 27 25291 19973
rect 25549 27 25595 19973
rect 25853 27 25899 19973
rect 26157 27 26203 19973
rect 26461 27 26507 19973
rect 26765 27 26811 19973
rect 27069 27 27115 19973
rect 27373 27 27419 19973
rect 27677 27 27723 19973
rect 27981 27 28027 19973
rect 28285 27 28331 19973
rect 28589 27 28635 19973
rect 28893 27 28939 19973
rect 29197 27 29243 19973
rect 29501 27 29547 19973
rect 29805 27 29851 19973
rect 30109 27 30155 19973
rect 30413 27 30459 19973
<< psubdiff >>
rect -152 19973 -64 20000
rect -152 27 -131 19973
rect -85 27 -64 19973
rect -152 0 -64 27
<< psubdiffcont >>
rect -131 27 -85 19973
<< polysilicon >>
rect 88 20000 288 20044
rect 392 20000 592 20044
rect 696 20000 896 20044
rect 1000 20000 1200 20044
rect 1304 20000 1504 20044
rect 1608 20000 1808 20044
rect 1912 20000 2112 20044
rect 2216 20000 2416 20044
rect 2520 20000 2720 20044
rect 2824 20000 3024 20044
rect 3128 20000 3328 20044
rect 3432 20000 3632 20044
rect 3736 20000 3936 20044
rect 4040 20000 4240 20044
rect 4344 20000 4544 20044
rect 4648 20000 4848 20044
rect 4952 20000 5152 20044
rect 5256 20000 5456 20044
rect 5560 20000 5760 20044
rect 5864 20000 6064 20044
rect 6168 20000 6368 20044
rect 6472 20000 6672 20044
rect 6776 20000 6976 20044
rect 7080 20000 7280 20044
rect 7384 20000 7584 20044
rect 7688 20000 7888 20044
rect 7992 20000 8192 20044
rect 8296 20000 8496 20044
rect 8600 20000 8800 20044
rect 8904 20000 9104 20044
rect 9208 20000 9408 20044
rect 9512 20000 9712 20044
rect 9816 20000 10016 20044
rect 10120 20000 10320 20044
rect 10424 20000 10624 20044
rect 10728 20000 10928 20044
rect 11032 20000 11232 20044
rect 11336 20000 11536 20044
rect 11640 20000 11840 20044
rect 11944 20000 12144 20044
rect 12248 20000 12448 20044
rect 12552 20000 12752 20044
rect 12856 20000 13056 20044
rect 13160 20000 13360 20044
rect 13464 20000 13664 20044
rect 13768 20000 13968 20044
rect 14072 20000 14272 20044
rect 14376 20000 14576 20044
rect 14680 20000 14880 20044
rect 14984 20000 15184 20044
rect 15288 20000 15488 20044
rect 15592 20000 15792 20044
rect 15896 20000 16096 20044
rect 16200 20000 16400 20044
rect 16504 20000 16704 20044
rect 16808 20000 17008 20044
rect 17112 20000 17312 20044
rect 17416 20000 17616 20044
rect 17720 20000 17920 20044
rect 18024 20000 18224 20044
rect 18328 20000 18528 20044
rect 18632 20000 18832 20044
rect 18936 20000 19136 20044
rect 19240 20000 19440 20044
rect 19544 20000 19744 20044
rect 19848 20000 20048 20044
rect 20152 20000 20352 20044
rect 20456 20000 20656 20044
rect 20760 20000 20960 20044
rect 21064 20000 21264 20044
rect 21368 20000 21568 20044
rect 21672 20000 21872 20044
rect 21976 20000 22176 20044
rect 22280 20000 22480 20044
rect 22584 20000 22784 20044
rect 22888 20000 23088 20044
rect 23192 20000 23392 20044
rect 23496 20000 23696 20044
rect 23800 20000 24000 20044
rect 24104 20000 24304 20044
rect 24408 20000 24608 20044
rect 24712 20000 24912 20044
rect 25016 20000 25216 20044
rect 25320 20000 25520 20044
rect 25624 20000 25824 20044
rect 25928 20000 26128 20044
rect 26232 20000 26432 20044
rect 26536 20000 26736 20044
rect 26840 20000 27040 20044
rect 27144 20000 27344 20044
rect 27448 20000 27648 20044
rect 27752 20000 27952 20044
rect 28056 20000 28256 20044
rect 28360 20000 28560 20044
rect 28664 20000 28864 20044
rect 28968 20000 29168 20044
rect 29272 20000 29472 20044
rect 29576 20000 29776 20044
rect 29880 20000 30080 20044
rect 30184 20000 30384 20044
rect 88 -44 288 0
rect 392 -44 592 0
rect 696 -44 896 0
rect 1000 -44 1200 0
rect 1304 -44 1504 0
rect 1608 -44 1808 0
rect 1912 -44 2112 0
rect 2216 -44 2416 0
rect 2520 -44 2720 0
rect 2824 -44 3024 0
rect 3128 -44 3328 0
rect 3432 -44 3632 0
rect 3736 -44 3936 0
rect 4040 -44 4240 0
rect 4344 -44 4544 0
rect 4648 -44 4848 0
rect 4952 -44 5152 0
rect 5256 -44 5456 0
rect 5560 -44 5760 0
rect 5864 -44 6064 0
rect 6168 -44 6368 0
rect 6472 -44 6672 0
rect 6776 -44 6976 0
rect 7080 -44 7280 0
rect 7384 -44 7584 0
rect 7688 -44 7888 0
rect 7992 -44 8192 0
rect 8296 -44 8496 0
rect 8600 -44 8800 0
rect 8904 -44 9104 0
rect 9208 -44 9408 0
rect 9512 -44 9712 0
rect 9816 -44 10016 0
rect 10120 -44 10320 0
rect 10424 -44 10624 0
rect 10728 -44 10928 0
rect 11032 -44 11232 0
rect 11336 -44 11536 0
rect 11640 -44 11840 0
rect 11944 -44 12144 0
rect 12248 -44 12448 0
rect 12552 -44 12752 0
rect 12856 -44 13056 0
rect 13160 -44 13360 0
rect 13464 -44 13664 0
rect 13768 -44 13968 0
rect 14072 -44 14272 0
rect 14376 -44 14576 0
rect 14680 -44 14880 0
rect 14984 -44 15184 0
rect 15288 -44 15488 0
rect 15592 -44 15792 0
rect 15896 -44 16096 0
rect 16200 -44 16400 0
rect 16504 -44 16704 0
rect 16808 -44 17008 0
rect 17112 -44 17312 0
rect 17416 -44 17616 0
rect 17720 -44 17920 0
rect 18024 -44 18224 0
rect 18328 -44 18528 0
rect 18632 -44 18832 0
rect 18936 -44 19136 0
rect 19240 -44 19440 0
rect 19544 -44 19744 0
rect 19848 -44 20048 0
rect 20152 -44 20352 0
rect 20456 -44 20656 0
rect 20760 -44 20960 0
rect 21064 -44 21264 0
rect 21368 -44 21568 0
rect 21672 -44 21872 0
rect 21976 -44 22176 0
rect 22280 -44 22480 0
rect 22584 -44 22784 0
rect 22888 -44 23088 0
rect 23192 -44 23392 0
rect 23496 -44 23696 0
rect 23800 -44 24000 0
rect 24104 -44 24304 0
rect 24408 -44 24608 0
rect 24712 -44 24912 0
rect 25016 -44 25216 0
rect 25320 -44 25520 0
rect 25624 -44 25824 0
rect 25928 -44 26128 0
rect 26232 -44 26432 0
rect 26536 -44 26736 0
rect 26840 -44 27040 0
rect 27144 -44 27344 0
rect 27448 -44 27648 0
rect 27752 -44 27952 0
rect 28056 -44 28256 0
rect 28360 -44 28560 0
rect 28664 -44 28864 0
rect 28968 -44 29168 0
rect 29272 -44 29472 0
rect 29576 -44 29776 0
rect 29880 -44 30080 0
rect 30184 -44 30384 0
<< metal1 >>
rect -152 19973 -64 20000
rect -152 27 -131 19973
rect -85 27 -64 19973
rect -152 0 -64 27
rect -2 19973 74 20002
rect -2 27 13 19973
rect 59 27 74 19973
rect -2 -2 74 27
rect 302 19973 378 20002
rect 302 27 317 19973
rect 363 27 378 19973
rect 302 -2 378 27
rect 606 19973 682 20002
rect 606 27 621 19973
rect 667 27 682 19973
rect 606 -2 682 27
rect 910 19973 986 20002
rect 910 27 925 19973
rect 971 27 986 19973
rect 910 -2 986 27
rect 1214 19973 1290 20002
rect 1214 27 1229 19973
rect 1275 27 1290 19973
rect 1214 -2 1290 27
rect 1518 19973 1594 20002
rect 1518 27 1533 19973
rect 1579 27 1594 19973
rect 1518 -2 1594 27
rect 1822 19973 1898 20002
rect 1822 27 1837 19973
rect 1883 27 1898 19973
rect 1822 -2 1898 27
rect 2126 19973 2202 20002
rect 2126 27 2141 19973
rect 2187 27 2202 19973
rect 2126 -2 2202 27
rect 2430 19973 2506 20002
rect 2430 27 2445 19973
rect 2491 27 2506 19973
rect 2430 -2 2506 27
rect 2734 19973 2810 20002
rect 2734 27 2749 19973
rect 2795 27 2810 19973
rect 2734 -2 2810 27
rect 3038 19973 3114 20002
rect 3038 27 3053 19973
rect 3099 27 3114 19973
rect 3038 -2 3114 27
rect 3342 19973 3418 20002
rect 3342 27 3357 19973
rect 3403 27 3418 19973
rect 3342 -2 3418 27
rect 3646 19973 3722 20002
rect 3646 27 3661 19973
rect 3707 27 3722 19973
rect 3646 -2 3722 27
rect 3950 19973 4026 20002
rect 3950 27 3965 19973
rect 4011 27 4026 19973
rect 3950 -2 4026 27
rect 4254 19973 4330 20002
rect 4254 27 4269 19973
rect 4315 27 4330 19973
rect 4254 -2 4330 27
rect 4558 19973 4634 20002
rect 4558 27 4573 19973
rect 4619 27 4634 19973
rect 4558 -2 4634 27
rect 4862 19973 4938 20002
rect 4862 27 4877 19973
rect 4923 27 4938 19973
rect 4862 -2 4938 27
rect 5166 19973 5242 20002
rect 5166 27 5181 19973
rect 5227 27 5242 19973
rect 5166 -2 5242 27
rect 5470 19973 5546 20002
rect 5470 27 5485 19973
rect 5531 27 5546 19973
rect 5470 -2 5546 27
rect 5774 19973 5850 20002
rect 5774 27 5789 19973
rect 5835 27 5850 19973
rect 5774 -2 5850 27
rect 6078 19973 6154 20002
rect 6078 27 6093 19973
rect 6139 27 6154 19973
rect 6078 -2 6154 27
rect 6382 19973 6458 20002
rect 6382 27 6397 19973
rect 6443 27 6458 19973
rect 6382 -2 6458 27
rect 6686 19973 6762 20002
rect 6686 27 6701 19973
rect 6747 27 6762 19973
rect 6686 -2 6762 27
rect 6990 19973 7066 20002
rect 6990 27 7005 19973
rect 7051 27 7066 19973
rect 6990 -2 7066 27
rect 7294 19973 7370 20002
rect 7294 27 7309 19973
rect 7355 27 7370 19973
rect 7294 -2 7370 27
rect 7598 19973 7674 20002
rect 7598 27 7613 19973
rect 7659 27 7674 19973
rect 7598 -2 7674 27
rect 7902 19973 7978 20002
rect 7902 27 7917 19973
rect 7963 27 7978 19973
rect 7902 -2 7978 27
rect 8206 19973 8282 20002
rect 8206 27 8221 19973
rect 8267 27 8282 19973
rect 8206 -2 8282 27
rect 8510 19973 8586 20002
rect 8510 27 8525 19973
rect 8571 27 8586 19973
rect 8510 -2 8586 27
rect 8814 19973 8890 20002
rect 8814 27 8829 19973
rect 8875 27 8890 19973
rect 8814 -2 8890 27
rect 9118 19973 9194 20002
rect 9118 27 9133 19973
rect 9179 27 9194 19973
rect 9118 -2 9194 27
rect 9422 19973 9498 20002
rect 9422 27 9437 19973
rect 9483 27 9498 19973
rect 9422 -2 9498 27
rect 9726 19973 9802 20002
rect 9726 27 9741 19973
rect 9787 27 9802 19973
rect 9726 -2 9802 27
rect 10030 19973 10106 20002
rect 10030 27 10045 19973
rect 10091 27 10106 19973
rect 10030 -2 10106 27
rect 10334 19973 10410 20002
rect 10334 27 10349 19973
rect 10395 27 10410 19973
rect 10334 -2 10410 27
rect 10638 19973 10714 20002
rect 10638 27 10653 19973
rect 10699 27 10714 19973
rect 10638 -2 10714 27
rect 10942 19973 11018 20002
rect 10942 27 10957 19973
rect 11003 27 11018 19973
rect 10942 -2 11018 27
rect 11246 19973 11322 20002
rect 11246 27 11261 19973
rect 11307 27 11322 19973
rect 11246 -2 11322 27
rect 11550 19973 11626 20002
rect 11550 27 11565 19973
rect 11611 27 11626 19973
rect 11550 -2 11626 27
rect 11854 19973 11930 20002
rect 11854 27 11869 19973
rect 11915 27 11930 19973
rect 11854 -2 11930 27
rect 12158 19973 12234 20002
rect 12158 27 12173 19973
rect 12219 27 12234 19973
rect 12158 -2 12234 27
rect 12462 19973 12538 20002
rect 12462 27 12477 19973
rect 12523 27 12538 19973
rect 12462 -2 12538 27
rect 12766 19973 12842 20002
rect 12766 27 12781 19973
rect 12827 27 12842 19973
rect 12766 -2 12842 27
rect 13070 19973 13146 20002
rect 13070 27 13085 19973
rect 13131 27 13146 19973
rect 13070 -2 13146 27
rect 13374 19973 13450 20002
rect 13374 27 13389 19973
rect 13435 27 13450 19973
rect 13374 -2 13450 27
rect 13678 19973 13754 20002
rect 13678 27 13693 19973
rect 13739 27 13754 19973
rect 13678 -2 13754 27
rect 13982 19973 14058 20002
rect 13982 27 13997 19973
rect 14043 27 14058 19973
rect 13982 -2 14058 27
rect 14286 19973 14362 20002
rect 14286 27 14301 19973
rect 14347 27 14362 19973
rect 14286 -2 14362 27
rect 14590 19973 14666 20002
rect 14590 27 14605 19973
rect 14651 27 14666 19973
rect 14590 -2 14666 27
rect 14894 19973 14970 20002
rect 14894 27 14909 19973
rect 14955 27 14970 19973
rect 14894 -2 14970 27
rect 15198 19973 15274 20002
rect 15198 27 15213 19973
rect 15259 27 15274 19973
rect 15198 -2 15274 27
rect 15502 19973 15578 20002
rect 15502 27 15517 19973
rect 15563 27 15578 19973
rect 15502 -2 15578 27
rect 15806 19973 15882 20002
rect 15806 27 15821 19973
rect 15867 27 15882 19973
rect 15806 -2 15882 27
rect 16110 19973 16186 20002
rect 16110 27 16125 19973
rect 16171 27 16186 19973
rect 16110 -2 16186 27
rect 16414 19973 16490 20002
rect 16414 27 16429 19973
rect 16475 27 16490 19973
rect 16414 -2 16490 27
rect 16718 19973 16794 20002
rect 16718 27 16733 19973
rect 16779 27 16794 19973
rect 16718 -2 16794 27
rect 17022 19973 17098 20002
rect 17022 27 17037 19973
rect 17083 27 17098 19973
rect 17022 -2 17098 27
rect 17326 19973 17402 20002
rect 17326 27 17341 19973
rect 17387 27 17402 19973
rect 17326 -2 17402 27
rect 17630 19973 17706 20002
rect 17630 27 17645 19973
rect 17691 27 17706 19973
rect 17630 -2 17706 27
rect 17934 19973 18010 20002
rect 17934 27 17949 19973
rect 17995 27 18010 19973
rect 17934 -2 18010 27
rect 18238 19973 18314 20002
rect 18238 27 18253 19973
rect 18299 27 18314 19973
rect 18238 -2 18314 27
rect 18542 19973 18618 20002
rect 18542 27 18557 19973
rect 18603 27 18618 19973
rect 18542 -2 18618 27
rect 18846 19973 18922 20002
rect 18846 27 18861 19973
rect 18907 27 18922 19973
rect 18846 -2 18922 27
rect 19150 19973 19226 20002
rect 19150 27 19165 19973
rect 19211 27 19226 19973
rect 19150 -2 19226 27
rect 19454 19973 19530 20002
rect 19454 27 19469 19973
rect 19515 27 19530 19973
rect 19454 -2 19530 27
rect 19758 19973 19834 20002
rect 19758 27 19773 19973
rect 19819 27 19834 19973
rect 19758 -2 19834 27
rect 20062 19973 20138 20002
rect 20062 27 20077 19973
rect 20123 27 20138 19973
rect 20062 -2 20138 27
rect 20366 19973 20442 20002
rect 20366 27 20381 19973
rect 20427 27 20442 19973
rect 20366 -2 20442 27
rect 20670 19973 20746 20002
rect 20670 27 20685 19973
rect 20731 27 20746 19973
rect 20670 -2 20746 27
rect 20974 19973 21050 20002
rect 20974 27 20989 19973
rect 21035 27 21050 19973
rect 20974 -2 21050 27
rect 21278 19973 21354 20002
rect 21278 27 21293 19973
rect 21339 27 21354 19973
rect 21278 -2 21354 27
rect 21582 19973 21658 20002
rect 21582 27 21597 19973
rect 21643 27 21658 19973
rect 21582 -2 21658 27
rect 21886 19973 21962 20002
rect 21886 27 21901 19973
rect 21947 27 21962 19973
rect 21886 -2 21962 27
rect 22190 19973 22266 20002
rect 22190 27 22205 19973
rect 22251 27 22266 19973
rect 22190 -2 22266 27
rect 22494 19973 22570 20002
rect 22494 27 22509 19973
rect 22555 27 22570 19973
rect 22494 -2 22570 27
rect 22798 19973 22874 20002
rect 22798 27 22813 19973
rect 22859 27 22874 19973
rect 22798 -2 22874 27
rect 23102 19973 23178 20002
rect 23102 27 23117 19973
rect 23163 27 23178 19973
rect 23102 -2 23178 27
rect 23406 19973 23482 20002
rect 23406 27 23421 19973
rect 23467 27 23482 19973
rect 23406 -2 23482 27
rect 23710 19973 23786 20002
rect 23710 27 23725 19973
rect 23771 27 23786 19973
rect 23710 -2 23786 27
rect 24014 19973 24090 20002
rect 24014 27 24029 19973
rect 24075 27 24090 19973
rect 24014 -2 24090 27
rect 24318 19973 24394 20002
rect 24318 27 24333 19973
rect 24379 27 24394 19973
rect 24318 -2 24394 27
rect 24622 19973 24698 20002
rect 24622 27 24637 19973
rect 24683 27 24698 19973
rect 24622 -2 24698 27
rect 24926 19973 25002 20002
rect 24926 27 24941 19973
rect 24987 27 25002 19973
rect 24926 -2 25002 27
rect 25230 19973 25306 20002
rect 25230 27 25245 19973
rect 25291 27 25306 19973
rect 25230 -2 25306 27
rect 25534 19973 25610 20002
rect 25534 27 25549 19973
rect 25595 27 25610 19973
rect 25534 -2 25610 27
rect 25838 19973 25914 20002
rect 25838 27 25853 19973
rect 25899 27 25914 19973
rect 25838 -2 25914 27
rect 26142 19973 26218 20002
rect 26142 27 26157 19973
rect 26203 27 26218 19973
rect 26142 -2 26218 27
rect 26446 19973 26522 20002
rect 26446 27 26461 19973
rect 26507 27 26522 19973
rect 26446 -2 26522 27
rect 26750 19973 26826 20002
rect 26750 27 26765 19973
rect 26811 27 26826 19973
rect 26750 -2 26826 27
rect 27054 19973 27130 20002
rect 27054 27 27069 19973
rect 27115 27 27130 19973
rect 27054 -2 27130 27
rect 27358 19973 27434 20002
rect 27358 27 27373 19973
rect 27419 27 27434 19973
rect 27358 -2 27434 27
rect 27662 19973 27738 20002
rect 27662 27 27677 19973
rect 27723 27 27738 19973
rect 27662 -2 27738 27
rect 27966 19973 28042 20002
rect 27966 27 27981 19973
rect 28027 27 28042 19973
rect 27966 -2 28042 27
rect 28270 19973 28346 20002
rect 28270 27 28285 19973
rect 28331 27 28346 19973
rect 28270 -2 28346 27
rect 28574 19973 28650 20002
rect 28574 27 28589 19973
rect 28635 27 28650 19973
rect 28574 -2 28650 27
rect 28878 19973 28954 20002
rect 28878 27 28893 19973
rect 28939 27 28954 19973
rect 28878 -2 28954 27
rect 29182 19973 29258 20002
rect 29182 27 29197 19973
rect 29243 27 29258 19973
rect 29182 -2 29258 27
rect 29486 19973 29562 20002
rect 29486 27 29501 19973
rect 29547 27 29562 19973
rect 29486 -2 29562 27
rect 29790 19973 29866 20002
rect 29790 27 29805 19973
rect 29851 27 29866 19973
rect 29790 -2 29866 27
rect 30094 19973 30170 20002
rect 30094 27 30109 19973
rect 30155 27 30170 19973
rect 30094 -2 30170 27
rect 30398 19973 30474 20002
rect 30398 27 30413 19973
rect 30459 27 30474 19973
rect 30398 -2 30474 27
<< end >>
