magic
tech gf180mcuC
magscale 1 10
timestamp 1676577649
<< error_p >>
rect -66 0 -64 10000
rect 0 0 2 10000
<< nwell >>
rect -176 -86 25358 10086
<< pmos >>
rect 88 0 488 10000
rect 592 0 992 10000
rect 1096 0 1496 10000
rect 1600 0 2000 10000
rect 2104 0 2504 10000
rect 2608 0 3008 10000
rect 3112 0 3512 10000
rect 3616 0 4016 10000
rect 4120 0 4520 10000
rect 4624 0 5024 10000
rect 5128 0 5528 10000
rect 5632 0 6032 10000
rect 6136 0 6536 10000
rect 6640 0 7040 10000
rect 7144 0 7544 10000
rect 7648 0 8048 10000
rect 8152 0 8552 10000
rect 8656 0 9056 10000
rect 9160 0 9560 10000
rect 9664 0 10064 10000
rect 10168 0 10568 10000
rect 10672 0 11072 10000
rect 11176 0 11576 10000
rect 11680 0 12080 10000
rect 12184 0 12584 10000
rect 12688 0 13088 10000
rect 13192 0 13592 10000
rect 13696 0 14096 10000
rect 14200 0 14600 10000
rect 14704 0 15104 10000
rect 15208 0 15608 10000
rect 15712 0 16112 10000
rect 16216 0 16616 10000
rect 16720 0 17120 10000
rect 17224 0 17624 10000
rect 17728 0 18128 10000
rect 18232 0 18632 10000
rect 18736 0 19136 10000
rect 19240 0 19640 10000
rect 19744 0 20144 10000
rect 20248 0 20648 10000
rect 20752 0 21152 10000
rect 21256 0 21656 10000
rect 21760 0 22160 10000
rect 22264 0 22664 10000
rect 22768 0 23168 10000
rect 23272 0 23672 10000
rect 23776 0 24176 10000
rect 24280 0 24680 10000
rect 24784 0 25184 10000
<< pdiff >>
rect 0 9973 88 10000
rect 0 27 13 9973
rect 59 27 88 9973
rect 0 0 88 27
rect 488 9973 592 10000
rect 488 27 517 9973
rect 563 27 592 9973
rect 488 0 592 27
rect 992 9973 1096 10000
rect 992 27 1021 9973
rect 1067 27 1096 9973
rect 992 0 1096 27
rect 1496 9973 1600 10000
rect 1496 27 1525 9973
rect 1571 27 1600 9973
rect 1496 0 1600 27
rect 2000 9973 2104 10000
rect 2000 27 2029 9973
rect 2075 27 2104 9973
rect 2000 0 2104 27
rect 2504 9973 2608 10000
rect 2504 27 2533 9973
rect 2579 27 2608 9973
rect 2504 0 2608 27
rect 3008 9973 3112 10000
rect 3008 27 3037 9973
rect 3083 27 3112 9973
rect 3008 0 3112 27
rect 3512 9973 3616 10000
rect 3512 27 3541 9973
rect 3587 27 3616 9973
rect 3512 0 3616 27
rect 4016 9973 4120 10000
rect 4016 27 4045 9973
rect 4091 27 4120 9973
rect 4016 0 4120 27
rect 4520 9973 4624 10000
rect 4520 27 4549 9973
rect 4595 27 4624 9973
rect 4520 0 4624 27
rect 5024 9973 5128 10000
rect 5024 27 5053 9973
rect 5099 27 5128 9973
rect 5024 0 5128 27
rect 5528 9973 5632 10000
rect 5528 27 5557 9973
rect 5603 27 5632 9973
rect 5528 0 5632 27
rect 6032 9973 6136 10000
rect 6032 27 6061 9973
rect 6107 27 6136 9973
rect 6032 0 6136 27
rect 6536 9973 6640 10000
rect 6536 27 6565 9973
rect 6611 27 6640 9973
rect 6536 0 6640 27
rect 7040 9973 7144 10000
rect 7040 27 7069 9973
rect 7115 27 7144 9973
rect 7040 0 7144 27
rect 7544 9973 7648 10000
rect 7544 27 7573 9973
rect 7619 27 7648 9973
rect 7544 0 7648 27
rect 8048 9973 8152 10000
rect 8048 27 8077 9973
rect 8123 27 8152 9973
rect 8048 0 8152 27
rect 8552 9973 8656 10000
rect 8552 27 8581 9973
rect 8627 27 8656 9973
rect 8552 0 8656 27
rect 9056 9973 9160 10000
rect 9056 27 9085 9973
rect 9131 27 9160 9973
rect 9056 0 9160 27
rect 9560 9973 9664 10000
rect 9560 27 9589 9973
rect 9635 27 9664 9973
rect 9560 0 9664 27
rect 10064 9973 10168 10000
rect 10064 27 10093 9973
rect 10139 27 10168 9973
rect 10064 0 10168 27
rect 10568 9973 10672 10000
rect 10568 27 10597 9973
rect 10643 27 10672 9973
rect 10568 0 10672 27
rect 11072 9973 11176 10000
rect 11072 27 11101 9973
rect 11147 27 11176 9973
rect 11072 0 11176 27
rect 11576 9973 11680 10000
rect 11576 27 11605 9973
rect 11651 27 11680 9973
rect 11576 0 11680 27
rect 12080 9973 12184 10000
rect 12080 27 12109 9973
rect 12155 27 12184 9973
rect 12080 0 12184 27
rect 12584 9973 12688 10000
rect 12584 27 12613 9973
rect 12659 27 12688 9973
rect 12584 0 12688 27
rect 13088 9973 13192 10000
rect 13088 27 13117 9973
rect 13163 27 13192 9973
rect 13088 0 13192 27
rect 13592 9973 13696 10000
rect 13592 27 13621 9973
rect 13667 27 13696 9973
rect 13592 0 13696 27
rect 14096 9973 14200 10000
rect 14096 27 14125 9973
rect 14171 27 14200 9973
rect 14096 0 14200 27
rect 14600 9973 14704 10000
rect 14600 27 14629 9973
rect 14675 27 14704 9973
rect 14600 0 14704 27
rect 15104 9973 15208 10000
rect 15104 27 15133 9973
rect 15179 27 15208 9973
rect 15104 0 15208 27
rect 15608 9973 15712 10000
rect 15608 27 15637 9973
rect 15683 27 15712 9973
rect 15608 0 15712 27
rect 16112 9973 16216 10000
rect 16112 27 16141 9973
rect 16187 27 16216 9973
rect 16112 0 16216 27
rect 16616 9973 16720 10000
rect 16616 27 16645 9973
rect 16691 27 16720 9973
rect 16616 0 16720 27
rect 17120 9973 17224 10000
rect 17120 27 17149 9973
rect 17195 27 17224 9973
rect 17120 0 17224 27
rect 17624 9973 17728 10000
rect 17624 27 17653 9973
rect 17699 27 17728 9973
rect 17624 0 17728 27
rect 18128 9973 18232 10000
rect 18128 27 18157 9973
rect 18203 27 18232 9973
rect 18128 0 18232 27
rect 18632 9973 18736 10000
rect 18632 27 18661 9973
rect 18707 27 18736 9973
rect 18632 0 18736 27
rect 19136 9973 19240 10000
rect 19136 27 19165 9973
rect 19211 27 19240 9973
rect 19136 0 19240 27
rect 19640 9973 19744 10000
rect 19640 27 19669 9973
rect 19715 27 19744 9973
rect 19640 0 19744 27
rect 20144 9973 20248 10000
rect 20144 27 20173 9973
rect 20219 27 20248 9973
rect 20144 0 20248 27
rect 20648 9973 20752 10000
rect 20648 27 20677 9973
rect 20723 27 20752 9973
rect 20648 0 20752 27
rect 21152 9973 21256 10000
rect 21152 27 21181 9973
rect 21227 27 21256 9973
rect 21152 0 21256 27
rect 21656 9973 21760 10000
rect 21656 27 21685 9973
rect 21731 27 21760 9973
rect 21656 0 21760 27
rect 22160 9973 22264 10000
rect 22160 27 22189 9973
rect 22235 27 22264 9973
rect 22160 0 22264 27
rect 22664 9973 22768 10000
rect 22664 27 22693 9973
rect 22739 27 22768 9973
rect 22664 0 22768 27
rect 23168 9973 23272 10000
rect 23168 27 23197 9973
rect 23243 27 23272 9973
rect 23168 0 23272 27
rect 23672 9973 23776 10000
rect 23672 27 23701 9973
rect 23747 27 23776 9973
rect 23672 0 23776 27
rect 24176 9973 24280 10000
rect 24176 27 24205 9973
rect 24251 27 24280 9973
rect 24176 0 24280 27
rect 24680 9973 24784 10000
rect 24680 27 24709 9973
rect 24755 27 24784 9973
rect 24680 0 24784 27
rect 25184 9973 25272 10000
rect 25184 27 25213 9973
rect 25259 27 25272 9973
rect 25184 0 25272 27
<< pdiffc >>
rect 13 27 59 9973
rect 517 27 563 9973
rect 1021 27 1067 9973
rect 1525 27 1571 9973
rect 2029 27 2075 9973
rect 2533 27 2579 9973
rect 3037 27 3083 9973
rect 3541 27 3587 9973
rect 4045 27 4091 9973
rect 4549 27 4595 9973
rect 5053 27 5099 9973
rect 5557 27 5603 9973
rect 6061 27 6107 9973
rect 6565 27 6611 9973
rect 7069 27 7115 9973
rect 7573 27 7619 9973
rect 8077 27 8123 9973
rect 8581 27 8627 9973
rect 9085 27 9131 9973
rect 9589 27 9635 9973
rect 10093 27 10139 9973
rect 10597 27 10643 9973
rect 11101 27 11147 9973
rect 11605 27 11651 9973
rect 12109 27 12155 9973
rect 12613 27 12659 9973
rect 13117 27 13163 9973
rect 13621 27 13667 9973
rect 14125 27 14171 9973
rect 14629 27 14675 9973
rect 15133 27 15179 9973
rect 15637 27 15683 9973
rect 16141 27 16187 9973
rect 16645 27 16691 9973
rect 17149 27 17195 9973
rect 17653 27 17699 9973
rect 18157 27 18203 9973
rect 18661 27 18707 9973
rect 19165 27 19211 9973
rect 19669 27 19715 9973
rect 20173 27 20219 9973
rect 20677 27 20723 9973
rect 21181 27 21227 9973
rect 21685 27 21731 9973
rect 22189 27 22235 9973
rect 22693 27 22739 9973
rect 23197 27 23243 9973
rect 23701 27 23747 9973
rect 24205 27 24251 9973
rect 24709 27 24755 9973
rect 25213 27 25259 9973
<< nsubdiff >>
rect -152 9973 -64 10000
rect -152 27 -131 9973
rect -85 27 -64 9973
rect -152 0 -64 27
<< nsubdiffcont >>
rect -131 27 -85 9973
<< polysilicon >>
rect 88 10000 488 10044
rect 592 10000 992 10044
rect 1096 10000 1496 10044
rect 1600 10000 2000 10044
rect 2104 10000 2504 10044
rect 2608 10000 3008 10044
rect 3112 10000 3512 10044
rect 3616 10000 4016 10044
rect 4120 10000 4520 10044
rect 4624 10000 5024 10044
rect 5128 10000 5528 10044
rect 5632 10000 6032 10044
rect 6136 10000 6536 10044
rect 6640 10000 7040 10044
rect 7144 10000 7544 10044
rect 7648 10000 8048 10044
rect 8152 10000 8552 10044
rect 8656 10000 9056 10044
rect 9160 10000 9560 10044
rect 9664 10000 10064 10044
rect 10168 10000 10568 10044
rect 10672 10000 11072 10044
rect 11176 10000 11576 10044
rect 11680 10000 12080 10044
rect 12184 10000 12584 10044
rect 12688 10000 13088 10044
rect 13192 10000 13592 10044
rect 13696 10000 14096 10044
rect 14200 10000 14600 10044
rect 14704 10000 15104 10044
rect 15208 10000 15608 10044
rect 15712 10000 16112 10044
rect 16216 10000 16616 10044
rect 16720 10000 17120 10044
rect 17224 10000 17624 10044
rect 17728 10000 18128 10044
rect 18232 10000 18632 10044
rect 18736 10000 19136 10044
rect 19240 10000 19640 10044
rect 19744 10000 20144 10044
rect 20248 10000 20648 10044
rect 20752 10000 21152 10044
rect 21256 10000 21656 10044
rect 21760 10000 22160 10044
rect 22264 10000 22664 10044
rect 22768 10000 23168 10044
rect 23272 10000 23672 10044
rect 23776 10000 24176 10044
rect 24280 10000 24680 10044
rect 24784 10000 25184 10044
rect 88 -44 488 0
rect 592 -44 992 0
rect 1096 -44 1496 0
rect 1600 -44 2000 0
rect 2104 -44 2504 0
rect 2608 -44 3008 0
rect 3112 -44 3512 0
rect 3616 -44 4016 0
rect 4120 -44 4520 0
rect 4624 -44 5024 0
rect 5128 -44 5528 0
rect 5632 -44 6032 0
rect 6136 -44 6536 0
rect 6640 -44 7040 0
rect 7144 -44 7544 0
rect 7648 -44 8048 0
rect 8152 -44 8552 0
rect 8656 -44 9056 0
rect 9160 -44 9560 0
rect 9664 -44 10064 0
rect 10168 -44 10568 0
rect 10672 -44 11072 0
rect 11176 -44 11576 0
rect 11680 -44 12080 0
rect 12184 -44 12584 0
rect 12688 -44 13088 0
rect 13192 -44 13592 0
rect 13696 -44 14096 0
rect 14200 -44 14600 0
rect 14704 -44 15104 0
rect 15208 -44 15608 0
rect 15712 -44 16112 0
rect 16216 -44 16616 0
rect 16720 -44 17120 0
rect 17224 -44 17624 0
rect 17728 -44 18128 0
rect 18232 -44 18632 0
rect 18736 -44 19136 0
rect 19240 -44 19640 0
rect 19744 -44 20144 0
rect 20248 -44 20648 0
rect 20752 -44 21152 0
rect 21256 -44 21656 0
rect 21760 -44 22160 0
rect 22264 -44 22664 0
rect 22768 -44 23168 0
rect 23272 -44 23672 0
rect 23776 -44 24176 0
rect 24280 -44 24680 0
rect 24784 -44 25184 0
<< metal1 >>
rect -152 9973 -64 10000
rect -152 27 -131 9973
rect -85 27 -64 9973
rect -152 0 -64 27
rect -2 9973 74 10002
rect -2 27 13 9973
rect 59 27 74 9973
rect -2 -2 74 27
rect 502 9973 578 10002
rect 502 27 517 9973
rect 563 27 578 9973
rect 502 -2 578 27
rect 1006 9973 1082 10002
rect 1006 27 1021 9973
rect 1067 27 1082 9973
rect 1006 -2 1082 27
rect 1510 9973 1586 10002
rect 1510 27 1525 9973
rect 1571 27 1586 9973
rect 1510 -2 1586 27
rect 2014 9973 2090 10002
rect 2014 27 2029 9973
rect 2075 27 2090 9973
rect 2014 -2 2090 27
rect 2518 9973 2594 10002
rect 2518 27 2533 9973
rect 2579 27 2594 9973
rect 2518 -2 2594 27
rect 3022 9973 3098 10002
rect 3022 27 3037 9973
rect 3083 27 3098 9973
rect 3022 -2 3098 27
rect 3526 9973 3602 10002
rect 3526 27 3541 9973
rect 3587 27 3602 9973
rect 3526 -2 3602 27
rect 4030 9973 4106 10002
rect 4030 27 4045 9973
rect 4091 27 4106 9973
rect 4030 -2 4106 27
rect 4534 9973 4610 10002
rect 4534 27 4549 9973
rect 4595 27 4610 9973
rect 4534 -2 4610 27
rect 5038 9973 5114 10002
rect 5038 27 5053 9973
rect 5099 27 5114 9973
rect 5038 -2 5114 27
rect 5542 9973 5618 10002
rect 5542 27 5557 9973
rect 5603 27 5618 9973
rect 5542 -2 5618 27
rect 6046 9973 6122 10002
rect 6046 27 6061 9973
rect 6107 27 6122 9973
rect 6046 -2 6122 27
rect 6550 9973 6626 10002
rect 6550 27 6565 9973
rect 6611 27 6626 9973
rect 6550 -2 6626 27
rect 7054 9973 7130 10002
rect 7054 27 7069 9973
rect 7115 27 7130 9973
rect 7054 -2 7130 27
rect 7558 9973 7634 10002
rect 7558 27 7573 9973
rect 7619 27 7634 9973
rect 7558 -2 7634 27
rect 8062 9973 8138 10002
rect 8062 27 8077 9973
rect 8123 27 8138 9973
rect 8062 -2 8138 27
rect 8566 9973 8642 10002
rect 8566 27 8581 9973
rect 8627 27 8642 9973
rect 8566 -2 8642 27
rect 9070 9973 9146 10002
rect 9070 27 9085 9973
rect 9131 27 9146 9973
rect 9070 -2 9146 27
rect 9574 9973 9650 10002
rect 9574 27 9589 9973
rect 9635 27 9650 9973
rect 9574 -2 9650 27
rect 10078 9973 10154 10002
rect 10078 27 10093 9973
rect 10139 27 10154 9973
rect 10078 -2 10154 27
rect 10582 9973 10658 10002
rect 10582 27 10597 9973
rect 10643 27 10658 9973
rect 10582 -2 10658 27
rect 11086 9973 11162 10002
rect 11086 27 11101 9973
rect 11147 27 11162 9973
rect 11086 -2 11162 27
rect 11590 9973 11666 10002
rect 11590 27 11605 9973
rect 11651 27 11666 9973
rect 11590 -2 11666 27
rect 12094 9973 12170 10002
rect 12094 27 12109 9973
rect 12155 27 12170 9973
rect 12094 -2 12170 27
rect 12598 9973 12674 10002
rect 12598 27 12613 9973
rect 12659 27 12674 9973
rect 12598 -2 12674 27
rect 13102 9973 13178 10002
rect 13102 27 13117 9973
rect 13163 27 13178 9973
rect 13102 -2 13178 27
rect 13606 9973 13682 10002
rect 13606 27 13621 9973
rect 13667 27 13682 9973
rect 13606 -2 13682 27
rect 14110 9973 14186 10002
rect 14110 27 14125 9973
rect 14171 27 14186 9973
rect 14110 -2 14186 27
rect 14614 9973 14690 10002
rect 14614 27 14629 9973
rect 14675 27 14690 9973
rect 14614 -2 14690 27
rect 15118 9973 15194 10002
rect 15118 27 15133 9973
rect 15179 27 15194 9973
rect 15118 -2 15194 27
rect 15622 9973 15698 10002
rect 15622 27 15637 9973
rect 15683 27 15698 9973
rect 15622 -2 15698 27
rect 16126 9973 16202 10002
rect 16126 27 16141 9973
rect 16187 27 16202 9973
rect 16126 -2 16202 27
rect 16630 9973 16706 10002
rect 16630 27 16645 9973
rect 16691 27 16706 9973
rect 16630 -2 16706 27
rect 17134 9973 17210 10002
rect 17134 27 17149 9973
rect 17195 27 17210 9973
rect 17134 -2 17210 27
rect 17638 9973 17714 10002
rect 17638 27 17653 9973
rect 17699 27 17714 9973
rect 17638 -2 17714 27
rect 18142 9973 18218 10002
rect 18142 27 18157 9973
rect 18203 27 18218 9973
rect 18142 -2 18218 27
rect 18646 9973 18722 10002
rect 18646 27 18661 9973
rect 18707 27 18722 9973
rect 18646 -2 18722 27
rect 19150 9973 19226 10002
rect 19150 27 19165 9973
rect 19211 27 19226 9973
rect 19150 -2 19226 27
rect 19654 9973 19730 10002
rect 19654 27 19669 9973
rect 19715 27 19730 9973
rect 19654 -2 19730 27
rect 20158 9973 20234 10002
rect 20158 27 20173 9973
rect 20219 27 20234 9973
rect 20158 -2 20234 27
rect 20662 9973 20738 10002
rect 20662 27 20677 9973
rect 20723 27 20738 9973
rect 20662 -2 20738 27
rect 21166 9973 21242 10002
rect 21166 27 21181 9973
rect 21227 27 21242 9973
rect 21166 -2 21242 27
rect 21670 9973 21746 10002
rect 21670 27 21685 9973
rect 21731 27 21746 9973
rect 21670 -2 21746 27
rect 22174 9973 22250 10002
rect 22174 27 22189 9973
rect 22235 27 22250 9973
rect 22174 -2 22250 27
rect 22678 9973 22754 10002
rect 22678 27 22693 9973
rect 22739 27 22754 9973
rect 22678 -2 22754 27
rect 23182 9973 23258 10002
rect 23182 27 23197 9973
rect 23243 27 23258 9973
rect 23182 -2 23258 27
rect 23686 9973 23762 10002
rect 23686 27 23701 9973
rect 23747 27 23762 9973
rect 23686 -2 23762 27
rect 24190 9973 24266 10002
rect 24190 27 24205 9973
rect 24251 27 24266 9973
rect 24190 -2 24266 27
rect 24694 9973 24770 10002
rect 24694 27 24709 9973
rect 24755 27 24770 9973
rect 24694 -2 24770 27
rect 25198 9973 25274 10002
rect 25198 27 25213 9973
rect 25259 27 25274 9973
rect 25198 -2 25274 27
<< end >>
