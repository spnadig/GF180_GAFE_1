*********************************************************************************

** sch_path: /home/lmadhu/openmpw/pdk_1/Project_gf180_tp/xschem/Amplifiers/OTA_2stage.sch

.subckt OTA_2stage vout vin1 vin2 vdd vss vp

*.opin vout

*.ipin vin1

*.ipin vin2

*.iopin vdd

*.iopin vss

*.ipin vp

********************************************************************************

****Differential NMOS Input pairs 
****(multiplicity doesnot work in the model. Multiple NMOS cells (for m=18 and W/L= 100u/1u) should be written manually)

XM1 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM12 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM13 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM14 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM15 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM16 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM17 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM18 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM19 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM110 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM111 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM112 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM113 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM114 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM115 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM116 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM117 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM118 vx vin1 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1

XM2 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM22 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM23 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM24 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM25 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM26 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM27 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM28 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM29 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM210 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM211 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM212 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM213 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM214 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM215 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM216 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM217 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1
XM218 net1 vin2 vtail vss nfet_03v3 L=1u W=100u nf=500 m=1

*****PMOS active load pairs

XM3 vx vx vdd vdd pfet_03v3 L=2u W=50u nf=50 m=1

XM4 net1 vx vdd vdd pfet_03v3 L=2u W=50u nf=50 m=1


*****Tail current NMOS 

XM5 vtail vbias_tail vss vss nfet_03v3 L=1u W=60u nf=60 m=1

*****Current Mirror NMOS 

XM6 vbias_tail vbias_tail vss vss nfet_03v3 L=1u W=20u nf=1 m=1

*****Current Reference PMOS

XM7 vbias_tail vp vdd vdd pfet_03v3 L=2u W=10u nf=1 m=1


*****Second stage Amplifier 

****(multiplicity doesnot work in the model. Multiple NMOS cells (for m=7 and W/L= 100u/1u) should be written manually)

XM8 vout vbias_tail vss vss nfet_03v3 L=1u W=100u nf=1 m=1
XM82 vout vbias_tail vss vss nfet_03v3 L=1u W=100u nf=1 m=1
XM83 vout vbias_tail vss vss nfet_03v3 L=1u W=100u nf=1 m=1
XM84 vout vbias_tail vss vss nfet_03v3 L=1u W=100u nf=1 m=1
XM85 vout vbias_tail vss vss nfet_03v3 L=1u W=100u nf=1 m=1
XM86 vout vbias_tail vss vss nfet_03v3 L=1u W=100u nf=1 m=1
XM87 vout vbias_tail vss vss nfet_03v3 L=1u W=100u nf=1 m=1

****(multiplicity doesnot work in the model. Multiple PMOS cells (for m=4 and W/L= 100u/0.7u) should be written manually)

XM10 vout net1 vdd vdd pfet_03v3 L=0.7u W=100u nf=5 m=1
XM102 vout net1 vdd vdd pfet_03v3 L=0.7u W=100u nf=5 m=1
XM103 vout net1 vdd vdd pfet_03v3 L=0.7u W=100u nf=5 m=1
XM104 vout net1 vdd vdd pfet_03v3 L=0.7u W=100u nf=5 m=1

*****Load Cap
C1 vout GND 1p m=1

*****Miller Compensation cap
C2 net2 vout 3p m=1

R1 net1 net2 200 m=1

.ends

