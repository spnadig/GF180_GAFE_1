magic
tech gf180mcuC
magscale 1 10
timestamp 1676577649
<< error_p >>
rect -66 0 -64 12000
rect 0 0 2 12000
<< nmos >>
rect 88 0 288 12000
rect 392 0 592 12000
rect 696 0 896 12000
rect 1000 0 1200 12000
rect 1304 0 1504 12000
rect 1608 0 1808 12000
rect 1912 0 2112 12000
rect 2216 0 2416 12000
rect 2520 0 2720 12000
rect 2824 0 3024 12000
rect 3128 0 3328 12000
rect 3432 0 3632 12000
rect 3736 0 3936 12000
rect 4040 0 4240 12000
rect 4344 0 4544 12000
rect 4648 0 4848 12000
rect 4952 0 5152 12000
rect 5256 0 5456 12000
rect 5560 0 5760 12000
rect 5864 0 6064 12000
rect 6168 0 6368 12000
rect 6472 0 6672 12000
rect 6776 0 6976 12000
rect 7080 0 7280 12000
rect 7384 0 7584 12000
rect 7688 0 7888 12000
rect 7992 0 8192 12000
rect 8296 0 8496 12000
rect 8600 0 8800 12000
rect 8904 0 9104 12000
rect 9208 0 9408 12000
rect 9512 0 9712 12000
rect 9816 0 10016 12000
rect 10120 0 10320 12000
rect 10424 0 10624 12000
rect 10728 0 10928 12000
rect 11032 0 11232 12000
rect 11336 0 11536 12000
rect 11640 0 11840 12000
rect 11944 0 12144 12000
rect 12248 0 12448 12000
rect 12552 0 12752 12000
rect 12856 0 13056 12000
rect 13160 0 13360 12000
rect 13464 0 13664 12000
rect 13768 0 13968 12000
rect 14072 0 14272 12000
rect 14376 0 14576 12000
rect 14680 0 14880 12000
rect 14984 0 15184 12000
rect 15288 0 15488 12000
rect 15592 0 15792 12000
rect 15896 0 16096 12000
rect 16200 0 16400 12000
rect 16504 0 16704 12000
rect 16808 0 17008 12000
rect 17112 0 17312 12000
rect 17416 0 17616 12000
rect 17720 0 17920 12000
rect 18024 0 18224 12000
<< ndiff >>
rect 0 11973 88 12000
rect 0 27 13 11973
rect 59 27 88 11973
rect 0 0 88 27
rect 288 11973 392 12000
rect 288 27 317 11973
rect 363 27 392 11973
rect 288 0 392 27
rect 592 11973 696 12000
rect 592 27 621 11973
rect 667 27 696 11973
rect 592 0 696 27
rect 896 11973 1000 12000
rect 896 27 925 11973
rect 971 27 1000 11973
rect 896 0 1000 27
rect 1200 11973 1304 12000
rect 1200 27 1229 11973
rect 1275 27 1304 11973
rect 1200 0 1304 27
rect 1504 11973 1608 12000
rect 1504 27 1533 11973
rect 1579 27 1608 11973
rect 1504 0 1608 27
rect 1808 11973 1912 12000
rect 1808 27 1837 11973
rect 1883 27 1912 11973
rect 1808 0 1912 27
rect 2112 11973 2216 12000
rect 2112 27 2141 11973
rect 2187 27 2216 11973
rect 2112 0 2216 27
rect 2416 11973 2520 12000
rect 2416 27 2445 11973
rect 2491 27 2520 11973
rect 2416 0 2520 27
rect 2720 11973 2824 12000
rect 2720 27 2749 11973
rect 2795 27 2824 11973
rect 2720 0 2824 27
rect 3024 11973 3128 12000
rect 3024 27 3053 11973
rect 3099 27 3128 11973
rect 3024 0 3128 27
rect 3328 11973 3432 12000
rect 3328 27 3357 11973
rect 3403 27 3432 11973
rect 3328 0 3432 27
rect 3632 11973 3736 12000
rect 3632 27 3661 11973
rect 3707 27 3736 11973
rect 3632 0 3736 27
rect 3936 11973 4040 12000
rect 3936 27 3965 11973
rect 4011 27 4040 11973
rect 3936 0 4040 27
rect 4240 11973 4344 12000
rect 4240 27 4269 11973
rect 4315 27 4344 11973
rect 4240 0 4344 27
rect 4544 11973 4648 12000
rect 4544 27 4573 11973
rect 4619 27 4648 11973
rect 4544 0 4648 27
rect 4848 11973 4952 12000
rect 4848 27 4877 11973
rect 4923 27 4952 11973
rect 4848 0 4952 27
rect 5152 11973 5256 12000
rect 5152 27 5181 11973
rect 5227 27 5256 11973
rect 5152 0 5256 27
rect 5456 11973 5560 12000
rect 5456 27 5485 11973
rect 5531 27 5560 11973
rect 5456 0 5560 27
rect 5760 11973 5864 12000
rect 5760 27 5789 11973
rect 5835 27 5864 11973
rect 5760 0 5864 27
rect 6064 11973 6168 12000
rect 6064 27 6093 11973
rect 6139 27 6168 11973
rect 6064 0 6168 27
rect 6368 11973 6472 12000
rect 6368 27 6397 11973
rect 6443 27 6472 11973
rect 6368 0 6472 27
rect 6672 11973 6776 12000
rect 6672 27 6701 11973
rect 6747 27 6776 11973
rect 6672 0 6776 27
rect 6976 11973 7080 12000
rect 6976 27 7005 11973
rect 7051 27 7080 11973
rect 6976 0 7080 27
rect 7280 11973 7384 12000
rect 7280 27 7309 11973
rect 7355 27 7384 11973
rect 7280 0 7384 27
rect 7584 11973 7688 12000
rect 7584 27 7613 11973
rect 7659 27 7688 11973
rect 7584 0 7688 27
rect 7888 11973 7992 12000
rect 7888 27 7917 11973
rect 7963 27 7992 11973
rect 7888 0 7992 27
rect 8192 11973 8296 12000
rect 8192 27 8221 11973
rect 8267 27 8296 11973
rect 8192 0 8296 27
rect 8496 11973 8600 12000
rect 8496 27 8525 11973
rect 8571 27 8600 11973
rect 8496 0 8600 27
rect 8800 11973 8904 12000
rect 8800 27 8829 11973
rect 8875 27 8904 11973
rect 8800 0 8904 27
rect 9104 11973 9208 12000
rect 9104 27 9133 11973
rect 9179 27 9208 11973
rect 9104 0 9208 27
rect 9408 11973 9512 12000
rect 9408 27 9437 11973
rect 9483 27 9512 11973
rect 9408 0 9512 27
rect 9712 11973 9816 12000
rect 9712 27 9741 11973
rect 9787 27 9816 11973
rect 9712 0 9816 27
rect 10016 11973 10120 12000
rect 10016 27 10045 11973
rect 10091 27 10120 11973
rect 10016 0 10120 27
rect 10320 11973 10424 12000
rect 10320 27 10349 11973
rect 10395 27 10424 11973
rect 10320 0 10424 27
rect 10624 11973 10728 12000
rect 10624 27 10653 11973
rect 10699 27 10728 11973
rect 10624 0 10728 27
rect 10928 11973 11032 12000
rect 10928 27 10957 11973
rect 11003 27 11032 11973
rect 10928 0 11032 27
rect 11232 11973 11336 12000
rect 11232 27 11261 11973
rect 11307 27 11336 11973
rect 11232 0 11336 27
rect 11536 11973 11640 12000
rect 11536 27 11565 11973
rect 11611 27 11640 11973
rect 11536 0 11640 27
rect 11840 11973 11944 12000
rect 11840 27 11869 11973
rect 11915 27 11944 11973
rect 11840 0 11944 27
rect 12144 11973 12248 12000
rect 12144 27 12173 11973
rect 12219 27 12248 11973
rect 12144 0 12248 27
rect 12448 11973 12552 12000
rect 12448 27 12477 11973
rect 12523 27 12552 11973
rect 12448 0 12552 27
rect 12752 11973 12856 12000
rect 12752 27 12781 11973
rect 12827 27 12856 11973
rect 12752 0 12856 27
rect 13056 11973 13160 12000
rect 13056 27 13085 11973
rect 13131 27 13160 11973
rect 13056 0 13160 27
rect 13360 11973 13464 12000
rect 13360 27 13389 11973
rect 13435 27 13464 11973
rect 13360 0 13464 27
rect 13664 11973 13768 12000
rect 13664 27 13693 11973
rect 13739 27 13768 11973
rect 13664 0 13768 27
rect 13968 11973 14072 12000
rect 13968 27 13997 11973
rect 14043 27 14072 11973
rect 13968 0 14072 27
rect 14272 11973 14376 12000
rect 14272 27 14301 11973
rect 14347 27 14376 11973
rect 14272 0 14376 27
rect 14576 11973 14680 12000
rect 14576 27 14605 11973
rect 14651 27 14680 11973
rect 14576 0 14680 27
rect 14880 11973 14984 12000
rect 14880 27 14909 11973
rect 14955 27 14984 11973
rect 14880 0 14984 27
rect 15184 11973 15288 12000
rect 15184 27 15213 11973
rect 15259 27 15288 11973
rect 15184 0 15288 27
rect 15488 11973 15592 12000
rect 15488 27 15517 11973
rect 15563 27 15592 11973
rect 15488 0 15592 27
rect 15792 11973 15896 12000
rect 15792 27 15821 11973
rect 15867 27 15896 11973
rect 15792 0 15896 27
rect 16096 11973 16200 12000
rect 16096 27 16125 11973
rect 16171 27 16200 11973
rect 16096 0 16200 27
rect 16400 11973 16504 12000
rect 16400 27 16429 11973
rect 16475 27 16504 11973
rect 16400 0 16504 27
rect 16704 11973 16808 12000
rect 16704 27 16733 11973
rect 16779 27 16808 11973
rect 16704 0 16808 27
rect 17008 11973 17112 12000
rect 17008 27 17037 11973
rect 17083 27 17112 11973
rect 17008 0 17112 27
rect 17312 11973 17416 12000
rect 17312 27 17341 11973
rect 17387 27 17416 11973
rect 17312 0 17416 27
rect 17616 11973 17720 12000
rect 17616 27 17645 11973
rect 17691 27 17720 11973
rect 17616 0 17720 27
rect 17920 11973 18024 12000
rect 17920 27 17949 11973
rect 17995 27 18024 11973
rect 17920 0 18024 27
rect 18224 11973 18312 12000
rect 18224 27 18253 11973
rect 18299 27 18312 11973
rect 18224 0 18312 27
<< ndiffc >>
rect 13 27 59 11973
rect 317 27 363 11973
rect 621 27 667 11973
rect 925 27 971 11973
rect 1229 27 1275 11973
rect 1533 27 1579 11973
rect 1837 27 1883 11973
rect 2141 27 2187 11973
rect 2445 27 2491 11973
rect 2749 27 2795 11973
rect 3053 27 3099 11973
rect 3357 27 3403 11973
rect 3661 27 3707 11973
rect 3965 27 4011 11973
rect 4269 27 4315 11973
rect 4573 27 4619 11973
rect 4877 27 4923 11973
rect 5181 27 5227 11973
rect 5485 27 5531 11973
rect 5789 27 5835 11973
rect 6093 27 6139 11973
rect 6397 27 6443 11973
rect 6701 27 6747 11973
rect 7005 27 7051 11973
rect 7309 27 7355 11973
rect 7613 27 7659 11973
rect 7917 27 7963 11973
rect 8221 27 8267 11973
rect 8525 27 8571 11973
rect 8829 27 8875 11973
rect 9133 27 9179 11973
rect 9437 27 9483 11973
rect 9741 27 9787 11973
rect 10045 27 10091 11973
rect 10349 27 10395 11973
rect 10653 27 10699 11973
rect 10957 27 11003 11973
rect 11261 27 11307 11973
rect 11565 27 11611 11973
rect 11869 27 11915 11973
rect 12173 27 12219 11973
rect 12477 27 12523 11973
rect 12781 27 12827 11973
rect 13085 27 13131 11973
rect 13389 27 13435 11973
rect 13693 27 13739 11973
rect 13997 27 14043 11973
rect 14301 27 14347 11973
rect 14605 27 14651 11973
rect 14909 27 14955 11973
rect 15213 27 15259 11973
rect 15517 27 15563 11973
rect 15821 27 15867 11973
rect 16125 27 16171 11973
rect 16429 27 16475 11973
rect 16733 27 16779 11973
rect 17037 27 17083 11973
rect 17341 27 17387 11973
rect 17645 27 17691 11973
rect 17949 27 17995 11973
rect 18253 27 18299 11973
<< psubdiff >>
rect -152 11973 -64 12000
rect -152 27 -131 11973
rect -85 27 -64 11973
rect -152 0 -64 27
<< psubdiffcont >>
rect -131 27 -85 11973
<< polysilicon >>
rect 88 12000 288 12044
rect 392 12000 592 12044
rect 696 12000 896 12044
rect 1000 12000 1200 12044
rect 1304 12000 1504 12044
rect 1608 12000 1808 12044
rect 1912 12000 2112 12044
rect 2216 12000 2416 12044
rect 2520 12000 2720 12044
rect 2824 12000 3024 12044
rect 3128 12000 3328 12044
rect 3432 12000 3632 12044
rect 3736 12000 3936 12044
rect 4040 12000 4240 12044
rect 4344 12000 4544 12044
rect 4648 12000 4848 12044
rect 4952 12000 5152 12044
rect 5256 12000 5456 12044
rect 5560 12000 5760 12044
rect 5864 12000 6064 12044
rect 6168 12000 6368 12044
rect 6472 12000 6672 12044
rect 6776 12000 6976 12044
rect 7080 12000 7280 12044
rect 7384 12000 7584 12044
rect 7688 12000 7888 12044
rect 7992 12000 8192 12044
rect 8296 12000 8496 12044
rect 8600 12000 8800 12044
rect 8904 12000 9104 12044
rect 9208 12000 9408 12044
rect 9512 12000 9712 12044
rect 9816 12000 10016 12044
rect 10120 12000 10320 12044
rect 10424 12000 10624 12044
rect 10728 12000 10928 12044
rect 11032 12000 11232 12044
rect 11336 12000 11536 12044
rect 11640 12000 11840 12044
rect 11944 12000 12144 12044
rect 12248 12000 12448 12044
rect 12552 12000 12752 12044
rect 12856 12000 13056 12044
rect 13160 12000 13360 12044
rect 13464 12000 13664 12044
rect 13768 12000 13968 12044
rect 14072 12000 14272 12044
rect 14376 12000 14576 12044
rect 14680 12000 14880 12044
rect 14984 12000 15184 12044
rect 15288 12000 15488 12044
rect 15592 12000 15792 12044
rect 15896 12000 16096 12044
rect 16200 12000 16400 12044
rect 16504 12000 16704 12044
rect 16808 12000 17008 12044
rect 17112 12000 17312 12044
rect 17416 12000 17616 12044
rect 17720 12000 17920 12044
rect 18024 12000 18224 12044
rect 88 -44 288 0
rect 392 -44 592 0
rect 696 -44 896 0
rect 1000 -44 1200 0
rect 1304 -44 1504 0
rect 1608 -44 1808 0
rect 1912 -44 2112 0
rect 2216 -44 2416 0
rect 2520 -44 2720 0
rect 2824 -44 3024 0
rect 3128 -44 3328 0
rect 3432 -44 3632 0
rect 3736 -44 3936 0
rect 4040 -44 4240 0
rect 4344 -44 4544 0
rect 4648 -44 4848 0
rect 4952 -44 5152 0
rect 5256 -44 5456 0
rect 5560 -44 5760 0
rect 5864 -44 6064 0
rect 6168 -44 6368 0
rect 6472 -44 6672 0
rect 6776 -44 6976 0
rect 7080 -44 7280 0
rect 7384 -44 7584 0
rect 7688 -44 7888 0
rect 7992 -44 8192 0
rect 8296 -44 8496 0
rect 8600 -44 8800 0
rect 8904 -44 9104 0
rect 9208 -44 9408 0
rect 9512 -44 9712 0
rect 9816 -44 10016 0
rect 10120 -44 10320 0
rect 10424 -44 10624 0
rect 10728 -44 10928 0
rect 11032 -44 11232 0
rect 11336 -44 11536 0
rect 11640 -44 11840 0
rect 11944 -44 12144 0
rect 12248 -44 12448 0
rect 12552 -44 12752 0
rect 12856 -44 13056 0
rect 13160 -44 13360 0
rect 13464 -44 13664 0
rect 13768 -44 13968 0
rect 14072 -44 14272 0
rect 14376 -44 14576 0
rect 14680 -44 14880 0
rect 14984 -44 15184 0
rect 15288 -44 15488 0
rect 15592 -44 15792 0
rect 15896 -44 16096 0
rect 16200 -44 16400 0
rect 16504 -44 16704 0
rect 16808 -44 17008 0
rect 17112 -44 17312 0
rect 17416 -44 17616 0
rect 17720 -44 17920 0
rect 18024 -44 18224 0
<< metal1 >>
rect -152 11973 -64 12000
rect -152 27 -131 11973
rect -85 27 -64 11973
rect -152 0 -64 27
rect -2 11973 74 12002
rect -2 27 13 11973
rect 59 27 74 11973
rect -2 -2 74 27
rect 302 11973 378 12002
rect 302 27 317 11973
rect 363 27 378 11973
rect 302 -2 378 27
rect 606 11973 682 12002
rect 606 27 621 11973
rect 667 27 682 11973
rect 606 -2 682 27
rect 910 11973 986 12002
rect 910 27 925 11973
rect 971 27 986 11973
rect 910 -2 986 27
rect 1214 11973 1290 12002
rect 1214 27 1229 11973
rect 1275 27 1290 11973
rect 1214 -2 1290 27
rect 1518 11973 1594 12002
rect 1518 27 1533 11973
rect 1579 27 1594 11973
rect 1518 -2 1594 27
rect 1822 11973 1898 12002
rect 1822 27 1837 11973
rect 1883 27 1898 11973
rect 1822 -2 1898 27
rect 2126 11973 2202 12002
rect 2126 27 2141 11973
rect 2187 27 2202 11973
rect 2126 -2 2202 27
rect 2430 11973 2506 12002
rect 2430 27 2445 11973
rect 2491 27 2506 11973
rect 2430 -2 2506 27
rect 2734 11973 2810 12002
rect 2734 27 2749 11973
rect 2795 27 2810 11973
rect 2734 -2 2810 27
rect 3038 11973 3114 12002
rect 3038 27 3053 11973
rect 3099 27 3114 11973
rect 3038 -2 3114 27
rect 3342 11973 3418 12002
rect 3342 27 3357 11973
rect 3403 27 3418 11973
rect 3342 -2 3418 27
rect 3646 11973 3722 12002
rect 3646 27 3661 11973
rect 3707 27 3722 11973
rect 3646 -2 3722 27
rect 3950 11973 4026 12002
rect 3950 27 3965 11973
rect 4011 27 4026 11973
rect 3950 -2 4026 27
rect 4254 11973 4330 12002
rect 4254 27 4269 11973
rect 4315 27 4330 11973
rect 4254 -2 4330 27
rect 4558 11973 4634 12002
rect 4558 27 4573 11973
rect 4619 27 4634 11973
rect 4558 -2 4634 27
rect 4862 11973 4938 12002
rect 4862 27 4877 11973
rect 4923 27 4938 11973
rect 4862 -2 4938 27
rect 5166 11973 5242 12002
rect 5166 27 5181 11973
rect 5227 27 5242 11973
rect 5166 -2 5242 27
rect 5470 11973 5546 12002
rect 5470 27 5485 11973
rect 5531 27 5546 11973
rect 5470 -2 5546 27
rect 5774 11973 5850 12002
rect 5774 27 5789 11973
rect 5835 27 5850 11973
rect 5774 -2 5850 27
rect 6078 11973 6154 12002
rect 6078 27 6093 11973
rect 6139 27 6154 11973
rect 6078 -2 6154 27
rect 6382 11973 6458 12002
rect 6382 27 6397 11973
rect 6443 27 6458 11973
rect 6382 -2 6458 27
rect 6686 11973 6762 12002
rect 6686 27 6701 11973
rect 6747 27 6762 11973
rect 6686 -2 6762 27
rect 6990 11973 7066 12002
rect 6990 27 7005 11973
rect 7051 27 7066 11973
rect 6990 -2 7066 27
rect 7294 11973 7370 12002
rect 7294 27 7309 11973
rect 7355 27 7370 11973
rect 7294 -2 7370 27
rect 7598 11973 7674 12002
rect 7598 27 7613 11973
rect 7659 27 7674 11973
rect 7598 -2 7674 27
rect 7902 11973 7978 12002
rect 7902 27 7917 11973
rect 7963 27 7978 11973
rect 7902 -2 7978 27
rect 8206 11973 8282 12002
rect 8206 27 8221 11973
rect 8267 27 8282 11973
rect 8206 -2 8282 27
rect 8510 11973 8586 12002
rect 8510 27 8525 11973
rect 8571 27 8586 11973
rect 8510 -2 8586 27
rect 8814 11973 8890 12002
rect 8814 27 8829 11973
rect 8875 27 8890 11973
rect 8814 -2 8890 27
rect 9118 11973 9194 12002
rect 9118 27 9133 11973
rect 9179 27 9194 11973
rect 9118 -2 9194 27
rect 9422 11973 9498 12002
rect 9422 27 9437 11973
rect 9483 27 9498 11973
rect 9422 -2 9498 27
rect 9726 11973 9802 12002
rect 9726 27 9741 11973
rect 9787 27 9802 11973
rect 9726 -2 9802 27
rect 10030 11973 10106 12002
rect 10030 27 10045 11973
rect 10091 27 10106 11973
rect 10030 -2 10106 27
rect 10334 11973 10410 12002
rect 10334 27 10349 11973
rect 10395 27 10410 11973
rect 10334 -2 10410 27
rect 10638 11973 10714 12002
rect 10638 27 10653 11973
rect 10699 27 10714 11973
rect 10638 -2 10714 27
rect 10942 11973 11018 12002
rect 10942 27 10957 11973
rect 11003 27 11018 11973
rect 10942 -2 11018 27
rect 11246 11973 11322 12002
rect 11246 27 11261 11973
rect 11307 27 11322 11973
rect 11246 -2 11322 27
rect 11550 11973 11626 12002
rect 11550 27 11565 11973
rect 11611 27 11626 11973
rect 11550 -2 11626 27
rect 11854 11973 11930 12002
rect 11854 27 11869 11973
rect 11915 27 11930 11973
rect 11854 -2 11930 27
rect 12158 11973 12234 12002
rect 12158 27 12173 11973
rect 12219 27 12234 11973
rect 12158 -2 12234 27
rect 12462 11973 12538 12002
rect 12462 27 12477 11973
rect 12523 27 12538 11973
rect 12462 -2 12538 27
rect 12766 11973 12842 12002
rect 12766 27 12781 11973
rect 12827 27 12842 11973
rect 12766 -2 12842 27
rect 13070 11973 13146 12002
rect 13070 27 13085 11973
rect 13131 27 13146 11973
rect 13070 -2 13146 27
rect 13374 11973 13450 12002
rect 13374 27 13389 11973
rect 13435 27 13450 11973
rect 13374 -2 13450 27
rect 13678 11973 13754 12002
rect 13678 27 13693 11973
rect 13739 27 13754 11973
rect 13678 -2 13754 27
rect 13982 11973 14058 12002
rect 13982 27 13997 11973
rect 14043 27 14058 11973
rect 13982 -2 14058 27
rect 14286 11973 14362 12002
rect 14286 27 14301 11973
rect 14347 27 14362 11973
rect 14286 -2 14362 27
rect 14590 11973 14666 12002
rect 14590 27 14605 11973
rect 14651 27 14666 11973
rect 14590 -2 14666 27
rect 14894 11973 14970 12002
rect 14894 27 14909 11973
rect 14955 27 14970 11973
rect 14894 -2 14970 27
rect 15198 11973 15274 12002
rect 15198 27 15213 11973
rect 15259 27 15274 11973
rect 15198 -2 15274 27
rect 15502 11973 15578 12002
rect 15502 27 15517 11973
rect 15563 27 15578 11973
rect 15502 -2 15578 27
rect 15806 11973 15882 12002
rect 15806 27 15821 11973
rect 15867 27 15882 11973
rect 15806 -2 15882 27
rect 16110 11973 16186 12002
rect 16110 27 16125 11973
rect 16171 27 16186 11973
rect 16110 -2 16186 27
rect 16414 11973 16490 12002
rect 16414 27 16429 11973
rect 16475 27 16490 11973
rect 16414 -2 16490 27
rect 16718 11973 16794 12002
rect 16718 27 16733 11973
rect 16779 27 16794 11973
rect 16718 -2 16794 27
rect 17022 11973 17098 12002
rect 17022 27 17037 11973
rect 17083 27 17098 11973
rect 17022 -2 17098 27
rect 17326 11973 17402 12002
rect 17326 27 17341 11973
rect 17387 27 17402 11973
rect 17326 -2 17402 27
rect 17630 11973 17706 12002
rect 17630 27 17645 11973
rect 17691 27 17706 11973
rect 17630 -2 17706 27
rect 17934 11973 18010 12002
rect 17934 27 17949 11973
rect 17995 27 18010 11973
rect 17934 -2 18010 27
rect 18238 11973 18314 12002
rect 18238 27 18253 11973
rect 18299 27 18314 11973
rect 18238 -2 18314 27
<< end >>
