VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO TopLevel_oscillator_macro
  CLASS BLOCK ;
  FOREIGN TopLevel_oscillator_macro ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 570.000 ;
  PIN VP
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 284.715 528.845 330.490 559.750 ;
    END
  END VP
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 371.565 528.845 417.340 559.750 ;
    END
  END GND
  PIN ASIG5V
    PORT
      LAYER Metal5 ;
        RECT -112.600 123.490 -112.590 123.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -27.600 123.490 -27.590 123.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 14.480 123.085 89.480 123.515 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 99.480 123.085 174.480 123.515 ;
    END
  END ASIG5V
  PIN CLK_EN
    PORT
      LAYER Metal2 ;
        RECT 29.560 528.845 75.335 559.750 ;
    END
  END CLK_EN
  PIN AND_OUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.860 528.845 160.635 559.750 ;
    END
  END AND_OUT
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.445 528.845 245.220 559.750 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 14.320 78.310 429.640 429.980 ;
      LAYER Metal2 ;
        RECT 14.480 528.545 29.260 529.365 ;
        RECT 75.635 528.545 114.560 529.365 ;
        RECT 160.935 528.545 199.145 529.365 ;
        RECT 245.520 528.545 429.480 529.365 ;
        RECT 14.480 12.770 429.480 528.545 ;
      LAYER Metal3 ;
        RECT 14.480 12.770 429.480 529.365 ;
      LAYER Metal4 ;
        RECT 14.480 528.545 284.415 529.365 ;
        RECT 330.790 528.545 371.265 529.365 ;
        RECT 417.640 528.545 429.480 529.365 ;
        RECT 14.480 12.770 429.480 528.545 ;
      LAYER Metal5 ;
        RECT 14.480 124.015 429.480 529.365 ;
        RECT 89.980 122.585 98.980 124.015 ;
        RECT 174.980 122.585 429.480 124.015 ;
        RECT 14.480 12.770 429.480 122.585 ;
  END
END TopLevel_oscillator_macro
END LIBRARY

