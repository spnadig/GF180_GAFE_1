(*blackbox*)
module OTA_2stage_macro (
    inout vdd,
    inout vss,
    output vout,
    input vin1,
    input vin2,
    input vp
);
endmodule // OTA_2stage
