VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OTA_2stage_macro
  CLASS BLOCK ;
  FOREIGN OTA_2stage_macro ;
  ORIGIN 0.000 0.000 ;
  SIZE 1804.180 BY 1218.995 ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 106.565 349.955 187.040 409.555 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 45.090 628.080 109.565 720.005 ;
    END
  END vdd
  OBS
      LAYER Metal1 ;
        RECT 10.530 720.305 1782.660 1153.455 ;
        RECT 10.530 627.780 44.790 720.305 ;
        RECT 109.865 627.780 1782.660 720.305 ;
        RECT 10.530 409.855 1782.660 627.780 ;
        RECT 10.530 349.655 106.265 409.855 ;
        RECT 187.340 349.655 1782.660 409.855 ;
        RECT 10.530 3.905 1782.660 349.655 ;
      LAYER Metal2 ;
        RECT 10.690 32.950 1695.285 1218.995 ;
      LAYER Metal3 ;
        RECT 10.690 112.505 1732.275 1218.995 ;
      LAYER Metal4 ;
        RECT 10.690 112.505 1799.790 1218.995 ;
      LAYER Metal5 ;
        RECT 10.690 112.505 1798.240 1218.995 ;
  END
END OTA_2stage_macro
END LIBRARY

