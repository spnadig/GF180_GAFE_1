* SPICE3 file created from OTA_2stage.ext - technology: gf180mcuC

.subckt pfet a_3112_n44# a_14200_n44# a_4624_n44# a_15712_n44# a_10064_0# a_18128_0#
+ a_11072_0# a_19136_0# a_6136_n44# a_17224_n44# a_12080_0# a_7648_n44# a_18736_n44#
+ a_2504_0# a_9160_n44# a_3512_0# w_n176_n86# a_10672_n44# a_4520_0# a_20752_n44#
+ a_12184_n44# a_1096_n44# a_992_0# a_13696_n44# a_10568_0# a_3008_0# a_22264_n44#
+ a_4016_0# a_11576_0# a_23776_n44# a_12584_0# a_5024_0# a_13592_0# a_6032_0# a_488_0#
+ a_7040_0# a_2104_n44# a_3616_n44# a_14704_n44# a_6640_n44# a_5128_n44# a_16216_n44#
+ a_13088_0# a_17728_n44# a_19240_n44# a_14096_0# a_8152_n44# a_9664_n44# a_5528_0#
+ a_6536_0# a_7544_0# a_11176_n44# a_8552_0# a_12688_n44# a_9560_0# a_14600_0# a_20144_0#
+ a_21256_n44# a_22768_n44# a_21152_0# a_24280_n44# a_22160_0# a_8048_0# a_9056_0#
+ a_2608_n44# a_88_n44# a_4120_n44# a_15104_0# a_5632_n44# a_16720_n44# a_16112_0#
+ a_15208_n44# a_17120_0# a_20648_0# a_7144_n44# a_18232_n44# a_8656_n44# a_19744_n44#
+ a_21656_0# a_22664_0# a_11680_n44# a_0_0# a_23672_0# a_24680_0# a_1496_0# a_10168_n44#
+ a_21760_n44# a_592_n44# a_13192_n44# a_15608_0# a_20248_n44# a_16616_0# a_23272_n44#
+ a_2000_0# a_17624_0# a_23168_0# a_24784_n44# a_18632_0# a_24176_0# a_1600_n44# a_19640_0#
+ VSUBS a_25184_0#
X0 a_8552_0# a_8152_n44# a_8048_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X1 a_10064_0# a_9664_n44# a_9560_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X2 a_15104_0# a_14704_n44# a_14600_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X3 a_5528_0# a_5128_n44# a_5024_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X4 a_7040_0# a_6640_n44# a_6536_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X5 a_2504_0# a_2104_n44# a_2000_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X6 a_4016_0# a_3616_n44# a_3512_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X7 a_22664_0# a_22264_n44# a_22160_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X8 a_24176_0# a_23776_n44# a_23672_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X9 a_14096_0# a_13696_n44# a_13592_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X10 a_12584_0# a_12184_n44# a_12080_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X11 a_21152_0# a_20752_n44# a_20648_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X12 a_11072_0# a_10672_n44# a_10568_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X13 a_1496_0# a_1096_n44# a_992_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X14 a_19136_0# a_18736_n44# a_18632_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X15 a_17624_0# a_17224_n44# a_17120_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X16 a_16112_0# a_15712_n44# a_15608_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X17 a_6536_0# a_6136_n44# a_6032_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X18 a_8048_0# a_7648_n44# a_7544_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X19 a_9560_0# a_9160_n44# a_9056_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X20 a_14600_0# a_14200_n44# a_14096_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X21 a_5024_0# a_4624_n44# a_4520_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X22 a_25184_0# a_24784_n44# a_24680_0# w_n176_n86# pfet_03v3 ad=22p pd=100.88u as=13p ps=50.52u w=50u l=2u
X23 a_3512_0# a_3112_n44# a_3008_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X24 a_20648_0# a_20248_n44# a_20144_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X25 a_23672_0# a_23272_n44# a_23168_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X26 a_2000_0# a_1600_n44# a_1496_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X27 a_13592_0# a_13192_n44# a_13088_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X28 a_10568_0# a_10168_n44# a_10064_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X29 a_22160_0# a_21760_n44# a_21656_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X30 a_12080_0# a_11680_n44# a_11576_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X31 a_20144_0# a_19744_n44# a_19640_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X32 a_18632_0# a_18232_n44# a_18128_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X33 a_488_0# a_88_n44# a_0_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=22p ps=100.88u w=50u l=2u
X34 a_15608_0# a_15208_n44# a_15104_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X35 a_9056_0# a_8656_n44# a_8552_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X36 a_17120_0# a_16720_n44# a_16616_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X37 a_7544_0# a_7144_n44# a_7040_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X38 a_6032_0# a_5632_n44# a_5528_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X39 a_3008_0# a_2608_n44# a_2504_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X40 a_4520_0# a_4120_n44# a_4016_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X41 a_23168_0# a_22768_n44# a_22664_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X42 a_24680_0# a_24280_n44# a_24176_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X43 a_21656_0# a_21256_n44# a_21152_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X44 a_13088_0# a_12688_n44# a_12584_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X45 a_11576_0# a_11176_n44# a_11072_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X46 a_992_0# a_592_n44# a_488_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X47 a_19640_0# a_19240_n44# a_19136_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X48 a_16616_0# a_16216_n44# a_16112_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
X49 a_18128_0# a_17728_n44# a_17624_0# w_n176_n86# pfet_03v3 ad=13p pd=50.52u as=13p ps=50.52u w=50u l=2u
C0 w_n176_n86# a_0_0# 4.68fF
C1 w_n176_n86# VSUBS 780.45fF
.ends

.subckt nfet$2 a_29776_0# a_592_0# a_15792_0# a_27752_n44# a_23800_n44# a_4952_n44#
+ a_27648_0# a_13664_0# a_20960_0# a_16400_0# a_11536_0# a_15288_n44# a_11336_n44#
+ a_1000_n44# a_5760_0# a_3632_0# a_21368_n44# a_18632_n44# a_28560_0# a_1504_0# a_23696_0#
+ a_28664_n44# a_24712_n44# a_5864_n44# a_1912_n44# a_19136_0# a_26432_0# a_22280_n44#
+ a_8496_0# a_21568_0# a_24304_0# a_10320_0# a_17008_0# a_6368_0# a_12248_n44# a_9104_0#
+ a_19544_n44# a_29168_0# a_15184_0# a_22480_0# a_13160_n44# a_29576_n44# a_25624_n44#
+ a_6776_n44# a_2824_n44# a_7280_0# a_13056_0# a_20352_0# a_23192_n44# a_5152_0# a_9208_n44#
+ a_17920_0# a_3024_0# a_n152_0# a_16504_n44# a_392_n44# a_23088_0# a_30384_0# a_14072_n44#
+ a_10120_n44# a_10928_0# a_26536_n44# a_7688_n44# a_3736_n44# a_20152_n44# a_27952_0#
+ a_30184_n44# a_14984_n44# a_18528_0# a_25824_0# a_11840_0# a_7888_0# a_17416_n44#
+ a_11032_n44# a_27448_n44# a_4648_n44# a_19440_0# a_21064_n44# a_14576_0# a_21872_0#
+ a_17312_0# a_28360_n44# a_15896_n44# a_11944_n44# a_5560_n44# a_6672_0# a_12448_0#
+ a_21976_n44# a_18328_n44# a_4544_0# a_29472_0# a_2416_0# a_24408_n44# a_1608_n44#
+ a_27344_0# a_19240_n44# a_13360_0# a_8904_n44# a_25216_0# a_29272_n44# a_11232_0#
+ a_25320_n44# a_12856_n44# a_6472_n44# a_2520_n44# a_22888_n44# a_16096_0# a_23392_0#
+ a_1200_0# a_8192_0# a_21264_0# a_16200_n44# a_24000_0# a_9816_n44# a_896_0# a_6064_0#
+ a_26232_n44# a_13768_n44# a_7384_n44# a_3432_n44# a_18832_0# a_13968_0# a_16704_0#
+ a_14680_n44# a_8800_0# a_20760_n44# a_17112_n44# a_3936_0# a_28864_0# a_1808_0#
+ a_14880_0# a_27144_n44# a_10728_n44# a_8296_n44# a_4344_n44# a_26736_0# a_12752_0#
+ a_24608_0# a_30080_0# a_10624_0# a_15592_n44# a_11640_n44# a_88_n44# a_9408_0# a_2720_0#
+ a_21672_n44# a_18024_n44# a_288_0# a_22784_0# a_15488_0# a_25520_0# a_28056_n44#
+ a_18224_0# a_24104_n44# a_5256_n44# a_1304_n44# a_7584_0# a_20656_0# a_18936_n44#
+ a_8600_n44# a_5456_0# a_12552_n44# a_28968_n44# a_3328_0# a_22584_n44# a_28256_0#
+ a_14272_0# a_26128_0# a_29880_n44# a_12144_0# a_0_0# a_25016_n44# a_6168_n44# a_2216_n44#
+ a_19848_n44# a_4240_0# a_10016_0# a_9512_n44# a_13464_n44# a_7080_n44# a_2112_0#
+ a_25928_n44# a_27040_0# a_23496_n44# a_22176_0# a_7992_n44# a_20048_0# a_26840_n44#
+ a_3128_n44# a_19744_0# a_16808_n44# a_696_n44# a_17616_0# a_24912_0# a_14376_n44#
+ a_10424_n44# a_4040_n44# a_6976_0# a_9712_0# a_20456_n44# a_17720_n44# a_4848_0#
X0 a_27648_0# a_27448_n44# a_27344_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X1 a_1808_0# a_1608_n44# a_1504_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X2 a_11232_0# a_11032_n44# a_10928_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X3 a_17616_0# a_17416_n44# a_17312_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X4 a_5760_0# a_5560_n44# a_5456_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X5 a_30384_0# a_30184_n44# a_30080_0# a_n152_0# nfet_03v3 ad=44p pd=200.88u as=26p ps=100.52u w=100u l=1000n
X6 a_15184_0# a_14984_n44# a_14880_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X7 a_20352_0# a_20152_n44# a_20048_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X8 a_26736_0# a_26536_n44# a_26432_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X9 a_4848_0# a_4648_n44# a_4544_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X10 a_10320_0# a_10120_n44# a_10016_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X11 a_14272_0# a_14072_n44# a_13968_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X12 a_16704_0# a_16504_n44# a_16400_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X13 a_23392_0# a_23192_n44# a_23088_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X14 a_3936_0# a_3736_n44# a_3632_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X15 a_29776_0# a_29576_n44# a_29472_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X16 a_25824_0# a_25624_n44# a_25520_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X17 a_7888_0# a_7688_n44# a_7584_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X18 a_13360_0# a_13160_n44# a_13056_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X19 a_19744_0# a_19544_n44# a_19440_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X20 a_12448_0# a_12248_n44# a_12144_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X21 a_9408_0# a_9208_n44# a_9104_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X22 a_22480_0# a_22280_n44# a_22176_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X23 a_3024_0# a_2824_n44# a_2720_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X24 a_28864_0# a_28664_n44# a_28560_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X25 a_24912_0# a_24712_n44# a_24608_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X26 a_6976_0# a_6776_n44# a_6672_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X27 a_21568_0# a_21368_n44# a_21264_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X28 a_18832_0# a_18632_n44# a_18528_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X29 a_15488_0# a_15288_n44# a_15184_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X30 a_11536_0# a_11336_n44# a_11232_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X31 a_27952_0# a_27752_n44# a_27648_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X32 a_24000_0# a_23800_n44# a_23696_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X33 a_6064_0# a_5864_n44# a_5760_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X34 a_2112_0# a_1912_n44# a_1808_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X35 a_20656_0# a_20456_n44# a_20352_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X36 a_17920_0# a_17720_n44# a_17616_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X37 a_1200_0# a_1000_n44# a_896_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X38 a_14576_0# a_14376_n44# a_14272_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X39 a_10624_0# a_10424_n44# a_10320_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X40 a_17008_0# a_16808_n44# a_16704_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X41 a_27040_0# a_26840_n44# a_26736_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X42 a_5152_0# a_4952_n44# a_4848_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X43 a_23696_0# a_23496_n44# a_23392_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X44 a_26128_0# a_25928_n44# a_25824_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X45 a_4240_0# a_4040_n44# a_3936_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X46 a_13664_0# a_13464_n44# a_13360_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X47 a_20048_0# a_19848_n44# a_19744_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X48 a_25216_0# a_25016_n44# a_24912_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X49 a_3328_0# a_3128_n44# a_3024_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X50 a_592_0# a_392_n44# a_288_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X51 a_30080_0# a_29880_n44# a_29776_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X52 a_8192_0# a_7992_n44# a_7888_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X53 a_22784_0# a_22584_n44# a_22480_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X54 a_29168_0# a_28968_n44# a_28864_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X55 a_12752_0# a_12552_n44# a_12448_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X56 a_7280_0# a_7080_n44# a_6976_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X57 a_9712_0# a_9512_n44# a_9408_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X58 a_19136_0# a_18936_n44# a_18832_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X59 a_24304_0# a_24104_n44# a_24000_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X60 a_6368_0# a_6168_n44# a_6064_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X61 a_2416_0# a_2216_n44# a_2112_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X62 a_288_0# a_88_n44# a_0_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=44p ps=200.88u w=100u l=1000n
X63 a_28256_0# a_28056_n44# a_27952_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X64 a_21872_0# a_21672_n44# a_21568_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X65 a_18224_0# a_18024_n44# a_17920_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X66 a_15792_0# a_15592_n44# a_15488_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X67 a_11840_0# a_11640_n44# a_11536_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X68 a_8800_0# a_8600_n44# a_8496_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X69 a_1504_0# a_1304_n44# a_1200_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X70 a_27344_0# a_27144_n44# a_27040_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X71 a_10928_0# a_10728_n44# a_10624_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X72 a_5456_0# a_5256_n44# a_5152_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X73 a_20960_0# a_20760_n44# a_20656_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X74 a_17312_0# a_17112_n44# a_17008_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X75 a_14880_0# a_14680_n44# a_14576_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X76 a_26432_0# a_26232_n44# a_26128_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X77 a_13968_0# a_13768_n44# a_13664_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X78 a_8496_0# a_8296_n44# a_8192_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X79 a_4544_0# a_4344_n44# a_4240_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X80 a_16400_0# a_16200_n44# a_16096_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X81 a_896_0# a_696_n44# a_592_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X82 a_23088_0# a_22888_n44# a_22784_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X83 a_25520_0# a_25320_n44# a_25216_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X84 a_13056_0# a_12856_n44# a_12752_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X85 a_7584_0# a_7384_n44# a_7280_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X86 a_3632_0# a_3432_n44# a_3328_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X87 a_29472_0# a_29272_n44# a_29168_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X88 a_10016_0# a_9816_n44# a_9712_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X89 a_19440_0# a_19240_n44# a_19136_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X90 a_24608_0# a_24408_n44# a_24304_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X91 a_22176_0# a_21976_n44# a_21872_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X92 a_18528_0# a_18328_n44# a_18224_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X93 a_12144_0# a_11944_n44# a_11840_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X94 a_6672_0# a_6472_n44# a_6368_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X95 a_2720_0# a_2520_n44# a_2416_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X96 a_28560_0# a_28360_n44# a_28256_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X97 a_16096_0# a_15896_n44# a_15792_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X98 a_9104_0# a_8904_n44# a_8800_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
X99 a_21264_0# a_21064_n44# a_20960_0# a_n152_0# nfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=1000n
C0 a_0_0# a_n152_0# 9.38fF
.ends

.subckt pfet$4 a_8036_0# a_23408_0# a_19852_n44# a_332_n44# a_4376_0# a_17308_0# a_13648_0#
+ a_576_n44# a_12184_0# a_472_0# a_19608_n44# a_18632_n44# a_24140_0# a_18876_n44#
+ a_6572_0# a_19504_0# a_21944_0# a_15844_0# a_18040_0# a_20480_0# a_17412_n44# a_14380_0#
+ a_17656_n44# a_16680_n44# a_16436_n44# a_15460_n44# w_n176_n86# a_1204_0# a_7548_0#
+ a_6084_0# a_19016_0# a_21456_0# a_15216_n44# a_14240_n44# a_3888_0# a_15356_0# a_23512_n44#
+ a_14484_n44# a_11800_n44# a_11696_0# a_3400_0# a_13020_n44# a_9744_0# a_23756_n44#
+ a_22780_n44# a_8280_0# a_23652_0# a_13264_n44# a_17552_0# a_22536_n44# a_21560_n44#
+ a_13892_0# a_10824_n44# a_12044_n44# a_9604_n44# a_21316_n44# a_20340_n44# a_12288_n44#
+ a_9848_n44# a_8872_n44# a_20584_n44# a_9256_0# a_11068_n44# a_10092_n44# a_18528_0#
+ a_20968_0# a_23164_0# a_8628_n44# a_7652_n44# a_5596_0# a_17064_0# a_14868_0# a_7896_n44#
+ a_7408_n44# a_6432_n44# a_2912_0# a_10720_0# a_6676_n44# a_7792_0# a_19260_0# a_5212_n44#
+ a_5456_n44# a_4480_n44# a_4236_n44# a_3260_n44# a_2424_0# a_8768_0# a_10232_0# a_22676_0#
+ a_3016_n44# a_2040_n44# a_16576_0# a_2284_n44# a_4620_0# a_820_n44# a_18772_0# a_1064_n44#
+ a_11208_0# a_22188_0# a_16088_0# a_17900_n44# a_4132_0# a_19120_n44# a_1936_0# a_13404_0#
+ a_19748_0# a_24384_0# a_18284_0# a_19364_n44# a_16924_n44# a_21700_0# a_15600_0#
+ a_18144_n44# a_11940_0# a_18388_n44# a_15704_n44# a_5108_0# a_1448_0# a_15948_n44#
+ a_14972_n44# a_17168_n44# a_16192_n44# a_14728_n44# a_13752_n44# a_7304_0# a_21212_0#
+ a_24000_n44# a_2180_0# a_3644_0# a_12916_0# a_15112_0# a_13996_n44# a_88_n44# a_9988_0#
+ a_11452_0# a_23896_0# a_24244_n44# a_13508_n44# a_12532_n44# a_17796_0# a_9500_0#
+ a_21804_n44# a_12776_n44# a_5840_0# a_23024_n44# a_11312_n44# a_23268_n44# a_22292_n44#
+ a_10580_n44# a_19992_0# a_11556_n44# a_9360_n44# a_3156_0# a_20828_n44# a_12428_0#
+ a_22048_n44# a_21072_n44# a_10336_n44# a_716_0# a_6920_n44# a_9116_n44# a_8140_n44#
+ a_6816_0# a_9012_0# a_5352_0# a_20724_0# a_8384_n44# a_5700_n44# a_14624_0# a_0_0#
+ a_20096_n44# a_1692_0# a_13160_0# a_5944_n44# a_10964_0# a_7164_n44# a_22920_0#
+ a_4724_n44# a_16820_0# a_228_0# a_4968_n44# a_3992_n44# a_6328_0# a_6188_n44# a_3504_n44#
+ a_20236_0# a_2668_0# a_14136_0# a_3748_n44# a_2772_n44# a_10476_0# a_8524_0# a_2528_n44#
+ a_1552_n44# a_7060_0# a_22432_0# a_4864_0# a_16332_0# a_12672_0# a_1796_n44# a_1308_n44#
+ VSUBS a_960_0#
X0 a_2424_0# a_2284_n44# a_2180_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X1 a_3156_0# a_3016_n44# a_2912_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X2 a_2180_0# a_2040_n44# a_1936_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X3 a_4376_0# a_4236_n44# a_4132_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X4 a_3400_0# a_3260_n44# a_3156_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X5 a_11208_0# a_11068_n44# a_10964_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X6 a_10232_0# a_10092_n44# a_9988_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X7 a_5596_0# a_5456_n44# a_5352_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X8 a_4620_0# a_4480_n44# a_4376_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X9 a_20724_0# a_20584_n44# a_20480_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X10 a_5352_0# a_5212_n44# a_5108_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X11 a_21456_0# a_21316_n44# a_21212_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X12 a_20480_0# a_20340_n44# a_20236_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X13 a_12428_0# a_12288_n44# a_12184_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X14 a_6816_0# a_6676_n44# a_6572_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X15 a_12184_0# a_12044_n44# a_11940_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X16 a_7548_0# a_7408_n44# a_7304_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X17 a_6572_0# a_6432_n44# a_6328_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X18 a_22676_0# a_22536_n44# a_22432_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X19 a_21700_0# a_21560_n44# a_21456_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X20 a_10964_0# a_10824_n44# a_10720_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X21 a_8036_0# a_7896_n44# a_7792_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X22 a_13404_0# a_13264_n44# a_13160_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X23 a_8768_0# a_8628_n44# a_8524_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X24 a_7792_0# a_7652_n44# a_7548_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X25 a_23896_0# a_23756_n44# a_23652_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X26 a_22920_0# a_22780_n44# a_22676_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X27 a_13160_0# a_13020_n44# a_12916_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X28 a_23652_0# a_23512_n44# a_23408_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X29 a_14624_0# a_14484_n44# a_14380_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X30 a_11940_0# a_11800_n44# a_11696_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X31 a_9988_0# a_9848_n44# a_9744_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X32 a_9012_0# a_8872_n44# a_8768_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X33 a_15356_0# a_15216_n44# a_15112_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X34 a_14380_0# a_14240_n44# a_14136_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X35 a_9744_0# a_9604_n44# a_9500_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X36 a_16576_0# a_16436_n44# a_16332_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X37 a_15600_0# a_15460_n44# a_15356_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X38 a_17796_0# a_17656_n44# a_17552_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X39 a_16820_0# a_16680_n44# a_16576_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X40 a_17552_0# a_17412_n44# a_17308_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X41 a_19016_0# a_18876_n44# a_18772_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X42 a_960_0# a_820_n44# a_716_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X43 a_19748_0# a_19608_n44# a_19504_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X44 a_18772_0# a_18632_n44# a_18528_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X45 a_19992_0# a_19852_n44# a_19748_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X46 a_1448_0# a_1308_n44# a_1204_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X47 a_1936_0# a_1796_n44# a_1692_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X48 a_2668_0# a_2528_n44# a_2424_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X49 a_1692_0# a_1552_n44# a_1448_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X50 a_20236_0# a_20096_n44# a_19992_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X51 a_3888_0# a_3748_n44# a_3644_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X52 a_2912_0# a_2772_n44# a_2668_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X53 a_6328_0# a_6188_n44# a_6084_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X54 a_3644_0# a_3504_n44# a_3400_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X55 a_5108_0# a_4968_n44# a_4864_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X56 a_4132_0# a_3992_n44# a_3888_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X57 a_22188_0# a_22048_n44# a_21944_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X58 a_21212_0# a_21072_n44# a_20968_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X59 a_10476_0# a_10336_n44# a_10232_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X60 a_4864_0# a_4724_n44# a_4620_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X61 a_20968_0# a_20828_n44# a_20724_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X62 a_7304_0# a_7164_n44# a_7060_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X63 a_23408_0# a_23268_n44# a_23164_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X64 a_22432_0# a_22292_n44# a_22188_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X65 a_11696_0# a_11556_n44# a_11452_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X66 a_10720_0# a_10580_n44# a_10476_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X67 a_6084_0# a_5944_n44# a_5840_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X68 a_228_0# a_88_n44# a_0_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=44p ps=200.88u w=100u l=700n
X69 a_23164_0# a_23024_n44# a_22920_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X70 a_11452_0# a_11312_n44# a_11208_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X71 a_8524_0# a_8384_n44# a_8280_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X72 a_5840_0# a_5700_n44# a_5596_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X73 a_21944_0# a_21804_n44# a_21700_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X74 a_12916_0# a_12776_n44# a_12672_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X75 a_9256_0# a_9116_n44# a_9012_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X76 a_24384_0# a_24244_n44# a_24140_0# w_n176_n86# pfet_03v3 ad=44p pd=200.88u as=26p ps=100.52u w=100u l=700n
X77 a_13648_0# a_13508_n44# a_13404_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X78 a_12672_0# a_12532_n44# a_12428_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X79 a_8280_0# a_8140_n44# a_8036_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X80 a_7060_0# a_6920_n44# a_6816_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X81 a_14136_0# a_13996_n44# a_13892_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X82 a_24140_0# a_24000_n44# a_23896_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X83 a_9500_0# a_9360_n44# a_9256_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X84 a_14868_0# a_14728_n44# a_14624_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X85 a_13892_0# a_13752_n44# a_13648_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X86 a_17308_0# a_17168_n44# a_17064_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X87 a_16332_0# a_16192_n44# a_16088_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X88 a_16088_0# a_15948_n44# a_15844_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X89 a_15112_0# a_14972_n44# a_14868_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X90 a_716_0# a_576_n44# a_472_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X91 a_18528_0# a_18388_n44# a_18284_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X92 a_15844_0# a_15704_n44# a_15600_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X93 a_472_0# a_332_n44# a_228_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X94 a_18284_0# a_18144_n44# a_18040_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X95 a_17064_0# a_16924_n44# a_16820_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X96 a_19504_0# a_19364_n44# a_19260_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X97 a_19260_0# a_19120_n44# a_19016_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X98 a_18040_0# a_17900_n44# a_17796_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
X99 a_1204_0# a_1064_n44# a_960_0# w_n176_n86# pfet_03v3 ad=26p pd=100.52u as=26p ps=100.52u w=100u l=700n
C0 a_19748_0# a_19992_0# 3.49fF
C1 a_16332_0# a_16088_0# 3.49fF
C2 a_2180_0# a_1936_0# 3.49fF
C3 a_2180_0# a_2424_0# 3.49fF
C4 a_18528_0# a_18772_0# 3.49fF
C5 a_8036_0# a_8280_0# 3.49fF
C6 a_3644_0# a_3400_0# 3.49fF
C7 a_2424_0# a_2668_0# 3.49fF
C8 a_19260_0# a_19016_0# 3.49fF
C9 a_22432_0# a_22676_0# 3.49fF
C10 a_12672_0# a_12916_0# 3.49fF
C11 a_8280_0# a_8524_0# 3.49fF
C12 a_15844_0# a_16088_0# 3.49fF
C13 a_17796_0# a_18040_0# 3.49fF
C14 a_9744_0# a_9500_0# 3.49fF
C15 a_228_0# a_0_0# 3.49fF
C16 a_22676_0# a_22920_0# 3.49fF
C17 a_10476_0# a_10720_0# 3.49fF
C18 a_5840_0# a_5596_0# 3.49fF
C19 a_20968_0# a_21212_0# 3.49fF
C20 a_6572_0# a_6328_0# 3.49fF
C21 a_5840_0# a_6084_0# 3.49fF
C22 a_14380_0# a_14624_0# 3.49fF
C23 a_4864_0# a_4620_0# 3.49fF
C24 a_19260_0# a_19504_0# 3.49fF
C25 a_5352_0# a_5596_0# 3.49fF
C26 a_0_0# w_n176_n86# 9.36fF
C27 a_10476_0# a_10232_0# 3.49fF
C28 a_21212_0# a_21456_0# 3.49fF
C29 a_1936_0# a_1692_0# 3.49fF
C30 a_20236_0# a_19992_0# 3.49fF
C31 a_21944_0# a_22188_0# 3.49fF
C32 a_14868_0# a_15112_0# 3.49fF
C33 a_6572_0# a_6816_0# 3.49fF
C34 a_23408_0# a_23652_0# 3.49fF
C35 a_12184_0# a_12428_0# 3.49fF
C36 a_16820_0# a_16576_0# 3.49fF
C37 a_21456_0# a_21700_0# 3.49fF
C38 a_3644_0# a_3888_0# 3.49fF
C39 a_1204_0# a_960_0# 3.49fF
C40 a_10720_0# a_10964_0# 3.49fF
C41 a_15844_0# a_15600_0# 3.49fF
C42 a_23652_0# a_23896_0# 3.49fF
C43 a_19748_0# a_19504_0# 3.49fF
C44 a_11696_0# a_11940_0# 3.49fF
C45 a_2912_0# a_2668_0# 3.49fF
C46 a_23896_0# a_24140_0# 3.49fF
C47 a_8036_0# a_7792_0# 3.49fF
C48 a_21700_0# a_21944_0# 3.49fF
C49 a_17796_0# a_17552_0# 3.49fF
C50 a_20480_0# a_20236_0# 3.49fF
C51 a_17064_0# a_17308_0# 3.49fF
C52 a_7060_0# a_6816_0# 3.49fF
C53 a_20724_0# a_20968_0# 3.49fF
C54 a_18040_0# a_18284_0# 3.49fF
C55 a_13892_0# a_14136_0# 3.49fF
C56 a_24140_0# a_24384_0# 3.49fF
C57 a_716_0# a_472_0# 3.49fF
C58 a_14380_0# a_14136_0# 3.49fF
C59 a_12672_0# a_12428_0# 3.49fF
C60 a_7304_0# a_7060_0# 3.49fF
C61 a_8768_0# a_8524_0# 3.49fF
C62 a_23164_0# a_23408_0# 3.49fF
C63 a_19016_0# a_18772_0# 3.49fF
C64 a_14868_0# a_14624_0# 3.49fF
C65 a_12184_0# a_11940_0# 3.49fF
C66 a_16332_0# a_16576_0# 3.49fF
C67 a_4132_0# a_3888_0# 3.49fF
C68 a_4132_0# a_4376_0# 3.49fF
C69 a_17308_0# a_17552_0# 3.49fF
C70 a_8768_0# a_9012_0# 3.49fF
C71 a_7548_0# a_7304_0# 3.49fF
C72 a_9500_0# a_9256_0# 3.49fF
C73 a_13160_0# a_12916_0# 3.49fF
C74 a_11696_0# a_11452_0# 3.49fF
C75 a_15356_0# a_15112_0# 3.49fF
C76 a_18528_0# a_18284_0# 3.49fF
C77 a_5108_0# a_4864_0# 3.49fF
C78 a_11208_0# a_10964_0# 3.49fF
C79 a_20480_0# a_20724_0# 3.49fF
C80 a_4376_0# a_4620_0# 3.49fF
C81 a_3156_0# a_2912_0# 3.49fF
C82 a_1448_0# a_1204_0# 3.49fF
C83 a_15600_0# a_15356_0# 3.49fF
C84 a_228_0# a_472_0# 3.49fF
C85 a_7548_0# a_7792_0# 3.49fF
C86 a_1448_0# a_1692_0# 3.49fF
C87 a_13648_0# a_13892_0# 3.49fF
C88 a_9012_0# a_9256_0# 3.49fF
C89 a_5352_0# a_5108_0# 3.49fF
C90 a_17064_0# a_16820_0# 3.49fF
C91 a_13404_0# a_13160_0# 3.49fF
C92 a_3400_0# a_3156_0# 3.49fF
C93 a_11452_0# a_11208_0# 3.49fF
C94 a_9988_0# a_10232_0# 3.49fF
C95 a_6084_0# a_6328_0# 3.49fF
C96 a_9988_0# a_9744_0# 3.49fF
C97 a_13648_0# a_13404_0# 3.49fF
C98 a_960_0# a_716_0# 3.49fF
C99 a_22188_0# a_22432_0# 3.49fF
C100 a_23164_0# a_22920_0# 3.49fF
C101 w_n176_n86# VSUBS 1499.28fF
.ends

.subckt pfet$2 w_n176_n86# a_488_0# a_88_n44# a_0_0# VSUBS
X0 a_488_0# a_88_n44# a_0_0# w_n176_n86# pfet_03v3 ad=4.4p pd=20.88u as=4.4p ps=20.88u w=10u l=2u
C0 w_n176_n86# VSUBS 5.73fF
.ends

.subckt nfet a_592_0# a_15792_0# a_4952_n44# a_13664_0# a_16400_0# a_11336_n44# a_15288_n44#
+ a_11536_0# a_1000_n44# a_5760_0# a_3632_0# a_1504_0# a_5864_n44# a_1912_n44# a_8496_0#
+ a_10320_0# a_17008_0# a_12248_n44# a_6368_0# a_9104_0# a_13160_n44# a_15184_0# a_6776_n44#
+ a_2824_n44# a_7280_0# a_13056_0# a_9208_n44# a_5152_0# a_17920_0# a_3024_0# a_n152_0#
+ a_16504_n44# a_392_n44# a_10120_n44# a_14072_n44# a_7688_n44# a_10928_0# a_3736_n44#
+ a_14984_n44# a_11840_0# a_7888_0# a_17416_n44# a_11032_n44# a_4648_n44# a_14576_0#
+ a_15896_n44# a_17312_0# a_11944_n44# a_5560_n44# a_6672_0# a_12448_0# a_4544_0#
+ a_2416_0# a_1608_n44# a_13360_0# a_8904_n44# a_12856_n44# a_11232_0# a_6472_n44#
+ a_2520_n44# a_1200_0# a_16096_0# a_16200_n44# a_8192_0# a_9816_n44# a_896_0# a_13768_n44#
+ a_6064_0# a_7384_n44# a_3432_n44# a_13968_0# a_16704_0# a_14680_n44# a_8800_0# a_17112_n44#
+ a_3936_0# a_8296_n44# a_10728_n44# a_1808_0# a_14880_0# a_4344_n44# a_12752_0# a_11640_n44#
+ a_15592_n44# a_10624_0# a_88_n44# a_9408_0# a_18024_n44# a_2720_0# a_288_0# a_15488_0#
+ a_18224_0# a_5256_n44# a_1304_n44# a_7584_0# a_8600_n44# a_12552_n44# a_5456_0#
+ a_3328_0# a_14272_0# a_0_0# a_12144_0# a_6168_n44# a_2216_n44# a_9512_n44# a_4240_0#
+ a_10016_0# a_13464_n44# a_7080_n44# a_2112_0# a_7992_n44# a_3128_n44# a_16808_n44#
+ a_696_n44# a_10424_n44# a_14376_n44# a_17616_0# a_4040_n44# a_6976_0# a_9712_0#
+ a_17720_n44# a_4848_0#
X0 a_1808_0# a_1608_n44# a_1504_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X1 a_11232_0# a_11032_n44# a_10928_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X2 a_17616_0# a_17416_n44# a_17312_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X3 a_5760_0# a_5560_n44# a_5456_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X4 a_15184_0# a_14984_n44# a_14880_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X5 a_4848_0# a_4648_n44# a_4544_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X6 a_10320_0# a_10120_n44# a_10016_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X7 a_14272_0# a_14072_n44# a_13968_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X8 a_16704_0# a_16504_n44# a_16400_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X9 a_3936_0# a_3736_n44# a_3632_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X10 a_7888_0# a_7688_n44# a_7584_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X11 a_13360_0# a_13160_n44# a_13056_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X12 a_9408_0# a_9208_n44# a_9104_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X13 a_12448_0# a_12248_n44# a_12144_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X14 a_3024_0# a_2824_n44# a_2720_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X15 a_6976_0# a_6776_n44# a_6672_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X16 a_11536_0# a_11336_n44# a_11232_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X17 a_15488_0# a_15288_n44# a_15184_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X18 a_2112_0# a_1912_n44# a_1808_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X19 a_6064_0# a_5864_n44# a_5760_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X20 a_1200_0# a_1000_n44# a_896_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X21 a_10624_0# a_10424_n44# a_10320_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X22 a_14576_0# a_14376_n44# a_14272_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X23 a_17920_0# a_17720_n44# a_17616_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X24 a_17008_0# a_16808_n44# a_16704_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X25 a_5152_0# a_4952_n44# a_4848_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X26 a_4240_0# a_4040_n44# a_3936_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X27 a_13664_0# a_13464_n44# a_13360_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X28 a_3328_0# a_3128_n44# a_3024_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X29 a_592_0# a_392_n44# a_288_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X30 a_8192_0# a_7992_n44# a_7888_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X31 a_7280_0# a_7080_n44# a_6976_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X32 a_9712_0# a_9512_n44# a_9408_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X33 a_12752_0# a_12552_n44# a_12448_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X34 a_288_0# a_88_n44# a_0_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=26.4p ps=120.88u w=60u l=1000n
X35 a_2416_0# a_2216_n44# a_2112_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X36 a_6368_0# a_6168_n44# a_6064_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X37 a_18224_0# a_18024_n44# a_17920_0# a_n152_0# nfet_03v3 ad=26.4p pd=120.88u as=15.6p ps=60.52u w=60u l=1000n
X38 a_8800_0# a_8600_n44# a_8496_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X39 a_11840_0# a_11640_n44# a_11536_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X40 a_15792_0# a_15592_n44# a_15488_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X41 a_1504_0# a_1304_n44# a_1200_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X42 a_5456_0# a_5256_n44# a_5152_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X43 a_10928_0# a_10728_n44# a_10624_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X44 a_17312_0# a_17112_n44# a_17008_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X45 a_14880_0# a_14680_n44# a_14576_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X46 a_4544_0# a_4344_n44# a_4240_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X47 a_8496_0# a_8296_n44# a_8192_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X48 a_13968_0# a_13768_n44# a_13664_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X49 a_896_0# a_696_n44# a_592_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X50 a_16400_0# a_16200_n44# a_16096_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X51 a_3632_0# a_3432_n44# a_3328_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X52 a_7584_0# a_7384_n44# a_7280_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X53 a_10016_0# a_9816_n44# a_9712_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X54 a_13056_0# a_12856_n44# a_12752_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X55 a_2720_0# a_2520_n44# a_2416_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X56 a_6672_0# a_6472_n44# a_6368_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X57 a_12144_0# a_11944_n44# a_11840_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X58 a_9104_0# a_8904_n44# a_8800_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
X59 a_16096_0# a_15896_n44# a_15792_0# a_n152_0# nfet_03v3 ad=15.6p pd=60.52u as=15.6p ps=60.52u w=60u l=1000n
C0 a_0_0# a_n152_0# 5.64fF
.ends

.subckt nfet$4 a_n152_0# a_88_n44# a_288_0# a_0_0#
X0 a_288_0# a_88_n44# a_0_0# a_n152_0# nfet_03v3 ad=8.8p pd=40.88u as=8.8p ps=40.88u w=20u l=1000n
.ends

.subckt OTA_2stage vout vss vin1 vin2 vp vdd
Xpfet_0 a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096# vdd vdd
+ vdd vdd a_155465_201096# a_155465_201096# vdd a_155465_201096# a_155465_201096#
+ a_213587_216449# a_155465_201096# a_213587_216449# vdd a_155465_201096# a_213587_216449#
+ a_155465_201096# a_155465_201096# a_155465_201096# vdd a_155465_201096# a_213587_216449#
+ vdd a_155465_201096# vdd a_213587_216449# a_155465_201096# a_213587_216449# vdd
+ a_213587_216449# vdd a_213587_216449# vdd a_155465_201096# a_155465_201096# a_155465_201096#
+ a_155465_201096# a_155465_201096# a_155465_201096# vdd a_155465_201096# a_155465_201096#
+ vdd a_155465_201096# a_155465_201096# a_213587_216449# a_213587_216449# a_213587_216449#
+ a_155465_201096# a_213587_216449# a_155465_201096# a_213587_216449# a_213587_216449#
+ vdd a_155465_201096# a_155465_201096# vdd a_155465_201096# vdd vdd vdd a_155465_201096#
+ a_155465_201096# a_155465_201096# vdd a_155465_201096# a_155465_201096# vdd a_155465_201096#
+ vdd a_213587_216449# a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096#
+ a_213587_216449# a_213587_216449# a_155465_201096# vdd a_213587_216449# a_213587_216449#
+ a_213587_216449# a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096#
+ a_213587_216449# a_155465_201096# a_213587_216449# a_155465_201096# vdd a_213587_216449#
+ vdd a_155465_201096# a_213587_216449# vdd a_155465_201096# a_213587_216449# vss
+ vdd pfet
Xnfet$2_37 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_26 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_15 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_2 vss vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vout vout
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss vout vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vout vout
+ a_49909_45330# vss vout vss vss vss vout a_49909_45330# vss a_49909_45330# vss vss
+ vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss
+ vout vout a_49909_45330# vout a_49909_45330# vout vss vss a_49909_45330# a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# vss a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vss a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss a_49909_45330# vss vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330# a_49909_45330#
+ vout vout vss a_49909_45330# a_49909_45330# vss a_49909_45330# vss a_49909_45330#
+ vout a_49909_45330# vout a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout vss vout vss a_49909_45330# vout a_49909_45330# vout vss
+ a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vss vout a_49909_45330#
+ vout a_49909_45330# a_49909_45330# vout vout vss vout a_49909_45330# a_49909_45330#
+ a_49909_45330# a_49909_45330# vss vss vout vout vout a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# vout vout vss a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# vout a_49909_45330# vout a_49909_45330# vout a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# a_49909_45330# vss vss a_49909_45330#
+ a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330# vss nfet$2
Xpfet_1 a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096# vdd vdd
+ vdd vdd a_155465_201096# a_155465_201096# vdd a_155465_201096# a_155465_201096#
+ a_155465_201096# a_155465_201096# a_155465_201096# vdd a_155465_201096# a_155465_201096#
+ a_155465_201096# a_155465_201096# a_155465_201096# vdd a_155465_201096# a_155465_201096#
+ vdd a_155465_201096# vdd a_155465_201096# a_155465_201096# a_155465_201096# vdd
+ a_155465_201096# vdd a_155465_201096# vdd a_155465_201096# a_155465_201096# a_155465_201096#
+ a_155465_201096# a_155465_201096# a_155465_201096# vdd a_155465_201096# a_155465_201096#
+ vdd a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096#
+ a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096#
+ vdd a_155465_201096# a_155465_201096# vdd a_155465_201096# vdd vdd vdd a_155465_201096#
+ a_155465_201096# a_155465_201096# vdd a_155465_201096# a_155465_201096# vdd a_155465_201096#
+ vdd a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096#
+ a_155465_201096# a_155465_201096# a_155465_201096# vdd a_155465_201096# a_155465_201096#
+ a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096#
+ a_155465_201096# a_155465_201096# a_155465_201096# a_155465_201096# vdd a_155465_201096#
+ vdd a_155465_201096# a_155465_201096# vdd a_155465_201096# a_155465_201096# vss
+ vdd pfet
Xnfet$2_38 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_27 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_16 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_4 vss vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vout vout
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss vout vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vout vout
+ a_49909_45330# vss vout vss vss vss vout a_49909_45330# vss a_49909_45330# vss vss
+ vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss
+ vout vout a_49909_45330# vout a_49909_45330# vout vss vss a_49909_45330# a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# vss a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vss a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss a_49909_45330# vss vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330# a_49909_45330#
+ vout vout vss a_49909_45330# a_49909_45330# vss a_49909_45330# vss a_49909_45330#
+ vout a_49909_45330# vout a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout vss vout vss a_49909_45330# vout a_49909_45330# vout vss
+ a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vss vout a_49909_45330#
+ vout a_49909_45330# a_49909_45330# vout vout vss vout a_49909_45330# a_49909_45330#
+ a_49909_45330# a_49909_45330# vss vss vout vout vout a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# vout vout vss a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# vout a_49909_45330# vout a_49909_45330# vout a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# a_49909_45330# vss vss a_49909_45330#
+ a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330# vss nfet$2
Xnfet$2_3 vss vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vout vout
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss vout vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vout vout
+ a_49909_45330# vss vout vss vss vss vout a_49909_45330# vss a_49909_45330# vss vss
+ vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss
+ vout vout a_49909_45330# vout a_49909_45330# vout vss vss a_49909_45330# a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# vss a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vss a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss a_49909_45330# vss vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330# a_49909_45330#
+ vout vout vss a_49909_45330# a_49909_45330# vss a_49909_45330# vss a_49909_45330#
+ vout a_49909_45330# vout a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout vss vout vss a_49909_45330# vout a_49909_45330# vout vss
+ a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vss vout a_49909_45330#
+ vout a_49909_45330# a_49909_45330# vout vout vss vout a_49909_45330# a_49909_45330#
+ a_49909_45330# a_49909_45330# vss vss vout vout vout a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# vout vout vss a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# vout a_49909_45330# vout a_49909_45330# vout a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# a_49909_45330# vss vss a_49909_45330#
+ a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330# vss nfet$2
Xnfet$2_39 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_28 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_17 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_5 vss vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vout vout
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss vout vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vout vout
+ a_49909_45330# vss vout vss vss vss vout a_49909_45330# vss a_49909_45330# vss vss
+ vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss
+ vout vout a_49909_45330# vout a_49909_45330# vout vss vss a_49909_45330# a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# vss a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vss a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss a_49909_45330# vss vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330# a_49909_45330#
+ vout vout vss a_49909_45330# a_49909_45330# vss a_49909_45330# vss a_49909_45330#
+ vout a_49909_45330# vout a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout vss vout vss a_49909_45330# vout a_49909_45330# vout vss
+ a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vss vout a_49909_45330#
+ vout a_49909_45330# a_49909_45330# vout vout vss vout a_49909_45330# a_49909_45330#
+ a_49909_45330# a_49909_45330# vss vss vout vout vout a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# vout vout vss a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# vout a_49909_45330# vout a_49909_45330# vout a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# a_49909_45330# vss vss a_49909_45330#
+ a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330# vss nfet$2
Xnfet$2_29 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_19 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_18 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_6 vss vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vout vout
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss vout vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vout vout
+ a_49909_45330# vss vout vss vss vss vout a_49909_45330# vss a_49909_45330# vss vss
+ vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss
+ vout vout a_49909_45330# vout a_49909_45330# vout vss vss a_49909_45330# a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# vss a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vss a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss a_49909_45330# vss vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330# a_49909_45330#
+ vout vout vss a_49909_45330# a_49909_45330# vss a_49909_45330# vss a_49909_45330#
+ vout a_49909_45330# vout a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout vss vout vss a_49909_45330# vout a_49909_45330# vout vss
+ a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vss vout a_49909_45330#
+ vout a_49909_45330# a_49909_45330# vout vout vss vout a_49909_45330# a_49909_45330#
+ a_49909_45330# a_49909_45330# vss vss vout vout vout a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# vout vout vss a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# vout a_49909_45330# vout a_49909_45330# vout a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# a_49909_45330# vss vss a_49909_45330#
+ a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330# vss nfet$2
Xnfet$2_7 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_8 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xpfet$4_0 vout vdd a_213587_216449# a_213587_216449# vdd vout vdd a_213587_216449#
+ vdd vdd a_213587_216449# a_213587_216449# vout a_213587_216449# vout vdd vdd vout
+ vdd vdd a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# vdd vout vout vout vdd vdd a_213587_216449# a_213587_216449# vdd
+ vout a_213587_216449# a_213587_216449# a_213587_216449# vdd vdd a_213587_216449#
+ vdd a_213587_216449# a_213587_216449# vdd vout a_213587_216449# vdd a_213587_216449#
+ a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ vdd a_213587_216449# a_213587_216449# vdd vdd vout a_213587_216449# a_213587_216449#
+ vout vdd vout a_213587_216449# a_213587_216449# a_213587_216449# vdd vdd a_213587_216449#
+ vdd vout a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ vdd vdd vdd vout a_213587_216449# a_213587_216449# vdd a_213587_216449# vout a_213587_216449#
+ vout a_213587_216449# vdd vout vdd a_213587_216449# vout a_213587_216449# vdd vout
+ vout vdd vout a_213587_216449# a_213587_216449# vout vdd a_213587_216449# vout a_213587_216449#
+ a_213587_216449# vout vdd a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# vdd vout a_213587_216449# vout vout vout vdd a_213587_216449#
+ a_213587_216449# vout vout vdd a_213587_216449# a_213587_216449# a_213587_216449#
+ vout vout a_213587_216449# a_213587_216449# vdd a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# a_213587_216449# vdd a_213587_216449# a_213587_216449#
+ vout a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449# vout
+ a_213587_216449# a_213587_216449# a_213587_216449# vdd vout vdd vout a_213587_216449#
+ a_213587_216449# vdd vdd a_213587_216449# vout vdd a_213587_216449# vout a_213587_216449#
+ vdd a_213587_216449# vout vout a_213587_216449# a_213587_216449# vdd a_213587_216449#
+ a_213587_216449# vout vout vdd a_213587_216449# a_213587_216449# vout vout a_213587_216449#
+ a_213587_216449# vout vdd vdd vout vdd a_213587_216449# a_213587_216449# vss vdd
+ pfet$4
Xnfet$2_9 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xpfet$4_1 vout vdd a_213587_216449# a_213587_216449# vdd vout vdd a_213587_216449#
+ vdd vdd a_213587_216449# a_213587_216449# vout a_213587_216449# vout vdd vdd vout
+ vdd vdd a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# vdd vout vout vout vdd vdd a_213587_216449# a_213587_216449# vdd
+ vout a_213587_216449# a_213587_216449# a_213587_216449# vdd vdd a_213587_216449#
+ vdd a_213587_216449# a_213587_216449# vdd vout a_213587_216449# vdd a_213587_216449#
+ a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ vdd a_213587_216449# a_213587_216449# vdd vdd vout a_213587_216449# a_213587_216449#
+ vout vdd vout a_213587_216449# a_213587_216449# a_213587_216449# vdd vdd a_213587_216449#
+ vdd vout a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ vdd vdd vdd vout a_213587_216449# a_213587_216449# vdd a_213587_216449# vout a_213587_216449#
+ vout a_213587_216449# vdd vout vdd a_213587_216449# vout a_213587_216449# vdd vout
+ vout vdd vout a_213587_216449# a_213587_216449# vout vdd a_213587_216449# vout a_213587_216449#
+ a_213587_216449# vout vdd a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# vdd vout a_213587_216449# vout vout vout vdd a_213587_216449#
+ a_213587_216449# vout vout vdd a_213587_216449# a_213587_216449# a_213587_216449#
+ vout vout a_213587_216449# a_213587_216449# vdd a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# a_213587_216449# vdd a_213587_216449# a_213587_216449#
+ vout a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449# vout
+ a_213587_216449# a_213587_216449# a_213587_216449# vdd vout vdd vout a_213587_216449#
+ a_213587_216449# vdd vdd a_213587_216449# vout vdd a_213587_216449# vout a_213587_216449#
+ vdd a_213587_216449# vout vout a_213587_216449# a_213587_216449# vdd a_213587_216449#
+ a_213587_216449# vout vout vdd a_213587_216449# a_213587_216449# vout vout a_213587_216449#
+ a_213587_216449# vout vdd vdd vout vdd a_213587_216449# a_213587_216449# vss vdd
+ pfet$4
Xpfet$4_2 vout vdd a_213587_216449# a_213587_216449# vdd vout vdd a_213587_216449#
+ vdd vdd a_213587_216449# a_213587_216449# vout a_213587_216449# vout vdd vdd vout
+ vdd vdd a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# vdd vout vout vout vdd vdd a_213587_216449# a_213587_216449# vdd
+ vout a_213587_216449# a_213587_216449# a_213587_216449# vdd vdd a_213587_216449#
+ vdd a_213587_216449# a_213587_216449# vdd vout a_213587_216449# vdd a_213587_216449#
+ a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ vdd a_213587_216449# a_213587_216449# vdd vdd vout a_213587_216449# a_213587_216449#
+ vout vdd vout a_213587_216449# a_213587_216449# a_213587_216449# vdd vdd a_213587_216449#
+ vdd vout a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ vdd vdd vdd vout a_213587_216449# a_213587_216449# vdd a_213587_216449# vout a_213587_216449#
+ vout a_213587_216449# vdd vout vdd a_213587_216449# vout a_213587_216449# vdd vout
+ vout vdd vout a_213587_216449# a_213587_216449# vout vdd a_213587_216449# vout a_213587_216449#
+ a_213587_216449# vout vdd a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# vdd vout a_213587_216449# vout vout vout vdd a_213587_216449#
+ a_213587_216449# vout vout vdd a_213587_216449# a_213587_216449# a_213587_216449#
+ vout vout a_213587_216449# a_213587_216449# vdd a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# a_213587_216449# vdd a_213587_216449# a_213587_216449#
+ vout a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449# vout
+ a_213587_216449# a_213587_216449# a_213587_216449# vdd vout vdd vout a_213587_216449#
+ a_213587_216449# vdd vdd a_213587_216449# vout vdd a_213587_216449# vout a_213587_216449#
+ vdd a_213587_216449# vout vout a_213587_216449# a_213587_216449# vdd a_213587_216449#
+ a_213587_216449# vout vout vdd a_213587_216449# a_213587_216449# vout vout a_213587_216449#
+ a_213587_216449# vout vdd vdd vout vdd a_213587_216449# a_213587_216449# vss vdd
+ pfet$4
Xpfet$2_0 vdd a_49909_45330# vp vdd vss pfet$2
Xpfet$4_3 vout vdd a_213587_216449# a_213587_216449# vdd vout vdd a_213587_216449#
+ vdd vdd a_213587_216449# a_213587_216449# vout a_213587_216449# vout vdd vdd vout
+ vdd vdd a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# vdd vout vout vout vdd vdd a_213587_216449# a_213587_216449# vdd
+ vout a_213587_216449# a_213587_216449# a_213587_216449# vdd vdd a_213587_216449#
+ vdd a_213587_216449# a_213587_216449# vdd vout a_213587_216449# vdd a_213587_216449#
+ a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ vdd a_213587_216449# a_213587_216449# vdd vdd vout a_213587_216449# a_213587_216449#
+ vout vdd vout a_213587_216449# a_213587_216449# a_213587_216449# vdd vdd a_213587_216449#
+ vdd vout a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ vdd vdd vdd vout a_213587_216449# a_213587_216449# vdd a_213587_216449# vout a_213587_216449#
+ vout a_213587_216449# vdd vout vdd a_213587_216449# vout a_213587_216449# vdd vout
+ vout vdd vout a_213587_216449# a_213587_216449# vout vdd a_213587_216449# vout a_213587_216449#
+ a_213587_216449# vout vdd a_213587_216449# a_213587_216449# a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# vdd vout a_213587_216449# vout vout vout vdd a_213587_216449#
+ a_213587_216449# vout vout vdd a_213587_216449# a_213587_216449# a_213587_216449#
+ vout vout a_213587_216449# a_213587_216449# vdd a_213587_216449# a_213587_216449#
+ a_213587_216449# a_213587_216449# a_213587_216449# vdd a_213587_216449# a_213587_216449#
+ vout a_213587_216449# vout a_213587_216449# a_213587_216449# a_213587_216449# vout
+ a_213587_216449# a_213587_216449# a_213587_216449# vdd vout vdd vout a_213587_216449#
+ a_213587_216449# vdd vdd a_213587_216449# vout vdd a_213587_216449# vout a_213587_216449#
+ vdd a_213587_216449# vout vout a_213587_216449# a_213587_216449# vdd a_213587_216449#
+ a_213587_216449# vout vout vdd a_213587_216449# a_213587_216449# vout vout a_213587_216449#
+ a_213587_216449# vout vdd vdd vout vdd a_213587_216449# a_213587_216449# vss vdd
+ pfet$4
Xnfet_0 vss vss a_49909_45330# vss vss a_49909_45330# a_49909_45330# vss a_49909_45330#
+ vss vss vss a_49909_45330# a_49909_45330# vss vss vss a_49909_45330# vss vss a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vss vss a_49909_45330# vss vss vss vss a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss a_49909_45330# a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# vss a_49909_45330# vss a_49909_45330#
+ a_49909_45330# vss vss vss vss a_49909_45330# vss a_49909_45330# a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vss vss a_49909_45330# vss a_49909_45330# vss
+ a_49909_45330# vss a_49909_45330# a_49909_45330# vss vss a_49909_45330# vss a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vss vss a_49909_45330# vss a_49909_45330# a_49909_45330#
+ vss a_49909_45330# vss a_49909_45330# vss vss vss vss a_49909_45330# a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vss vss vss vss vss a_49909_45330# a_49909_45330#
+ a_49909_45330# vss vss a_49909_45330# a_49909_45330# vss a_49909_45330# a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss a_49909_45330# vss
+ vss a_49909_45330# vss nfet
Xnfet$2_40 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_41 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_30 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_42 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_32 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_31 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_21 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_20 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_10 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$4_0 vss a_49909_45330# a_49909_45330# vss nfet$4
Xnfet$2_33 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_22 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_11 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_34 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_23 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_12 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_35 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_24 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_13 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_0 vss vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vout vout
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss vout vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vout vout
+ a_49909_45330# vss vout vss vss vss vout a_49909_45330# vss a_49909_45330# vss vss
+ vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss
+ vout vout a_49909_45330# vout a_49909_45330# vout vss vss a_49909_45330# a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# vss a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vss a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss a_49909_45330# vss vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330# a_49909_45330#
+ vout vout vss a_49909_45330# a_49909_45330# vss a_49909_45330# vss a_49909_45330#
+ vout a_49909_45330# vout a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout vss vout vss a_49909_45330# vout a_49909_45330# vout vss
+ a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vss vout a_49909_45330#
+ vout a_49909_45330# a_49909_45330# vout vout vss vout a_49909_45330# a_49909_45330#
+ a_49909_45330# a_49909_45330# vss vss vout vout vout a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# vout vout vss a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# vout a_49909_45330# vout a_49909_45330# vout a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# a_49909_45330# vss vss a_49909_45330#
+ a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330# vss nfet$2
Xnfet$2_36 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_25 vss vss vss vin1 vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096#
+ vss vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss a_155465_201096# vss vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vin1 vss a_155465_201096# vss vss
+ vss a_155465_201096# vin1 vss vin1 vss vss vss vin1 vin1 vin1 vin1 vin1 vss a_155465_201096#
+ a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096# vss vss vin1 vin1 vss
+ vss vin1 vin1 vss vin1 vin1 vin1 vin1 vss vin1 vin1 a_155465_201096# a_155465_201096#
+ a_155465_201096# vss vin1 vin1 vin1 vin1 vss vin1 vss vss a_155465_201096# vin1
+ vin1 vin1 vin1 vss a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096#
+ vss vin1 vin1 vss vin1 vss vin1 a_155465_201096# vin1 a_155465_201096# vin1 vin1
+ vin1 vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vss vin1 a_155465_201096#
+ vin1 a_155465_201096# vss vin1 vin1 vin1 vin1 vss vss a_155465_201096# vin1 a_155465_201096#
+ vin1 vin1 a_155465_201096# a_155465_201096# vss a_155465_201096# vin1 vin1 vin1
+ vin1 vss vss a_155465_201096# a_155465_201096# a_155465_201096# vin1 vin1 vin1 a_155465_201096#
+ a_155465_201096# vin1 vin1 a_155465_201096# a_155465_201096# a_155465_201096# vss
+ vin1 vss vin1 vin1 vin1 a_155465_201096# vss vin1 vin1 vss vin1 vin1 a_155465_201096#
+ vin1 a_155465_201096# a_155465_201096# vss vin1 vss vss vin1 vin1 vin1 vin1 vss
+ a_155465_201096# vin1 vin1 vin1 a_155465_201096# vin1 a_155465_201096# vin1 a_155465_201096#
+ vin1 vss vin1 vin1 a_155465_201096# vin1 vin1 vss vss vin1 vin1 vin1 a_155465_201096#
+ vss vin1 vin1 vss nfet$2
Xnfet$2_14 vss vss vss vin2 vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449#
+ vss vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss a_213587_216449# vss vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vin2 vss a_213587_216449# vss vss
+ vss a_213587_216449# vin2 vss vin2 vss vss vss vin2 vin2 vin2 vin2 vin2 vss a_213587_216449#
+ a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449# vss vss vin2 vin2 vss
+ vss vin2 vin2 vss vin2 vin2 vin2 vin2 vss vin2 vin2 a_213587_216449# a_213587_216449#
+ a_213587_216449# vss vin2 vin2 vin2 vin2 vss vin2 vss vss a_213587_216449# vin2
+ vin2 vin2 vin2 vss a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449#
+ vss vin2 vin2 vss vin2 vss vin2 a_213587_216449# vin2 a_213587_216449# vin2 vin2
+ vin2 vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vss vin2 a_213587_216449#
+ vin2 a_213587_216449# vss vin2 vin2 vin2 vin2 vss vss a_213587_216449# vin2 a_213587_216449#
+ vin2 vin2 a_213587_216449# a_213587_216449# vss a_213587_216449# vin2 vin2 vin2
+ vin2 vss vss a_213587_216449# a_213587_216449# a_213587_216449# vin2 vin2 vin2 a_213587_216449#
+ a_213587_216449# vin2 vin2 a_213587_216449# a_213587_216449# a_213587_216449# vss
+ vin2 vss vin2 vin2 vin2 a_213587_216449# vss vin2 vin2 vss vin2 vin2 a_213587_216449#
+ vin2 a_213587_216449# a_213587_216449# vss vin2 vss vss vin2 vin2 vin2 vin2 vss
+ a_213587_216449# vin2 vin2 vin2 a_213587_216449# vin2 a_213587_216449# vin2 a_213587_216449#
+ vin2 vss vin2 vin2 a_213587_216449# vin2 vin2 vss vss vin2 vin2 vin2 a_213587_216449#
+ vss vin2 vin2 vss nfet$2
Xnfet$2_1 vss vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vout vout
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss vout vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vout vout
+ a_49909_45330# vss vout vss vss vss vout a_49909_45330# vss a_49909_45330# vss vss
+ vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss
+ vout vout a_49909_45330# vout a_49909_45330# vout vss vss a_49909_45330# a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# vss a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vss a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss a_49909_45330# vss vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330# a_49909_45330#
+ vout vout vss a_49909_45330# a_49909_45330# vss a_49909_45330# vss a_49909_45330#
+ vout a_49909_45330# vout a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout vss vout vss a_49909_45330# vout a_49909_45330# vout vss
+ a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vss vout a_49909_45330#
+ vout a_49909_45330# a_49909_45330# vout vout vss vout a_49909_45330# a_49909_45330#
+ a_49909_45330# a_49909_45330# vss vss vout vout vout a_49909_45330# a_49909_45330#
+ a_49909_45330# vout vout a_49909_45330# a_49909_45330# vout vout vout vss a_49909_45330#
+ vss a_49909_45330# a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# vout vout vss a_49909_45330#
+ vss vss a_49909_45330# a_49909_45330# a_49909_45330# a_49909_45330# vss vout a_49909_45330#
+ a_49909_45330# a_49909_45330# vout a_49909_45330# vout a_49909_45330# vout a_49909_45330#
+ vss a_49909_45330# a_49909_45330# vout a_49909_45330# a_49909_45330# vss vss a_49909_45330#
+ a_49909_45330# a_49909_45330# vout vss a_49909_45330# a_49909_45330# vss nfet$2
X0 a_213587_216449# a_141890_183202# vdd ppolyf_u r_width=39.75u r_length=25u
X1 vout a_141890_183202# cap_mim_2f0_m4m5_noshield c_width=100u c_length=125u
X2 vout a_141890_183202# cap_mim_2f0_m4m5_noshield c_width=100u c_length=125u
X3 vout a_141890_183202# cap_mim_2f0_m4m5_noshield c_width=100u c_length=125u
X4 vout vss cap_mim_2f0_m4m5_noshield c_width=125u c_length=100u
C0 a_155465_201096# m3_270065_28942# 62.15fF
C1 m1_336658_16084# vss 471.18fF
C2 a_143326_204039# m3_17923_28702# 46.25fF
C3 a_155465_201096# m3_17923_28702# 1698.21fF
C4 a_18229_167177# m3_17923_28702# 171.33fF
C5 vout m3_270065_28942# 2520.42fF
C6 a_155465_201096# m2_316327_22594# 227.43fF
C7 vout m1_270384_178745# 590.02fF
C8 a_49909_45330# m2_89552_16161# 42.08fF
C9 vin1 a_155465_201096# 866.53fF
C10 vout m3_17923_28702# 202.81fF
C11 m4_270065_28942# m5_271138_28942# 613.61fF
C12 a_155465_201096# m2_275886_12791# 232.66fF
C13 a_213587_216449# m3_270065_28942# 81.73fF
C14 vdd a_141890_183202# 70.14fF
C15 vdd a_49909_45330# 8.26fF
C16 vout m2_316327_22594# 161.10fF
C17 vin1 vout 171.32fF
C18 a_155465_201096# m2_247088_16161# 178.47fF
C19 a_213587_216449# m3_17923_28702# 5723.39fF
C20 vout m2_275886_12791# 395.49fF
C21 m4_17923_28702# m5_21063_28702# 68.31fF
C22 m3_270065_28942# m5_271138_28942# 3.67fF
C23 a_213587_216449# m2_316327_22594# 276.10fF
C24 vout m2_247088_16161# 229.39fF
C25 vin1 a_213587_216449# 404.71fF
C26 a_18229_167177# m1_22935_171882# 30.11fF
C27 a_155465_201096# m2_207566_53538# 291.80fF
C28 a_213587_216449# m2_275886_12791# 287.96fF
C29 vout m2_104013_15854# 1441.91fF
C30 m3_17923_28702# m5_21063_28702# 18.90fF
C31 m3_270065_28942# m4_270065_28942# 23.01fF
C32 vin2 vout 171.32fF
C33 a_19014_30903# vss 321.94fF
C34 a_213587_216449# m2_247088_16161# 264.27fF
C35 a_119209_165804# m2_68719_172226# 120.67fF
C36 m1_270384_178745# m4_270065_28942# 265.87fF
C37 vout m2_207566_53538# 70.81fF
C38 m1_22212_14629# m3_17923_28702# 984.86fF
C39 m3_17923_28702# m4_17923_28702# 505.63fF
C40 vin2 a_213587_216449# 1115.10fF
C41 a_213587_216449# m2_207566_53538# 416.41fF
C42 vdd a_143326_204039# 1028.24fF
C43 m1_336854_101883# vss 187.31fF
C44 vin1 m1_22212_14629# 203.76fF
C45 vdd a_155465_201096# 20.24fF
C46 a_155465_201096# m2_88082_114628# 523.99fF
C47 a_213587_216449# m2_156402_54151# 435.24fF
C48 vout m2_89552_16161# 61.99fF
C49 m2_104013_15854# m5_21063_28702# 7.63fF
C50 m2_316327_22594# m3_270065_28942# 4.51fF
C51 vin1 m3_270065_28942# 117.68fF
C52 a_213587_216449# m2_117187_51087# 288.50fF
C53 a_18229_167177# m2_68719_172226# 3.14fF
C54 a_269011_166588# m1_336854_101883# 20.20fF
C55 vdd vout 8.32fF
C56 m2_275886_12791# m3_270065_28942# 7.17fF
C57 vin1 m3_17923_28702# 622.23fF
C58 a_213587_216449# m2_89552_16161# 172.67fF
C59 m1_270384_178745# m2_275886_12791# 102.16fF
C60 m2_104013_15854# m4_17923_28702# 10.95fF
C61 vin1 m2_316327_22594# 252.66fF
C62 vdd a_213587_216449# 176.13fF
C63 vin1 m2_275886_12791# 294.30fF
C64 vin2 m3_270065_28942# 199.41fF
C65 m2_104013_15854# m3_17923_28702# 24.30fF
C66 vin1 m2_247088_16161# 224.45fF
C67 vin2 m3_17923_28702# 542.82fF
C68 a_335678_28942# m3_270065_28942# 98.24fF
C69 vin2 m2_316327_22594# 303.27fF
C70 m2_156402_54151# m3_17923_28702# 2418.42fF
C71 vin1 m2_207566_53538# 367.94fF
C72 vin2 m2_275886_12791# 294.30fF
C73 a_269011_166588# vss 168.16fF
C74 a_335678_28942# m2_316327_22594# 24.43fF
C75 a_335089_106785# m3_270065_28942# 121.33fF
C76 m2_117187_51087# m3_17923_28702# 1631.68fF
C77 vin2 m2_247088_16161# 224.45fF
C78 a_153914_166588# vss 119.06fF
C79 m2_89552_16161# m3_17923_28702# 1320.19fF
C80 a_335089_106785# m2_316327_22594# 48.33fF
C81 vdd m3_17923_28702# 1062.35fF
C82 vin2 m2_207566_53538# 367.94fF
C83 a_49909_45330# vss 519.17fF
C84 m1_336658_16084# m3_270065_28942# 148.80fF
C85 m2_68719_172226# m3_17923_28702# 1507.90fF
C86 vin1 m2_88082_114628# 683.82fF
C87 vin2 m2_156402_54151# 436.21fF
C88 vin2 m2_117187_51087# 294.92fF
C89 a_141890_183202# a_269011_166588# 3.09fF
C90 vdd m2_247088_16161# 39.75fF
C91 m1_336658_16084# m2_316327_22594# 364.61fF
C92 vin2 m2_89552_16161# 173.37fF
C93 a_119209_165804# vss 61.29fF
C94 vdd m2_207566_53538# 75.66fF
C95 m1_22935_171882# m2_68719_172226# 1161.30fF
C96 vin2 m1_336658_16084# 88.91fF
C97 a_19014_30903# m1_22212_14629# 2196.54fF
C98 a_155465_201096# vss 500.97fF
C99 a_18229_167177# vss 92.83fF
C100 a_335678_28942# m1_336658_16084# 830.04fF
C101 m1_336854_101883# m4_270065_28942# 3.47fF
C102 a_49909_45330# a_119209_165804# 86.96fF
C103 vout vss 650.28fF
C104 a_19014_30903# m3_17923_28702# 178.67fF
C105 vp m3_17923_28702# 148.69fF
C106 m1_336854_101883# m3_270065_28942# 128.70fF
C107 a_155465_201096# a_153914_166588# 477.37fF
C108 a_213587_216449# vss 1037.73fF
C109 vout a_269011_166588# 746.93fF
C110 m1_336854_101883# m2_316327_22594# 330.02fF
C111 a_155465_201096# a_141890_183202# 110.32fF
C112 a_49909_45330# a_155465_201096# 113.57fF
C113 a_49909_45330# a_18229_167177# 17.41fF
C114 a_213587_216449# a_153914_166588# 333.39fF
C115 vout a_141890_183202# 70.86fF
C116 m4_270065_28942# vss 68.57fF
C117 a_49909_45330# vout 80.13fF
C118 vp m1_22935_171882# 7.86fF
C119 m4_17923_28702# vss 4.82fF
C120 vin2 m1_336854_101883# 25.74fF
C121 a_213587_216449# a_141890_183202# 114.91fF
C122 a_49909_45330# a_213587_216449# 141.18fF
C123 m3_270065_28942# vss 1093.82fF
C124 a_269011_166588# m4_270065_28942# 80.45fF
C125 m1_270384_178745# vss 63.55fF
C126 m3_17923_28702# vss 5933.66fF
C127 m2_316327_22594# vss 575.21fF
C128 vin1 vss 1161.91fF
C129 vp vdd 3.96fF
C130 a_269011_166588# m1_270384_178745# 25.78fF
C131 m2_275886_12791# vss 910.51fF
C132 a_335089_106785# m1_336854_101883# 678.21fF
C133 a_141890_183202# m4_270065_28942# 19.37fF
C134 m2_247088_16161# vss 660.41fF
C135 a_153914_166588# m3_17923_28702# 84.60fF
C136 a_155465_201096# vout 137.28fF
C137 a_269011_166588# m2_275886_12791# 44.38fF
C138 m2_104013_15854# vss 1252.19fF
C139 a_49909_45330# m3_270065_28942# 49.05fF
C140 vin2 vss 1074.92fF
C141 a_141890_183202# m1_270384_178745# 144.59fF
C142 m2_207566_53538# vss 733.95fF
C143 a_141890_183202# m3_17923_28702# 541.56fF
C144 a_49909_45330# m3_17923_28702# 2674.39fF
C145 a_155465_201096# a_213587_216449# 326.06fF
C146 m2_156402_54151# vss 351.69fF
C147 a_49909_45330# m2_316327_22594# 89.44fF
C148 a_49909_45330# vin1 144.29fF
C149 a_213587_216449# vout 270.58fF
C150 m2_117187_51087# vss 311.50fF
C151 a_49909_45330# m2_275886_12791# 126.72fF
C152 a_335089_106785# vss 60.02fF
C153 a_153914_166588# m2_207566_53538# 24.41fF
C154 a_119209_165804# m3_17923_28702# 63.29fF
C155 m2_89552_16161# vss 246.84fF
C156 a_49909_45330# m2_247088_16161# 96.12fF
C157 m2_88082_114628# vss 710.32fF
C158 a_49909_45330# m2_104013_15854# 697.23fF
C159 a_49909_45330# vin2 144.29fF
C160 a_49909_45330# m1_22935_171882# 770.82fF
C161 vout m4_270065_28942# 174.27fF
C162 vss 0 4445.83fF
C189 a_141890_183202# 0 112.63fF
C193 vout 0 1204.34fF
C194 a_213587_216449# 0 1667.23fF
C195 vin2 0 5786.09fF
C196 a_155465_201096# 0 603.41fF
C197 vin1 0 5775.28fF
C198 a_49909_45330# 0 1371.98fF
C199 vdd 0 8560.55fF
C200 vp 0 1233.65fF
.ends

