(*blackbox*)
module OTA_2stage (
    inout vdd,
    inout vss,
    output vout,
    input vin1,
    input vin2,
    input vp
);
endmodule // OTA_2stage
