(*blackbox*)
module TopLevel_oscillator (
    inout VP,
    inout GND,
    output Y
);
endmodule // TopLevel_oscillator
