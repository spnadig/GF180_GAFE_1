magic
tech gf180mcuC
magscale 1 10
timestamp 1676577649
<< error_p >>
rect -66 0 -64 20000
rect 0 0 2 20000
<< nwell >>
rect -176 -86 24558 20086
<< pmos >>
rect 88 0 228 20000
rect 332 0 472 20000
rect 576 0 716 20000
rect 820 0 960 20000
rect 1064 0 1204 20000
rect 1308 0 1448 20000
rect 1552 0 1692 20000
rect 1796 0 1936 20000
rect 2040 0 2180 20000
rect 2284 0 2424 20000
rect 2528 0 2668 20000
rect 2772 0 2912 20000
rect 3016 0 3156 20000
rect 3260 0 3400 20000
rect 3504 0 3644 20000
rect 3748 0 3888 20000
rect 3992 0 4132 20000
rect 4236 0 4376 20000
rect 4480 0 4620 20000
rect 4724 0 4864 20000
rect 4968 0 5108 20000
rect 5212 0 5352 20000
rect 5456 0 5596 20000
rect 5700 0 5840 20000
rect 5944 0 6084 20000
rect 6188 0 6328 20000
rect 6432 0 6572 20000
rect 6676 0 6816 20000
rect 6920 0 7060 20000
rect 7164 0 7304 20000
rect 7408 0 7548 20000
rect 7652 0 7792 20000
rect 7896 0 8036 20000
rect 8140 0 8280 20000
rect 8384 0 8524 20000
rect 8628 0 8768 20000
rect 8872 0 9012 20000
rect 9116 0 9256 20000
rect 9360 0 9500 20000
rect 9604 0 9744 20000
rect 9848 0 9988 20000
rect 10092 0 10232 20000
rect 10336 0 10476 20000
rect 10580 0 10720 20000
rect 10824 0 10964 20000
rect 11068 0 11208 20000
rect 11312 0 11452 20000
rect 11556 0 11696 20000
rect 11800 0 11940 20000
rect 12044 0 12184 20000
rect 12288 0 12428 20000
rect 12532 0 12672 20000
rect 12776 0 12916 20000
rect 13020 0 13160 20000
rect 13264 0 13404 20000
rect 13508 0 13648 20000
rect 13752 0 13892 20000
rect 13996 0 14136 20000
rect 14240 0 14380 20000
rect 14484 0 14624 20000
rect 14728 0 14868 20000
rect 14972 0 15112 20000
rect 15216 0 15356 20000
rect 15460 0 15600 20000
rect 15704 0 15844 20000
rect 15948 0 16088 20000
rect 16192 0 16332 20000
rect 16436 0 16576 20000
rect 16680 0 16820 20000
rect 16924 0 17064 20000
rect 17168 0 17308 20000
rect 17412 0 17552 20000
rect 17656 0 17796 20000
rect 17900 0 18040 20000
rect 18144 0 18284 20000
rect 18388 0 18528 20000
rect 18632 0 18772 20000
rect 18876 0 19016 20000
rect 19120 0 19260 20000
rect 19364 0 19504 20000
rect 19608 0 19748 20000
rect 19852 0 19992 20000
rect 20096 0 20236 20000
rect 20340 0 20480 20000
rect 20584 0 20724 20000
rect 20828 0 20968 20000
rect 21072 0 21212 20000
rect 21316 0 21456 20000
rect 21560 0 21700 20000
rect 21804 0 21944 20000
rect 22048 0 22188 20000
rect 22292 0 22432 20000
rect 22536 0 22676 20000
rect 22780 0 22920 20000
rect 23024 0 23164 20000
rect 23268 0 23408 20000
rect 23512 0 23652 20000
rect 23756 0 23896 20000
rect 24000 0 24140 20000
rect 24244 0 24384 20000
<< pdiff >>
rect 0 19973 88 20000
rect 0 27 13 19973
rect 59 27 88 19973
rect 0 0 88 27
rect 228 19973 332 20000
rect 228 27 257 19973
rect 303 27 332 19973
rect 228 0 332 27
rect 472 19973 576 20000
rect 472 27 501 19973
rect 547 27 576 19973
rect 472 0 576 27
rect 716 19973 820 20000
rect 716 27 745 19973
rect 791 27 820 19973
rect 716 0 820 27
rect 960 19973 1064 20000
rect 960 27 989 19973
rect 1035 27 1064 19973
rect 960 0 1064 27
rect 1204 19973 1308 20000
rect 1204 27 1233 19973
rect 1279 27 1308 19973
rect 1204 0 1308 27
rect 1448 19973 1552 20000
rect 1448 27 1477 19973
rect 1523 27 1552 19973
rect 1448 0 1552 27
rect 1692 19973 1796 20000
rect 1692 27 1721 19973
rect 1767 27 1796 19973
rect 1692 0 1796 27
rect 1936 19973 2040 20000
rect 1936 27 1965 19973
rect 2011 27 2040 19973
rect 1936 0 2040 27
rect 2180 19973 2284 20000
rect 2180 27 2209 19973
rect 2255 27 2284 19973
rect 2180 0 2284 27
rect 2424 19973 2528 20000
rect 2424 27 2453 19973
rect 2499 27 2528 19973
rect 2424 0 2528 27
rect 2668 19973 2772 20000
rect 2668 27 2697 19973
rect 2743 27 2772 19973
rect 2668 0 2772 27
rect 2912 19973 3016 20000
rect 2912 27 2941 19973
rect 2987 27 3016 19973
rect 2912 0 3016 27
rect 3156 19973 3260 20000
rect 3156 27 3185 19973
rect 3231 27 3260 19973
rect 3156 0 3260 27
rect 3400 19973 3504 20000
rect 3400 27 3429 19973
rect 3475 27 3504 19973
rect 3400 0 3504 27
rect 3644 19973 3748 20000
rect 3644 27 3673 19973
rect 3719 27 3748 19973
rect 3644 0 3748 27
rect 3888 19973 3992 20000
rect 3888 27 3917 19973
rect 3963 27 3992 19973
rect 3888 0 3992 27
rect 4132 19973 4236 20000
rect 4132 27 4161 19973
rect 4207 27 4236 19973
rect 4132 0 4236 27
rect 4376 19973 4480 20000
rect 4376 27 4405 19973
rect 4451 27 4480 19973
rect 4376 0 4480 27
rect 4620 19973 4724 20000
rect 4620 27 4649 19973
rect 4695 27 4724 19973
rect 4620 0 4724 27
rect 4864 19973 4968 20000
rect 4864 27 4893 19973
rect 4939 27 4968 19973
rect 4864 0 4968 27
rect 5108 19973 5212 20000
rect 5108 27 5137 19973
rect 5183 27 5212 19973
rect 5108 0 5212 27
rect 5352 19973 5456 20000
rect 5352 27 5381 19973
rect 5427 27 5456 19973
rect 5352 0 5456 27
rect 5596 19973 5700 20000
rect 5596 27 5625 19973
rect 5671 27 5700 19973
rect 5596 0 5700 27
rect 5840 19973 5944 20000
rect 5840 27 5869 19973
rect 5915 27 5944 19973
rect 5840 0 5944 27
rect 6084 19973 6188 20000
rect 6084 27 6113 19973
rect 6159 27 6188 19973
rect 6084 0 6188 27
rect 6328 19973 6432 20000
rect 6328 27 6357 19973
rect 6403 27 6432 19973
rect 6328 0 6432 27
rect 6572 19973 6676 20000
rect 6572 27 6601 19973
rect 6647 27 6676 19973
rect 6572 0 6676 27
rect 6816 19973 6920 20000
rect 6816 27 6845 19973
rect 6891 27 6920 19973
rect 6816 0 6920 27
rect 7060 19973 7164 20000
rect 7060 27 7089 19973
rect 7135 27 7164 19973
rect 7060 0 7164 27
rect 7304 19973 7408 20000
rect 7304 27 7333 19973
rect 7379 27 7408 19973
rect 7304 0 7408 27
rect 7548 19973 7652 20000
rect 7548 27 7577 19973
rect 7623 27 7652 19973
rect 7548 0 7652 27
rect 7792 19973 7896 20000
rect 7792 27 7821 19973
rect 7867 27 7896 19973
rect 7792 0 7896 27
rect 8036 19973 8140 20000
rect 8036 27 8065 19973
rect 8111 27 8140 19973
rect 8036 0 8140 27
rect 8280 19973 8384 20000
rect 8280 27 8309 19973
rect 8355 27 8384 19973
rect 8280 0 8384 27
rect 8524 19973 8628 20000
rect 8524 27 8553 19973
rect 8599 27 8628 19973
rect 8524 0 8628 27
rect 8768 19973 8872 20000
rect 8768 27 8797 19973
rect 8843 27 8872 19973
rect 8768 0 8872 27
rect 9012 19973 9116 20000
rect 9012 27 9041 19973
rect 9087 27 9116 19973
rect 9012 0 9116 27
rect 9256 19973 9360 20000
rect 9256 27 9285 19973
rect 9331 27 9360 19973
rect 9256 0 9360 27
rect 9500 19973 9604 20000
rect 9500 27 9529 19973
rect 9575 27 9604 19973
rect 9500 0 9604 27
rect 9744 19973 9848 20000
rect 9744 27 9773 19973
rect 9819 27 9848 19973
rect 9744 0 9848 27
rect 9988 19973 10092 20000
rect 9988 27 10017 19973
rect 10063 27 10092 19973
rect 9988 0 10092 27
rect 10232 19973 10336 20000
rect 10232 27 10261 19973
rect 10307 27 10336 19973
rect 10232 0 10336 27
rect 10476 19973 10580 20000
rect 10476 27 10505 19973
rect 10551 27 10580 19973
rect 10476 0 10580 27
rect 10720 19973 10824 20000
rect 10720 27 10749 19973
rect 10795 27 10824 19973
rect 10720 0 10824 27
rect 10964 19973 11068 20000
rect 10964 27 10993 19973
rect 11039 27 11068 19973
rect 10964 0 11068 27
rect 11208 19973 11312 20000
rect 11208 27 11237 19973
rect 11283 27 11312 19973
rect 11208 0 11312 27
rect 11452 19973 11556 20000
rect 11452 27 11481 19973
rect 11527 27 11556 19973
rect 11452 0 11556 27
rect 11696 19973 11800 20000
rect 11696 27 11725 19973
rect 11771 27 11800 19973
rect 11696 0 11800 27
rect 11940 19973 12044 20000
rect 11940 27 11969 19973
rect 12015 27 12044 19973
rect 11940 0 12044 27
rect 12184 19973 12288 20000
rect 12184 27 12213 19973
rect 12259 27 12288 19973
rect 12184 0 12288 27
rect 12428 19973 12532 20000
rect 12428 27 12457 19973
rect 12503 27 12532 19973
rect 12428 0 12532 27
rect 12672 19973 12776 20000
rect 12672 27 12701 19973
rect 12747 27 12776 19973
rect 12672 0 12776 27
rect 12916 19973 13020 20000
rect 12916 27 12945 19973
rect 12991 27 13020 19973
rect 12916 0 13020 27
rect 13160 19973 13264 20000
rect 13160 27 13189 19973
rect 13235 27 13264 19973
rect 13160 0 13264 27
rect 13404 19973 13508 20000
rect 13404 27 13433 19973
rect 13479 27 13508 19973
rect 13404 0 13508 27
rect 13648 19973 13752 20000
rect 13648 27 13677 19973
rect 13723 27 13752 19973
rect 13648 0 13752 27
rect 13892 19973 13996 20000
rect 13892 27 13921 19973
rect 13967 27 13996 19973
rect 13892 0 13996 27
rect 14136 19973 14240 20000
rect 14136 27 14165 19973
rect 14211 27 14240 19973
rect 14136 0 14240 27
rect 14380 19973 14484 20000
rect 14380 27 14409 19973
rect 14455 27 14484 19973
rect 14380 0 14484 27
rect 14624 19973 14728 20000
rect 14624 27 14653 19973
rect 14699 27 14728 19973
rect 14624 0 14728 27
rect 14868 19973 14972 20000
rect 14868 27 14897 19973
rect 14943 27 14972 19973
rect 14868 0 14972 27
rect 15112 19973 15216 20000
rect 15112 27 15141 19973
rect 15187 27 15216 19973
rect 15112 0 15216 27
rect 15356 19973 15460 20000
rect 15356 27 15385 19973
rect 15431 27 15460 19973
rect 15356 0 15460 27
rect 15600 19973 15704 20000
rect 15600 27 15629 19973
rect 15675 27 15704 19973
rect 15600 0 15704 27
rect 15844 19973 15948 20000
rect 15844 27 15873 19973
rect 15919 27 15948 19973
rect 15844 0 15948 27
rect 16088 19973 16192 20000
rect 16088 27 16117 19973
rect 16163 27 16192 19973
rect 16088 0 16192 27
rect 16332 19973 16436 20000
rect 16332 27 16361 19973
rect 16407 27 16436 19973
rect 16332 0 16436 27
rect 16576 19973 16680 20000
rect 16576 27 16605 19973
rect 16651 27 16680 19973
rect 16576 0 16680 27
rect 16820 19973 16924 20000
rect 16820 27 16849 19973
rect 16895 27 16924 19973
rect 16820 0 16924 27
rect 17064 19973 17168 20000
rect 17064 27 17093 19973
rect 17139 27 17168 19973
rect 17064 0 17168 27
rect 17308 19973 17412 20000
rect 17308 27 17337 19973
rect 17383 27 17412 19973
rect 17308 0 17412 27
rect 17552 19973 17656 20000
rect 17552 27 17581 19973
rect 17627 27 17656 19973
rect 17552 0 17656 27
rect 17796 19973 17900 20000
rect 17796 27 17825 19973
rect 17871 27 17900 19973
rect 17796 0 17900 27
rect 18040 19973 18144 20000
rect 18040 27 18069 19973
rect 18115 27 18144 19973
rect 18040 0 18144 27
rect 18284 19973 18388 20000
rect 18284 27 18313 19973
rect 18359 27 18388 19973
rect 18284 0 18388 27
rect 18528 19973 18632 20000
rect 18528 27 18557 19973
rect 18603 27 18632 19973
rect 18528 0 18632 27
rect 18772 19973 18876 20000
rect 18772 27 18801 19973
rect 18847 27 18876 19973
rect 18772 0 18876 27
rect 19016 19973 19120 20000
rect 19016 27 19045 19973
rect 19091 27 19120 19973
rect 19016 0 19120 27
rect 19260 19973 19364 20000
rect 19260 27 19289 19973
rect 19335 27 19364 19973
rect 19260 0 19364 27
rect 19504 19973 19608 20000
rect 19504 27 19533 19973
rect 19579 27 19608 19973
rect 19504 0 19608 27
rect 19748 19973 19852 20000
rect 19748 27 19777 19973
rect 19823 27 19852 19973
rect 19748 0 19852 27
rect 19992 19973 20096 20000
rect 19992 27 20021 19973
rect 20067 27 20096 19973
rect 19992 0 20096 27
rect 20236 19973 20340 20000
rect 20236 27 20265 19973
rect 20311 27 20340 19973
rect 20236 0 20340 27
rect 20480 19973 20584 20000
rect 20480 27 20509 19973
rect 20555 27 20584 19973
rect 20480 0 20584 27
rect 20724 19973 20828 20000
rect 20724 27 20753 19973
rect 20799 27 20828 19973
rect 20724 0 20828 27
rect 20968 19973 21072 20000
rect 20968 27 20997 19973
rect 21043 27 21072 19973
rect 20968 0 21072 27
rect 21212 19973 21316 20000
rect 21212 27 21241 19973
rect 21287 27 21316 19973
rect 21212 0 21316 27
rect 21456 19973 21560 20000
rect 21456 27 21485 19973
rect 21531 27 21560 19973
rect 21456 0 21560 27
rect 21700 19973 21804 20000
rect 21700 27 21729 19973
rect 21775 27 21804 19973
rect 21700 0 21804 27
rect 21944 19973 22048 20000
rect 21944 27 21973 19973
rect 22019 27 22048 19973
rect 21944 0 22048 27
rect 22188 19973 22292 20000
rect 22188 27 22217 19973
rect 22263 27 22292 19973
rect 22188 0 22292 27
rect 22432 19973 22536 20000
rect 22432 27 22461 19973
rect 22507 27 22536 19973
rect 22432 0 22536 27
rect 22676 19973 22780 20000
rect 22676 27 22705 19973
rect 22751 27 22780 19973
rect 22676 0 22780 27
rect 22920 19973 23024 20000
rect 22920 27 22949 19973
rect 22995 27 23024 19973
rect 22920 0 23024 27
rect 23164 19973 23268 20000
rect 23164 27 23193 19973
rect 23239 27 23268 19973
rect 23164 0 23268 27
rect 23408 19973 23512 20000
rect 23408 27 23437 19973
rect 23483 27 23512 19973
rect 23408 0 23512 27
rect 23652 19973 23756 20000
rect 23652 27 23681 19973
rect 23727 27 23756 19973
rect 23652 0 23756 27
rect 23896 19973 24000 20000
rect 23896 27 23925 19973
rect 23971 27 24000 19973
rect 23896 0 24000 27
rect 24140 19973 24244 20000
rect 24140 27 24169 19973
rect 24215 27 24244 19973
rect 24140 0 24244 27
rect 24384 19973 24472 20000
rect 24384 27 24413 19973
rect 24459 27 24472 19973
rect 24384 0 24472 27
<< pdiffc >>
rect 13 27 59 19973
rect 257 27 303 19973
rect 501 27 547 19973
rect 745 27 791 19973
rect 989 27 1035 19973
rect 1233 27 1279 19973
rect 1477 27 1523 19973
rect 1721 27 1767 19973
rect 1965 27 2011 19973
rect 2209 27 2255 19973
rect 2453 27 2499 19973
rect 2697 27 2743 19973
rect 2941 27 2987 19973
rect 3185 27 3231 19973
rect 3429 27 3475 19973
rect 3673 27 3719 19973
rect 3917 27 3963 19973
rect 4161 27 4207 19973
rect 4405 27 4451 19973
rect 4649 27 4695 19973
rect 4893 27 4939 19973
rect 5137 27 5183 19973
rect 5381 27 5427 19973
rect 5625 27 5671 19973
rect 5869 27 5915 19973
rect 6113 27 6159 19973
rect 6357 27 6403 19973
rect 6601 27 6647 19973
rect 6845 27 6891 19973
rect 7089 27 7135 19973
rect 7333 27 7379 19973
rect 7577 27 7623 19973
rect 7821 27 7867 19973
rect 8065 27 8111 19973
rect 8309 27 8355 19973
rect 8553 27 8599 19973
rect 8797 27 8843 19973
rect 9041 27 9087 19973
rect 9285 27 9331 19973
rect 9529 27 9575 19973
rect 9773 27 9819 19973
rect 10017 27 10063 19973
rect 10261 27 10307 19973
rect 10505 27 10551 19973
rect 10749 27 10795 19973
rect 10993 27 11039 19973
rect 11237 27 11283 19973
rect 11481 27 11527 19973
rect 11725 27 11771 19973
rect 11969 27 12015 19973
rect 12213 27 12259 19973
rect 12457 27 12503 19973
rect 12701 27 12747 19973
rect 12945 27 12991 19973
rect 13189 27 13235 19973
rect 13433 27 13479 19973
rect 13677 27 13723 19973
rect 13921 27 13967 19973
rect 14165 27 14211 19973
rect 14409 27 14455 19973
rect 14653 27 14699 19973
rect 14897 27 14943 19973
rect 15141 27 15187 19973
rect 15385 27 15431 19973
rect 15629 27 15675 19973
rect 15873 27 15919 19973
rect 16117 27 16163 19973
rect 16361 27 16407 19973
rect 16605 27 16651 19973
rect 16849 27 16895 19973
rect 17093 27 17139 19973
rect 17337 27 17383 19973
rect 17581 27 17627 19973
rect 17825 27 17871 19973
rect 18069 27 18115 19973
rect 18313 27 18359 19973
rect 18557 27 18603 19973
rect 18801 27 18847 19973
rect 19045 27 19091 19973
rect 19289 27 19335 19973
rect 19533 27 19579 19973
rect 19777 27 19823 19973
rect 20021 27 20067 19973
rect 20265 27 20311 19973
rect 20509 27 20555 19973
rect 20753 27 20799 19973
rect 20997 27 21043 19973
rect 21241 27 21287 19973
rect 21485 27 21531 19973
rect 21729 27 21775 19973
rect 21973 27 22019 19973
rect 22217 27 22263 19973
rect 22461 27 22507 19973
rect 22705 27 22751 19973
rect 22949 27 22995 19973
rect 23193 27 23239 19973
rect 23437 27 23483 19973
rect 23681 27 23727 19973
rect 23925 27 23971 19973
rect 24169 27 24215 19973
rect 24413 27 24459 19973
<< nsubdiff >>
rect -152 19973 -64 20000
rect -152 27 -131 19973
rect -85 27 -64 19973
rect -152 0 -64 27
<< nsubdiffcont >>
rect -131 27 -85 19973
<< polysilicon >>
rect 88 20000 228 20044
rect 332 20000 472 20044
rect 576 20000 716 20044
rect 820 20000 960 20044
rect 1064 20000 1204 20044
rect 1308 20000 1448 20044
rect 1552 20000 1692 20044
rect 1796 20000 1936 20044
rect 2040 20000 2180 20044
rect 2284 20000 2424 20044
rect 2528 20000 2668 20044
rect 2772 20000 2912 20044
rect 3016 20000 3156 20044
rect 3260 20000 3400 20044
rect 3504 20000 3644 20044
rect 3748 20000 3888 20044
rect 3992 20000 4132 20044
rect 4236 20000 4376 20044
rect 4480 20000 4620 20044
rect 4724 20000 4864 20044
rect 4968 20000 5108 20044
rect 5212 20000 5352 20044
rect 5456 20000 5596 20044
rect 5700 20000 5840 20044
rect 5944 20000 6084 20044
rect 6188 20000 6328 20044
rect 6432 20000 6572 20044
rect 6676 20000 6816 20044
rect 6920 20000 7060 20044
rect 7164 20000 7304 20044
rect 7408 20000 7548 20044
rect 7652 20000 7792 20044
rect 7896 20000 8036 20044
rect 8140 20000 8280 20044
rect 8384 20000 8524 20044
rect 8628 20000 8768 20044
rect 8872 20000 9012 20044
rect 9116 20000 9256 20044
rect 9360 20000 9500 20044
rect 9604 20000 9744 20044
rect 9848 20000 9988 20044
rect 10092 20000 10232 20044
rect 10336 20000 10476 20044
rect 10580 20000 10720 20044
rect 10824 20000 10964 20044
rect 11068 20000 11208 20044
rect 11312 20000 11452 20044
rect 11556 20000 11696 20044
rect 11800 20000 11940 20044
rect 12044 20000 12184 20044
rect 12288 20000 12428 20044
rect 12532 20000 12672 20044
rect 12776 20000 12916 20044
rect 13020 20000 13160 20044
rect 13264 20000 13404 20044
rect 13508 20000 13648 20044
rect 13752 20000 13892 20044
rect 13996 20000 14136 20044
rect 14240 20000 14380 20044
rect 14484 20000 14624 20044
rect 14728 20000 14868 20044
rect 14972 20000 15112 20044
rect 15216 20000 15356 20044
rect 15460 20000 15600 20044
rect 15704 20000 15844 20044
rect 15948 20000 16088 20044
rect 16192 20000 16332 20044
rect 16436 20000 16576 20044
rect 16680 20000 16820 20044
rect 16924 20000 17064 20044
rect 17168 20000 17308 20044
rect 17412 20000 17552 20044
rect 17656 20000 17796 20044
rect 17900 20000 18040 20044
rect 18144 20000 18284 20044
rect 18388 20000 18528 20044
rect 18632 20000 18772 20044
rect 18876 20000 19016 20044
rect 19120 20000 19260 20044
rect 19364 20000 19504 20044
rect 19608 20000 19748 20044
rect 19852 20000 19992 20044
rect 20096 20000 20236 20044
rect 20340 20000 20480 20044
rect 20584 20000 20724 20044
rect 20828 20000 20968 20044
rect 21072 20000 21212 20044
rect 21316 20000 21456 20044
rect 21560 20000 21700 20044
rect 21804 20000 21944 20044
rect 22048 20000 22188 20044
rect 22292 20000 22432 20044
rect 22536 20000 22676 20044
rect 22780 20000 22920 20044
rect 23024 20000 23164 20044
rect 23268 20000 23408 20044
rect 23512 20000 23652 20044
rect 23756 20000 23896 20044
rect 24000 20000 24140 20044
rect 24244 20000 24384 20044
rect 88 -44 228 0
rect 332 -44 472 0
rect 576 -44 716 0
rect 820 -44 960 0
rect 1064 -44 1204 0
rect 1308 -44 1448 0
rect 1552 -44 1692 0
rect 1796 -44 1936 0
rect 2040 -44 2180 0
rect 2284 -44 2424 0
rect 2528 -44 2668 0
rect 2772 -44 2912 0
rect 3016 -44 3156 0
rect 3260 -44 3400 0
rect 3504 -44 3644 0
rect 3748 -44 3888 0
rect 3992 -44 4132 0
rect 4236 -44 4376 0
rect 4480 -44 4620 0
rect 4724 -44 4864 0
rect 4968 -44 5108 0
rect 5212 -44 5352 0
rect 5456 -44 5596 0
rect 5700 -44 5840 0
rect 5944 -44 6084 0
rect 6188 -44 6328 0
rect 6432 -44 6572 0
rect 6676 -44 6816 0
rect 6920 -44 7060 0
rect 7164 -44 7304 0
rect 7408 -44 7548 0
rect 7652 -44 7792 0
rect 7896 -44 8036 0
rect 8140 -44 8280 0
rect 8384 -44 8524 0
rect 8628 -44 8768 0
rect 8872 -44 9012 0
rect 9116 -44 9256 0
rect 9360 -44 9500 0
rect 9604 -44 9744 0
rect 9848 -44 9988 0
rect 10092 -44 10232 0
rect 10336 -44 10476 0
rect 10580 -44 10720 0
rect 10824 -44 10964 0
rect 11068 -44 11208 0
rect 11312 -44 11452 0
rect 11556 -44 11696 0
rect 11800 -44 11940 0
rect 12044 -44 12184 0
rect 12288 -44 12428 0
rect 12532 -44 12672 0
rect 12776 -44 12916 0
rect 13020 -44 13160 0
rect 13264 -44 13404 0
rect 13508 -44 13648 0
rect 13752 -44 13892 0
rect 13996 -44 14136 0
rect 14240 -44 14380 0
rect 14484 -44 14624 0
rect 14728 -44 14868 0
rect 14972 -44 15112 0
rect 15216 -44 15356 0
rect 15460 -44 15600 0
rect 15704 -44 15844 0
rect 15948 -44 16088 0
rect 16192 -44 16332 0
rect 16436 -44 16576 0
rect 16680 -44 16820 0
rect 16924 -44 17064 0
rect 17168 -44 17308 0
rect 17412 -44 17552 0
rect 17656 -44 17796 0
rect 17900 -44 18040 0
rect 18144 -44 18284 0
rect 18388 -44 18528 0
rect 18632 -44 18772 0
rect 18876 -44 19016 0
rect 19120 -44 19260 0
rect 19364 -44 19504 0
rect 19608 -44 19748 0
rect 19852 -44 19992 0
rect 20096 -44 20236 0
rect 20340 -44 20480 0
rect 20584 -44 20724 0
rect 20828 -44 20968 0
rect 21072 -44 21212 0
rect 21316 -44 21456 0
rect 21560 -44 21700 0
rect 21804 -44 21944 0
rect 22048 -44 22188 0
rect 22292 -44 22432 0
rect 22536 -44 22676 0
rect 22780 -44 22920 0
rect 23024 -44 23164 0
rect 23268 -44 23408 0
rect 23512 -44 23652 0
rect 23756 -44 23896 0
rect 24000 -44 24140 0
rect 24244 -44 24384 0
<< metal1 >>
rect -152 19973 -64 20000
rect -152 27 -131 19973
rect -85 27 -64 19973
rect -152 0 -64 27
rect -2 19973 74 20002
rect -2 27 13 19973
rect 59 27 74 19973
rect -2 -2 74 27
rect 242 19973 318 20002
rect 242 27 257 19973
rect 303 27 318 19973
rect 242 -2 318 27
rect 486 19973 562 20002
rect 486 27 501 19973
rect 547 27 562 19973
rect 486 -2 562 27
rect 730 19973 806 20002
rect 730 27 745 19973
rect 791 27 806 19973
rect 730 -2 806 27
rect 974 19973 1050 20002
rect 974 27 989 19973
rect 1035 27 1050 19973
rect 974 -2 1050 27
rect 1218 19973 1294 20002
rect 1218 27 1233 19973
rect 1279 27 1294 19973
rect 1218 -2 1294 27
rect 1462 19973 1538 20002
rect 1462 27 1477 19973
rect 1523 27 1538 19973
rect 1462 -2 1538 27
rect 1706 19973 1782 20002
rect 1706 27 1721 19973
rect 1767 27 1782 19973
rect 1706 -2 1782 27
rect 1950 19973 2026 20002
rect 1950 27 1965 19973
rect 2011 27 2026 19973
rect 1950 -2 2026 27
rect 2194 19973 2270 20002
rect 2194 27 2209 19973
rect 2255 27 2270 19973
rect 2194 -2 2270 27
rect 2438 19973 2514 20002
rect 2438 27 2453 19973
rect 2499 27 2514 19973
rect 2438 -2 2514 27
rect 2682 19973 2758 20002
rect 2682 27 2697 19973
rect 2743 27 2758 19973
rect 2682 -2 2758 27
rect 2926 19973 3002 20002
rect 2926 27 2941 19973
rect 2987 27 3002 19973
rect 2926 -2 3002 27
rect 3170 19973 3246 20002
rect 3170 27 3185 19973
rect 3231 27 3246 19973
rect 3170 -2 3246 27
rect 3414 19973 3490 20002
rect 3414 27 3429 19973
rect 3475 27 3490 19973
rect 3414 -2 3490 27
rect 3658 19973 3734 20002
rect 3658 27 3673 19973
rect 3719 27 3734 19973
rect 3658 -2 3734 27
rect 3902 19973 3978 20002
rect 3902 27 3917 19973
rect 3963 27 3978 19973
rect 3902 -2 3978 27
rect 4146 19973 4222 20002
rect 4146 27 4161 19973
rect 4207 27 4222 19973
rect 4146 -2 4222 27
rect 4390 19973 4466 20002
rect 4390 27 4405 19973
rect 4451 27 4466 19973
rect 4390 -2 4466 27
rect 4634 19973 4710 20002
rect 4634 27 4649 19973
rect 4695 27 4710 19973
rect 4634 -2 4710 27
rect 4878 19973 4954 20002
rect 4878 27 4893 19973
rect 4939 27 4954 19973
rect 4878 -2 4954 27
rect 5122 19973 5198 20002
rect 5122 27 5137 19973
rect 5183 27 5198 19973
rect 5122 -2 5198 27
rect 5366 19973 5442 20002
rect 5366 27 5381 19973
rect 5427 27 5442 19973
rect 5366 -2 5442 27
rect 5610 19973 5686 20002
rect 5610 27 5625 19973
rect 5671 27 5686 19973
rect 5610 -2 5686 27
rect 5854 19973 5930 20002
rect 5854 27 5869 19973
rect 5915 27 5930 19973
rect 5854 -2 5930 27
rect 6098 19973 6174 20002
rect 6098 27 6113 19973
rect 6159 27 6174 19973
rect 6098 -2 6174 27
rect 6342 19973 6418 20002
rect 6342 27 6357 19973
rect 6403 27 6418 19973
rect 6342 -2 6418 27
rect 6586 19973 6662 20002
rect 6586 27 6601 19973
rect 6647 27 6662 19973
rect 6586 -2 6662 27
rect 6830 19973 6906 20002
rect 6830 27 6845 19973
rect 6891 27 6906 19973
rect 6830 -2 6906 27
rect 7074 19973 7150 20002
rect 7074 27 7089 19973
rect 7135 27 7150 19973
rect 7074 -2 7150 27
rect 7318 19973 7394 20002
rect 7318 27 7333 19973
rect 7379 27 7394 19973
rect 7318 -2 7394 27
rect 7562 19973 7638 20002
rect 7562 27 7577 19973
rect 7623 27 7638 19973
rect 7562 -2 7638 27
rect 7806 19973 7882 20002
rect 7806 27 7821 19973
rect 7867 27 7882 19973
rect 7806 -2 7882 27
rect 8050 19973 8126 20002
rect 8050 27 8065 19973
rect 8111 27 8126 19973
rect 8050 -2 8126 27
rect 8294 19973 8370 20002
rect 8294 27 8309 19973
rect 8355 27 8370 19973
rect 8294 -2 8370 27
rect 8538 19973 8614 20002
rect 8538 27 8553 19973
rect 8599 27 8614 19973
rect 8538 -2 8614 27
rect 8782 19973 8858 20002
rect 8782 27 8797 19973
rect 8843 27 8858 19973
rect 8782 -2 8858 27
rect 9026 19973 9102 20002
rect 9026 27 9041 19973
rect 9087 27 9102 19973
rect 9026 -2 9102 27
rect 9270 19973 9346 20002
rect 9270 27 9285 19973
rect 9331 27 9346 19973
rect 9270 -2 9346 27
rect 9514 19973 9590 20002
rect 9514 27 9529 19973
rect 9575 27 9590 19973
rect 9514 -2 9590 27
rect 9758 19973 9834 20002
rect 9758 27 9773 19973
rect 9819 27 9834 19973
rect 9758 -2 9834 27
rect 10002 19973 10078 20002
rect 10002 27 10017 19973
rect 10063 27 10078 19973
rect 10002 -2 10078 27
rect 10246 19973 10322 20002
rect 10246 27 10261 19973
rect 10307 27 10322 19973
rect 10246 -2 10322 27
rect 10490 19973 10566 20002
rect 10490 27 10505 19973
rect 10551 27 10566 19973
rect 10490 -2 10566 27
rect 10734 19973 10810 20002
rect 10734 27 10749 19973
rect 10795 27 10810 19973
rect 10734 -2 10810 27
rect 10978 19973 11054 20002
rect 10978 27 10993 19973
rect 11039 27 11054 19973
rect 10978 -2 11054 27
rect 11222 19973 11298 20002
rect 11222 27 11237 19973
rect 11283 27 11298 19973
rect 11222 -2 11298 27
rect 11466 19973 11542 20002
rect 11466 27 11481 19973
rect 11527 27 11542 19973
rect 11466 -2 11542 27
rect 11710 19973 11786 20002
rect 11710 27 11725 19973
rect 11771 27 11786 19973
rect 11710 -2 11786 27
rect 11954 19973 12030 20002
rect 11954 27 11969 19973
rect 12015 27 12030 19973
rect 11954 -2 12030 27
rect 12198 19973 12274 20002
rect 12198 27 12213 19973
rect 12259 27 12274 19973
rect 12198 -2 12274 27
rect 12442 19973 12518 20002
rect 12442 27 12457 19973
rect 12503 27 12518 19973
rect 12442 -2 12518 27
rect 12686 19973 12762 20002
rect 12686 27 12701 19973
rect 12747 27 12762 19973
rect 12686 -2 12762 27
rect 12930 19973 13006 20002
rect 12930 27 12945 19973
rect 12991 27 13006 19973
rect 12930 -2 13006 27
rect 13174 19973 13250 20002
rect 13174 27 13189 19973
rect 13235 27 13250 19973
rect 13174 -2 13250 27
rect 13418 19973 13494 20002
rect 13418 27 13433 19973
rect 13479 27 13494 19973
rect 13418 -2 13494 27
rect 13662 19973 13738 20002
rect 13662 27 13677 19973
rect 13723 27 13738 19973
rect 13662 -2 13738 27
rect 13906 19973 13982 20002
rect 13906 27 13921 19973
rect 13967 27 13982 19973
rect 13906 -2 13982 27
rect 14150 19973 14226 20002
rect 14150 27 14165 19973
rect 14211 27 14226 19973
rect 14150 -2 14226 27
rect 14394 19973 14470 20002
rect 14394 27 14409 19973
rect 14455 27 14470 19973
rect 14394 -2 14470 27
rect 14638 19973 14714 20002
rect 14638 27 14653 19973
rect 14699 27 14714 19973
rect 14638 -2 14714 27
rect 14882 19973 14958 20002
rect 14882 27 14897 19973
rect 14943 27 14958 19973
rect 14882 -2 14958 27
rect 15126 19973 15202 20002
rect 15126 27 15141 19973
rect 15187 27 15202 19973
rect 15126 -2 15202 27
rect 15370 19973 15446 20002
rect 15370 27 15385 19973
rect 15431 27 15446 19973
rect 15370 -2 15446 27
rect 15614 19973 15690 20002
rect 15614 27 15629 19973
rect 15675 27 15690 19973
rect 15614 -2 15690 27
rect 15858 19973 15934 20002
rect 15858 27 15873 19973
rect 15919 27 15934 19973
rect 15858 -2 15934 27
rect 16102 19973 16178 20002
rect 16102 27 16117 19973
rect 16163 27 16178 19973
rect 16102 -2 16178 27
rect 16346 19973 16422 20002
rect 16346 27 16361 19973
rect 16407 27 16422 19973
rect 16346 -2 16422 27
rect 16590 19973 16666 20002
rect 16590 27 16605 19973
rect 16651 27 16666 19973
rect 16590 -2 16666 27
rect 16834 19973 16910 20002
rect 16834 27 16849 19973
rect 16895 27 16910 19973
rect 16834 -2 16910 27
rect 17078 19973 17154 20002
rect 17078 27 17093 19973
rect 17139 27 17154 19973
rect 17078 -2 17154 27
rect 17322 19973 17398 20002
rect 17322 27 17337 19973
rect 17383 27 17398 19973
rect 17322 -2 17398 27
rect 17566 19973 17642 20002
rect 17566 27 17581 19973
rect 17627 27 17642 19973
rect 17566 -2 17642 27
rect 17810 19973 17886 20002
rect 17810 27 17825 19973
rect 17871 27 17886 19973
rect 17810 -2 17886 27
rect 18054 19973 18130 20002
rect 18054 27 18069 19973
rect 18115 27 18130 19973
rect 18054 -2 18130 27
rect 18298 19973 18374 20002
rect 18298 27 18313 19973
rect 18359 27 18374 19973
rect 18298 -2 18374 27
rect 18542 19973 18618 20002
rect 18542 27 18557 19973
rect 18603 27 18618 19973
rect 18542 -2 18618 27
rect 18786 19973 18862 20002
rect 18786 27 18801 19973
rect 18847 27 18862 19973
rect 18786 -2 18862 27
rect 19030 19973 19106 20002
rect 19030 27 19045 19973
rect 19091 27 19106 19973
rect 19030 -2 19106 27
rect 19274 19973 19350 20002
rect 19274 27 19289 19973
rect 19335 27 19350 19973
rect 19274 -2 19350 27
rect 19518 19973 19594 20002
rect 19518 27 19533 19973
rect 19579 27 19594 19973
rect 19518 -2 19594 27
rect 19762 19973 19838 20002
rect 19762 27 19777 19973
rect 19823 27 19838 19973
rect 19762 -2 19838 27
rect 20006 19973 20082 20002
rect 20006 27 20021 19973
rect 20067 27 20082 19973
rect 20006 -2 20082 27
rect 20250 19973 20326 20002
rect 20250 27 20265 19973
rect 20311 27 20326 19973
rect 20250 -2 20326 27
rect 20494 19973 20570 20002
rect 20494 27 20509 19973
rect 20555 27 20570 19973
rect 20494 -2 20570 27
rect 20738 19973 20814 20002
rect 20738 27 20753 19973
rect 20799 27 20814 19973
rect 20738 -2 20814 27
rect 20982 19973 21058 20002
rect 20982 27 20997 19973
rect 21043 27 21058 19973
rect 20982 -2 21058 27
rect 21226 19973 21302 20002
rect 21226 27 21241 19973
rect 21287 27 21302 19973
rect 21226 -2 21302 27
rect 21470 19973 21546 20002
rect 21470 27 21485 19973
rect 21531 27 21546 19973
rect 21470 -2 21546 27
rect 21714 19973 21790 20002
rect 21714 27 21729 19973
rect 21775 27 21790 19973
rect 21714 -2 21790 27
rect 21958 19973 22034 20002
rect 21958 27 21973 19973
rect 22019 27 22034 19973
rect 21958 -2 22034 27
rect 22202 19973 22278 20002
rect 22202 27 22217 19973
rect 22263 27 22278 19973
rect 22202 -2 22278 27
rect 22446 19973 22522 20002
rect 22446 27 22461 19973
rect 22507 27 22522 19973
rect 22446 -2 22522 27
rect 22690 19973 22766 20002
rect 22690 27 22705 19973
rect 22751 27 22766 19973
rect 22690 -2 22766 27
rect 22934 19973 23010 20002
rect 22934 27 22949 19973
rect 22995 27 23010 19973
rect 22934 -2 23010 27
rect 23178 19973 23254 20002
rect 23178 27 23193 19973
rect 23239 27 23254 19973
rect 23178 -2 23254 27
rect 23422 19973 23498 20002
rect 23422 27 23437 19973
rect 23483 27 23498 19973
rect 23422 -2 23498 27
rect 23666 19973 23742 20002
rect 23666 27 23681 19973
rect 23727 27 23742 19973
rect 23666 -2 23742 27
rect 23910 19973 23986 20002
rect 23910 27 23925 19973
rect 23971 27 23986 19973
rect 23910 -2 23986 27
rect 24154 19973 24230 20002
rect 24154 27 24169 19973
rect 24215 27 24230 19973
rect 24154 -2 24230 27
rect 24398 19973 24474 20002
rect 24398 27 24413 19973
rect 24459 27 24474 19973
rect 24398 -2 24474 27
<< end >>
