* Extracted by KLayout with GF180 LVS runset on : 07/02/2023 19:17

.SUBCKT TopLevel_oscillator
X$1 \$5 \$3 \$1 \$2 inverter
X$2 \$4 \$5 \$1 \$2 inverter
X$3 \$3 \$4 \$1 \$2 inverter
.ENDS TopLevel_oscillator

.SUBCKT inverter \$1 \$2 \$3 \$4
M$1 \$3 \$1 \$2 \$3 pfet_03v3_dn L=5U W=0.5U AS=0.22P AD=0.22P PS=1.88U PD=1.88U
M$2 \$4 \$1 \$2 \$4 nfet_03v3_dn L=5U W=0.5U AS=0.22P AD=0.22P PS=1.88U PD=1.88U
.ENDS inverter
